//  A testbench for UART-RX_en_tb
`timescale 1us/1ns

module UART-RX_en_tb;
    reg RX;
    reg clk16;
    reg CDP;
    reg en;
    wire [7:0] DATA;
    wire DP;
    wire busy;

  \UART-RX  \UART-RX 0 (
    .RX(RX),
    .clk16(clk16),
    .CDP(CDP),
    .en(en),
    .DATA(DATA),
    .DP(DP),
    .busy(busy)
  );

    reg [12:0] patterns[0:7694];
    integer i;

    initial begin
      patterns[0] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[1] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[2] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[3] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[4] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[5] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[6] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[7] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[8] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[9] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[10] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[11] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[12] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[13] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[14] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[15] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[16] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[17] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[18] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[19] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[20] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[21] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[22] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[23] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[24] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[25] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[26] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[27] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[28] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[29] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[30] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[31] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[32] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[33] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[34] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[35] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[36] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[37] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[38] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[39] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[40] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[41] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[42] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[43] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[44] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[45] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[46] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[47] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[48] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[49] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[50] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[51] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[52] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[53] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[54] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[55] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[56] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[57] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[58] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[59] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[60] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[61] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[62] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[63] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[64] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[65] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[66] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[67] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[68] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[69] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[70] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[71] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[72] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[73] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[74] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[75] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[76] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[77] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[78] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[79] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[80] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[81] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[82] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[83] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[84] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[85] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[86] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[87] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[88] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[89] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[90] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[91] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[92] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[93] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[94] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[95] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[96] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[97] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[98] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[99] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[100] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[101] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[102] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[103] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[104] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[105] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[106] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[107] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[108] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[109] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[110] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[111] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[112] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[113] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[114] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[115] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[116] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[117] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[118] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[119] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[120] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[121] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[122] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[123] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[124] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[125] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[126] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[127] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[128] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[129] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[130] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[131] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[132] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[133] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[134] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[135] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[136] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[137] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[138] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[139] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[140] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[141] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[142] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[143] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[144] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[145] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[146] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[147] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[148] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[149] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[150] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[151] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[152] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[153] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[154] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[155] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[156] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[157] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[158] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[159] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[160] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[161] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[162] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[163] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[164] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[165] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[166] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[167] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[168] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[169] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[170] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[171] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[172] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[173] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[174] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[175] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[176] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[177] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[178] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[179] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[180] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[181] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[182] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[183] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[184] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[185] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[186] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[187] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[188] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[189] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[190] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[191] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[192] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[193] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[194] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[195] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[196] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[197] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[198] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[199] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[200] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[201] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[202] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[203] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[204] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[205] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[206] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[207] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[208] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[209] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[210] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[211] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[212] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[213] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[214] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[215] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[216] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[217] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[218] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[219] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[220] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[221] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[222] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[223] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[224] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[225] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[226] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[227] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[228] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[229] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[230] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[231] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[232] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[233] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[234] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[235] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[236] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[237] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[238] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[239] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[240] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[241] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[242] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[243] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[244] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[245] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[246] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[247] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[248] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[249] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[250] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[251] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[252] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[253] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[254] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[255] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[256] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[257] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[258] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[259] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[260] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[261] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[262] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[263] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[264] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[265] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[266] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[267] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[268] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[269] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[270] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[271] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[272] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[273] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[274] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[275] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[276] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[277] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[278] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[279] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[280] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[281] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[282] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[283] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[284] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[285] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[286] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[287] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[288] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[289] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[290] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[291] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[292] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[293] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[294] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[295] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[296] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[297] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[298] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[299] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[300] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[301] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[302] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[303] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[304] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[305] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[306] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[307] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[308] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[309] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[310] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[311] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[312] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[313] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[314] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[315] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[316] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[317] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[318] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[319] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[320] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[321] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[322] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[323] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[324] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[325] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[326] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[327] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[328] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[329] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[330] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[331] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[332] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[333] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[334] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[335] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[336] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[337] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[338] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[339] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[340] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[341] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[342] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[343] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[344] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[345] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[346] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[347] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[348] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[349] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[350] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[351] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[352] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[353] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[354] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[355] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[356] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[357] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[358] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[359] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[360] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[361] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[362] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[363] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[364] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[365] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[366] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[367] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[368] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[369] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[370] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[371] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[372] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[373] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[374] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[375] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[376] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[377] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[378] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[379] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[380] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[381] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[382] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[383] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[384] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[385] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[386] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[387] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[388] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[389] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[390] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[391] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[392] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[393] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[394] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[395] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[396] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[397] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[398] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[399] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[400] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[401] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[402] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[403] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[404] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[405] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[406] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[407] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[408] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[409] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[410] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[411] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[412] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[413] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[414] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[415] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[416] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[417] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[418] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[419] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[420] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[421] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[422] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[423] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[424] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[425] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[426] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[427] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[428] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[429] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[430] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[431] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[432] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[433] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[434] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[435] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[436] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[437] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[438] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[439] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[440] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[441] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[442] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[443] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[444] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[445] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[446] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[447] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[448] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[449] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[450] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[451] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[452] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[453] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[454] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[455] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[456] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[457] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[458] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[459] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[460] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[461] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[462] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[463] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[464] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[465] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[466] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[467] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[468] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[469] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[470] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[471] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[472] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[473] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[474] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[475] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[476] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[477] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[478] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[479] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[480] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[481] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[482] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[483] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[484] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[485] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[486] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[487] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[488] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[489] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[490] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[491] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[492] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[493] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[494] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[495] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[496] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[497] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[498] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[499] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[500] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[501] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[502] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[503] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[504] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[505] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[506] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[507] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[508] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[509] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[510] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[511] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[512] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[513] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[514] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[515] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[516] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[517] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[518] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[519] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[520] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[521] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[522] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[523] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[524] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[525] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[526] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[527] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[528] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[529] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[530] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[531] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[532] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[533] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[534] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[535] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[536] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[537] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[538] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[539] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[540] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[541] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[542] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[543] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[544] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[545] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[546] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[547] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[548] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[549] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[550] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[551] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[552] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[553] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[554] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[555] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[556] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[557] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[558] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[559] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[560] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[561] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[562] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[563] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[564] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[565] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[566] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[567] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[568] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[569] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[570] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[571] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[572] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[573] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[574] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[575] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[576] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[577] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[578] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[579] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[580] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[581] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[582] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[583] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[584] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[585] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[586] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[587] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[588] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[589] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[590] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[591] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[592] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[593] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[594] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[595] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[596] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[597] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[598] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[599] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[600] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[601] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[602] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[603] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[604] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[605] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[606] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[607] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[608] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[609] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[610] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[611] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[612] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[613] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[614] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[615] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[616] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[617] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[618] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[619] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[620] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[621] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[622] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[623] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[624] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[625] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[626] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[627] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[628] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[629] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[630] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[631] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[632] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[633] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[634] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[635] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[636] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[637] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[638] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[639] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[640] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[641] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[642] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[643] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[644] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[645] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[646] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[647] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[648] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[649] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[650] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[651] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[652] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[653] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[654] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[655] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[656] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[657] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[658] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[659] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[660] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[661] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[662] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[663] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[664] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[665] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[666] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[667] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[668] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[669] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[670] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[671] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[672] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[673] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[674] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[675] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[676] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[677] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[678] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[679] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[680] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[681] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[682] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[683] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[684] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[685] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[686] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[687] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[688] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[689] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[690] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[691] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[692] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[693] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[694] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[695] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[696] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[697] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[698] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[699] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[700] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[701] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[702] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[703] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[704] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[705] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[706] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[707] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[708] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[709] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[710] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[711] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[712] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[713] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[714] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[715] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[716] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[717] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[718] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[719] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[720] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[721] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[722] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[723] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[724] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[725] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[726] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[727] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[728] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[729] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[730] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[731] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[732] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[733] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[734] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[735] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[736] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[737] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[738] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[739] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[740] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[741] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[742] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[743] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[744] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[745] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[746] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[747] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[748] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[749] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[750] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[751] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[752] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[753] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[754] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[755] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[756] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[757] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[758] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[759] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[760] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[761] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[762] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[763] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[764] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[765] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[766] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[767] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[768] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[769] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[770] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[771] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[772] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[773] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[774] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[775] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[776] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[777] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[778] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[779] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[780] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[781] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[782] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[783] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[784] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[785] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[786] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[787] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[788] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[789] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[790] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[791] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[792] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[793] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[794] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[795] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[796] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[797] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[798] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[799] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[800] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[801] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[802] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[803] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[804] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[805] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[806] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[807] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[808] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[809] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[810] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[811] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[812] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[813] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[814] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[815] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[816] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[817] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[818] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[819] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[820] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[821] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[822] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[823] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[824] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[825] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[826] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[827] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[828] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[829] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[830] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[831] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[832] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[833] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[834] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[835] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[836] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[837] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[838] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[839] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[840] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[841] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[842] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[843] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[844] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[845] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[846] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[847] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[848] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[849] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[850] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[851] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[852] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[853] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[854] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[855] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[856] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[857] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[858] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[859] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[860] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[861] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[862] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[863] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[864] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[865] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[866] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[867] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[868] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[869] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[870] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[871] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[872] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[873] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[874] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[875] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[876] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[877] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[878] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[879] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[880] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[881] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[882] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[883] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[884] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[885] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[886] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[887] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[888] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[889] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[890] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[891] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[892] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[893] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[894] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[895] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[896] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[897] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[898] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[899] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[900] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[901] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[902] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[903] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[904] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[905] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[906] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[907] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[908] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[909] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[910] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[911] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[912] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[913] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[914] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[915] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[916] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[917] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[918] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[919] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[920] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[921] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[922] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[923] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[924] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[925] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[926] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[927] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[928] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[929] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[930] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[931] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[932] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[933] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[934] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[935] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[936] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[937] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[938] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[939] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[940] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[941] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[942] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[943] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[944] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[945] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[946] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[947] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[948] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[949] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[950] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[951] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[952] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[953] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[954] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[955] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[956] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[957] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[958] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[959] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[960] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[961] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[962] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[963] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[964] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[965] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[966] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[967] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[968] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[969] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[970] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[971] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[972] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[973] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[974] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[975] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[976] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[977] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[978] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[979] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[980] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[981] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[982] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[983] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[984] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[985] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[986] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[987] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[988] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[989] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[990] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[991] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[992] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[993] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[994] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[995] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[996] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[997] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[998] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[999] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1000] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1001] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1002] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1003] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1004] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1005] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1006] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1007] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1008] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1009] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1010] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1011] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1012] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1013] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1014] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1015] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1016] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1017] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1018] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1019] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1020] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1021] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1022] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1023] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[1024] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[1025] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[1026] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1027] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1028] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1029] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1030] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1031] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1032] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1033] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1034] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1035] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1036] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1037] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1038] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1039] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1040] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1041] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1042] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1043] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1044] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1045] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1046] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1047] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1048] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1049] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1050] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1051] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1052] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1053] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1054] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1055] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1056] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1057] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1058] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1059] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1060] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1061] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1062] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1063] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1064] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1065] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1066] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1067] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1068] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1069] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1070] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1071] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[1072] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[1073] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[1074] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1075] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1076] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1077] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1078] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1079] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1080] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1081] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1082] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1083] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1084] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1085] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1086] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1087] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1088] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1089] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1090] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1091] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1092] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1093] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1094] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1095] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1096] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1097] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1098] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1099] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1100] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1101] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1102] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1103] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1104] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1105] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1106] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1107] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1108] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1109] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1110] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1111] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1112] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1113] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1114] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1115] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1116] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1117] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1118] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1119] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[1120] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[1121] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[1122] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1123] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1124] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1125] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1126] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1127] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1128] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1129] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1130] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1131] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1132] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1133] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1134] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1135] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1136] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1137] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1138] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1139] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1140] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1141] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1142] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1143] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1144] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1145] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1146] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1147] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1148] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1149] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1150] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1151] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1152] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1153] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1154] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1155] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1156] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1157] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1158] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1159] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1160] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1161] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1162] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1163] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1164] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1165] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1166] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1167] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[1168] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[1169] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[1170] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1171] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1172] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1173] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1174] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1175] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1176] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1177] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1178] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1179] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1180] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1181] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1182] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1183] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1184] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1185] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1186] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1187] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1188] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1189] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1190] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1191] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1192] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1193] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1194] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1195] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1196] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1197] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1198] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1199] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1200] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1201] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1202] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1203] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1204] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1205] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1206] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1207] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1208] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1209] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1210] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1211] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1212] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1213] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1214] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1215] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[1216] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[1217] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[1218] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1219] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1220] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1221] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1222] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1223] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1224] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1225] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1226] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1227] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1228] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1229] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1230] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1231] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1232] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1233] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1234] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1235] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1236] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1237] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1238] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1239] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1240] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1241] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1242] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1243] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1244] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1245] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1246] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1247] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1248] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1249] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1250] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1251] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1252] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1253] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1254] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1255] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1256] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1257] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1258] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1259] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1260] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1261] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1262] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1263] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[1264] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[1265] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[1266] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1267] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1268] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1269] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1270] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1271] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1272] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1273] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1274] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1275] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1276] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1277] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1278] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1279] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1280] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1281] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1282] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1283] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1284] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1285] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1286] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1287] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1288] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1289] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1290] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1291] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1292] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1293] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1294] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1295] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1296] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1297] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1298] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1299] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1300] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1301] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1302] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1303] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1304] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1305] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1306] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1307] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1308] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1309] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1310] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1311] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[1312] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[1313] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[1314] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1315] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1316] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1317] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1318] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1319] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1320] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1321] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1322] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1323] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1324] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1325] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1326] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1327] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1328] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1329] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1330] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1331] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1332] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1333] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1334] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1335] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1336] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1337] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1338] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1339] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1340] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1341] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1342] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1343] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1344] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1345] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1346] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1347] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1348] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1349] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1350] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1351] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1352] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1353] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1354] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1355] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1356] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1357] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1358] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1359] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[1360] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[1361] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[1362] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1363] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1364] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1365] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1366] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1367] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1368] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1369] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1370] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1371] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1372] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1373] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1374] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1375] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1376] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1377] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1378] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1379] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1380] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1381] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1382] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1383] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1384] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1385] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1386] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1387] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1388] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1389] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1390] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1391] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1392] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1393] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1394] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1395] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1396] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1397] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1398] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1399] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1400] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1401] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1402] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1403] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1404] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1405] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1406] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1407] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[1408] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[1409] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[1410] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1411] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1412] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1413] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1414] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1415] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1416] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1417] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1418] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1419] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1420] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1421] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1422] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1423] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1424] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1425] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1426] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1427] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1428] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1429] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1430] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1431] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1432] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1433] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1434] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1435] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1436] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1437] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1438] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1439] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1440] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1441] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1442] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1443] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1444] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1445] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1446] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1447] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1448] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1449] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1450] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1451] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1452] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1453] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1454] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1455] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[1456] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[1457] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[1458] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1459] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1460] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1461] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1462] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1463] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1464] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1465] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1466] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1467] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1468] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1469] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1470] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1471] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1472] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1473] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1474] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1475] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1476] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1477] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1478] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1479] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1480] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1481] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1482] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1483] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1484] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1485] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1486] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1487] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1488] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1489] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1490] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1491] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1492] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1493] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1494] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1495] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1496] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1497] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1498] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1499] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1500] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1501] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1502] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1503] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[1504] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[1505] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[1506] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1507] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1508] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1509] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1510] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1511] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1512] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1513] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1514] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1515] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1516] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1517] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1518] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1519] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1520] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1521] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1522] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1523] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1524] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1525] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1526] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1527] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1528] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1529] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1530] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1531] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1532] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1533] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1534] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1535] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1536] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1537] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1538] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1539] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1540] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1541] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1542] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1543] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1544] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1545] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1546] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1547] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1548] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[1549] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[1550] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[1551] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[1552] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[1553] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[1554] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1555] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1556] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1557] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1558] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1559] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1560] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1561] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1562] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1563] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1564] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1565] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1566] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1567] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1568] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1569] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1570] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1571] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1572] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1573] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1574] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1575] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1576] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1577] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1578] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1579] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1580] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1581] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1582] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1583] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1584] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1585] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1586] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1587] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1588] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1589] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1590] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1591] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1592] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1593] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1594] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1595] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1596] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1597] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1598] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1599] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[1600] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[1601] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[1602] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1603] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1604] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1605] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1606] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1607] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1608] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1609] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1610] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1611] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1612] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1613] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1614] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1615] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1616] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1617] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1618] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1619] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1620] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1621] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1622] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1623] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1624] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1625] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1626] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1627] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1628] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1629] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1630] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1631] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1632] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1633] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1634] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1635] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1636] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1637] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1638] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1639] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1640] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1641] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1642] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1643] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1644] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1645] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1646] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1647] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[1648] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[1649] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[1650] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1651] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1652] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1653] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1654] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1655] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1656] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1657] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1658] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1659] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1660] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1661] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1662] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1663] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1664] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1665] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1666] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1667] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1668] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1669] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1670] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1671] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1672] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1673] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1674] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1675] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1676] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1677] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1678] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1679] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1680] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1681] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1682] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1683] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1684] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1685] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1686] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1687] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1688] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1689] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1690] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1691] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1692] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1693] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1694] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1695] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[1696] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[1697] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[1698] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1699] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1700] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1701] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1702] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1703] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1704] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1705] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1706] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1707] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1708] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1709] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1710] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1711] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1712] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1713] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1714] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1715] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1716] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1717] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1718] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1719] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1720] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1721] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1722] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1723] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1724] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1725] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1726] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1727] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1728] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1729] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1730] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1731] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1732] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1733] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1734] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1735] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1736] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1737] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1738] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1739] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1740] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1741] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1742] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1743] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[1744] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[1745] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[1746] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1747] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1748] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1749] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1750] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1751] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1752] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1753] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1754] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1755] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1756] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1757] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1758] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1759] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1760] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1761] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1762] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1763] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1764] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1765] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1766] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1767] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1768] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1769] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1770] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1771] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1772] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1773] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1774] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1775] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1776] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1777] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1778] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1779] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1780] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1781] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1782] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1783] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1784] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1785] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1786] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1787] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1788] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1789] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1790] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1791] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[1792] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[1793] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[1794] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1795] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1796] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1797] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1798] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1799] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1800] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1801] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1802] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1803] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1804] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1805] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1806] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1807] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1808] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1809] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1810] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1811] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1812] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1813] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1814] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1815] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1816] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1817] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1818] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1819] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1820] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1821] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1822] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1823] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1824] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1825] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1826] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1827] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1828] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1829] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1830] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1831] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1832] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1833] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1834] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1835] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1836] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1837] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1838] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1839] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[1840] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[1841] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[1842] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1843] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1844] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1845] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1846] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1847] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1848] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1849] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1850] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1851] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1852] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1853] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1854] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1855] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1856] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1857] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1858] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1859] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1860] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1861] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1862] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1863] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1864] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1865] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1866] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1867] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1868] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1869] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1870] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1871] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1872] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1873] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1874] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1875] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1876] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1877] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1878] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1879] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1880] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1881] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1882] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1883] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1884] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1885] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1886] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1887] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[1888] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[1889] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[1890] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1891] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1892] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1893] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1894] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1895] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1896] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1897] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1898] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1899] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1900] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1901] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1902] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1903] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1904] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1905] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1906] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1907] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1908] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1909] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1910] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1911] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1912] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1913] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1914] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1915] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1916] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1917] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1918] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1919] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1920] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1921] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1922] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1923] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1924] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1925] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1926] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1927] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1928] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1929] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1930] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1931] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1932] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1933] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1934] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1935] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[1936] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[1937] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[1938] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1939] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1940] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1941] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1942] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1943] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1944] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1945] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1946] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1947] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1948] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1949] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1950] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1951] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1952] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1953] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1954] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1955] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1956] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1957] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1958] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1959] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1960] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1961] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1962] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1963] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1964] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1965] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1966] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1967] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1968] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1969] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1970] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1971] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1972] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1973] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1974] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1975] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1976] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1977] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1978] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1979] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1980] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1981] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1982] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1983] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[1984] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[1985] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[1986] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1987] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1988] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1989] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1990] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1991] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1992] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1993] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1994] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1995] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1996] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[1997] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[1998] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[1999] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2000] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2001] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2002] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2003] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2004] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2005] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2006] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2007] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2008] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2009] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2010] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2011] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2012] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2013] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2014] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2015] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2016] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2017] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2018] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2019] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2020] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2021] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2022] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2023] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2024] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2025] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2026] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2027] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2028] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2029] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2030] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2031] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[2032] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[2033] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[2034] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2035] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2036] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2037] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2038] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2039] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2040] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2041] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2042] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2043] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2044] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2045] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2046] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2047] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2048] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2049] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2050] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2051] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2052] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2053] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2054] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2055] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2056] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2057] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2058] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2059] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2060] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2061] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2062] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2063] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2064] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2065] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2066] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2067] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2068] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2069] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2070] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2071] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2072] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2073] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2074] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2075] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2076] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2077] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2078] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2079] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[2080] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[2081] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[2082] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2083] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2084] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2085] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2086] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2087] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2088] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2089] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2090] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2091] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2092] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2093] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2094] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2095] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2096] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2097] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2098] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2099] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2100] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2101] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2102] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2103] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2104] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2105] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2106] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2107] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2108] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2109] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2110] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2111] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2112] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2113] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2114] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2115] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2116] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2117] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2118] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2119] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2120] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2121] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2122] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2123] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2124] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2125] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2126] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2127] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[2128] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[2129] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[2130] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2131] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2132] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2133] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2134] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2135] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2136] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2137] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2138] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2139] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2140] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2141] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2142] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2143] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2144] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2145] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2146] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2147] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2148] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2149] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2150] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2151] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2152] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2153] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2154] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2155] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2156] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2157] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2158] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2159] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2160] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2161] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2162] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2163] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2164] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2165] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2166] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2167] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2168] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2169] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2170] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2171] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2172] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2173] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2174] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2175] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[2176] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[2177] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[2178] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2179] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2180] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2181] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2182] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2183] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2184] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2185] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2186] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2187] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2188] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2189] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2190] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2191] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2192] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2193] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2194] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2195] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2196] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2197] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2198] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2199] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2200] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2201] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2202] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2203] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2204] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2205] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2206] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2207] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2208] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2209] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2210] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2211] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2212] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2213] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2214] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2215] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2216] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2217] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2218] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2219] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2220] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2221] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2222] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2223] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[2224] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[2225] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[2226] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2227] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2228] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2229] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2230] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2231] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2232] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2233] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2234] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2235] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2236] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2237] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2238] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2239] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2240] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2241] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2242] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2243] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2244] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2245] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2246] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2247] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2248] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2249] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2250] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2251] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2252] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2253] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2254] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2255] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2256] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2257] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2258] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2259] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2260] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2261] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2262] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2263] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2264] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2265] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2266] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2267] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2268] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2269] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2270] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2271] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[2272] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[2273] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[2274] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2275] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2276] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2277] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2278] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2279] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2280] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2281] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2282] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2283] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2284] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2285] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2286] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2287] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2288] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2289] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2290] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2291] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2292] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2293] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2294] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2295] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2296] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2297] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2298] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2299] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2300] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2301] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2302] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2303] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2304] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2305] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2306] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2307] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2308] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2309] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2310] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2311] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2312] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2313] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2314] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2315] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2316] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[2317] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[2318] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[2319] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[2320] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[2321] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[2322] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2323] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2324] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2325] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2326] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2327] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2328] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2329] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2330] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2331] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2332] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2333] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2334] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2335] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2336] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2337] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2338] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2339] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2340] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2341] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2342] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2343] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2344] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2345] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2346] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2347] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2348] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2349] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2350] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2351] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2352] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2353] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2354] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2355] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2356] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2357] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2358] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2359] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2360] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2361] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2362] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2363] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2364] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2365] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2366] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2367] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[2368] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[2369] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[2370] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2371] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2372] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2373] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2374] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2375] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2376] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2377] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2378] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2379] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2380] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2381] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2382] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2383] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2384] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2385] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2386] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2387] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2388] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2389] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2390] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2391] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2392] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2393] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2394] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2395] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2396] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2397] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2398] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2399] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2400] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2401] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2402] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2403] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2404] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2405] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2406] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2407] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2408] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2409] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2410] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2411] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2412] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2413] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2414] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2415] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[2416] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[2417] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[2418] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2419] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2420] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2421] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2422] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2423] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2424] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2425] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2426] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2427] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2428] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2429] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2430] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2431] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2432] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2433] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2434] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2435] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2436] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2437] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2438] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2439] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2440] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2441] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2442] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2443] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2444] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2445] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2446] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2447] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2448] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2449] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2450] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2451] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2452] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2453] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2454] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2455] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2456] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2457] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2458] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2459] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2460] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2461] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2462] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2463] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[2464] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[2465] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[2466] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2467] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2468] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2469] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2470] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2471] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2472] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2473] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2474] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2475] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2476] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2477] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2478] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2479] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2480] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2481] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2482] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2483] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2484] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2485] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2486] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2487] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2488] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2489] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2490] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2491] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2492] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2493] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2494] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2495] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2496] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2497] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2498] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2499] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2500] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2501] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2502] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2503] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2504] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2505] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2506] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2507] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2508] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2509] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2510] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2511] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[2512] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[2513] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[2514] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2515] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2516] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2517] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2518] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2519] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2520] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2521] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2522] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2523] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2524] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2525] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2526] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2527] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2528] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2529] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2530] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2531] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2532] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2533] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2534] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2535] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2536] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2537] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2538] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2539] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2540] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2541] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2542] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2543] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2544] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2545] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2546] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2547] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2548] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2549] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2550] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2551] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2552] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2553] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2554] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2555] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2556] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2557] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2558] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2559] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[2560] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[2561] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[2562] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2563] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2564] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2565] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2566] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2567] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2568] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2569] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2570] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2571] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2572] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2573] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2574] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2575] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2576] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2577] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2578] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2579] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2580] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2581] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2582] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2583] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2584] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2585] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2586] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2587] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2588] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2589] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2590] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2591] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2592] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2593] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2594] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2595] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2596] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2597] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2598] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2599] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2600] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2601] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2602] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2603] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2604] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2605] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2606] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2607] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[2608] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[2609] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[2610] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2611] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2612] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2613] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2614] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2615] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2616] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2617] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2618] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2619] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2620] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2621] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2622] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2623] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2624] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2625] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2626] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2627] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2628] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2629] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2630] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2631] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2632] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2633] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2634] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2635] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2636] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2637] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2638] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2639] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2640] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2641] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2642] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2643] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2644] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2645] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2646] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2647] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2648] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2649] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2650] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2651] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2652] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2653] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2654] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2655] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[2656] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[2657] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[2658] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2659] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2660] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2661] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2662] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2663] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2664] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2665] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2666] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2667] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2668] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2669] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2670] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2671] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2672] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2673] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2674] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2675] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2676] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2677] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2678] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2679] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2680] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2681] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2682] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2683] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2684] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2685] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2686] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2687] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2688] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2689] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2690] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2691] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2692] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2693] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2694] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2695] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2696] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2697] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2698] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2699] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2700] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2701] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2702] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2703] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[2704] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[2705] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[2706] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2707] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2708] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2709] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2710] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2711] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2712] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2713] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2714] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2715] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2716] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2717] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2718] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2719] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2720] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2721] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2722] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2723] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2724] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2725] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2726] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2727] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2728] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2729] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2730] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2731] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2732] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2733] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2734] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2735] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2736] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2737] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2738] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2739] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2740] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2741] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2742] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2743] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2744] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2745] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2746] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2747] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2748] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2749] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2750] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2751] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[2752] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[2753] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[2754] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2755] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2756] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2757] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2758] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2759] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2760] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2761] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2762] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2763] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2764] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2765] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2766] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2767] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2768] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2769] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2770] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2771] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2772] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2773] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2774] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2775] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2776] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2777] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2778] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2779] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2780] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2781] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2782] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2783] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2784] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2785] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2786] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2787] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2788] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2789] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2790] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2791] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2792] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2793] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2794] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2795] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2796] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2797] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2798] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2799] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[2800] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[2801] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[2802] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2803] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2804] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2805] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2806] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2807] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2808] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2809] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2810] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2811] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2812] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2813] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2814] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2815] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2816] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2817] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2818] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2819] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2820] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2821] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2822] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2823] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2824] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2825] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2826] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2827] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2828] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2829] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2830] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2831] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2832] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2833] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2834] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2835] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2836] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2837] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2838] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2839] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2840] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2841] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2842] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2843] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2844] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2845] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2846] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2847] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[2848] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[2849] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[2850] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2851] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2852] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2853] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2854] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2855] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2856] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2857] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2858] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2859] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2860] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2861] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2862] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2863] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2864] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2865] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2866] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2867] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2868] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2869] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2870] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2871] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2872] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2873] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2874] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2875] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2876] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2877] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2878] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2879] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2880] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2881] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2882] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2883] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2884] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2885] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2886] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2887] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2888] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2889] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2890] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2891] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2892] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2893] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2894] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2895] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[2896] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[2897] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[2898] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2899] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2900] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2901] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2902] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2903] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2904] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2905] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2906] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2907] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2908] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2909] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2910] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2911] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2912] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2913] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2914] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2915] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2916] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2917] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2918] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2919] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2920] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2921] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2922] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2923] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2924] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2925] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2926] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2927] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2928] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2929] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2930] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2931] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2932] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2933] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2934] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2935] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2936] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2937] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2938] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2939] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2940] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2941] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2942] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2943] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[2944] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[2945] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[2946] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2947] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2948] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2949] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2950] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2951] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2952] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2953] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2954] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2955] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2956] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2957] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2958] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2959] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2960] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2961] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2962] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2963] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2964] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2965] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2966] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2967] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2968] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2969] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2970] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2971] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2972] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2973] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2974] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2975] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2976] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2977] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2978] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2979] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2980] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2981] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2982] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2983] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2984] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2985] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2986] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2987] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2988] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2989] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2990] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2991] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[2992] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[2993] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[2994] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2995] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2996] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[2997] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[2998] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[2999] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3000] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3001] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3002] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3003] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3004] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3005] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3006] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3007] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3008] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3009] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3010] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3011] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3012] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3013] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3014] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3015] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3016] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3017] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3018] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3019] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3020] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3021] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3022] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3023] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3024] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3025] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3026] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3027] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3028] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3029] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3030] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3031] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3032] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3033] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3034] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3035] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3036] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3037] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3038] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3039] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[3040] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[3041] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[3042] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3043] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3044] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3045] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3046] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3047] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3048] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3049] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3050] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3051] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3052] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3053] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3054] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3055] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3056] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3057] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3058] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3059] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3060] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3061] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3062] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3063] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3064] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3065] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3066] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3067] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3068] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3069] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3070] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3071] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3072] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3073] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3074] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3075] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3076] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3077] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3078] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3079] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3080] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3081] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3082] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3083] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3084] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3085] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3086] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3087] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[3088] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[3089] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[3090] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3091] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3092] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3093] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3094] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3095] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3096] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3097] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3098] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3099] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3100] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3101] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3102] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3103] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3104] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3105] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3106] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3107] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3108] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3109] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3110] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3111] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3112] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3113] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3114] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3115] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3116] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3117] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3118] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3119] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3120] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3121] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3122] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3123] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3124] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3125] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3126] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3127] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3128] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3129] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3130] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3131] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3132] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3133] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3134] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3135] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[3136] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[3137] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[3138] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3139] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3140] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3141] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3142] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3143] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3144] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3145] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3146] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3147] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3148] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3149] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3150] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3151] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3152] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3153] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3154] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3155] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3156] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3157] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3158] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3159] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3160] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3161] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3162] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3163] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3164] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3165] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3166] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3167] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3168] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3169] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3170] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3171] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3172] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3173] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3174] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3175] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3176] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3177] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3178] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3179] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3180] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3181] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3182] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3183] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[3184] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[3185] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[3186] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3187] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3188] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3189] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3190] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3191] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3192] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3193] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3194] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3195] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3196] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3197] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3198] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3199] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3200] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3201] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3202] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3203] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3204] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3205] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3206] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3207] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3208] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3209] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3210] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3211] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3212] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3213] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3214] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3215] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3216] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3217] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3218] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3219] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3220] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3221] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3222] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3223] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3224] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3225] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3226] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3227] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3228] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3229] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3230] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3231] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[3232] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[3233] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[3234] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3235] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3236] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3237] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3238] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3239] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3240] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3241] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3242] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3243] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3244] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3245] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3246] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3247] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3248] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3249] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3250] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3251] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3252] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3253] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3254] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3255] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3256] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3257] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3258] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3259] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3260] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3261] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3262] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3263] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3264] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3265] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3266] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3267] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3268] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3269] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3270] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3271] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3272] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3273] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3274] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3275] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3276] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3277] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3278] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3279] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[3280] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[3281] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[3282] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3283] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3284] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3285] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3286] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3287] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3288] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3289] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3290] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3291] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3292] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3293] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3294] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3295] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3296] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3297] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3298] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3299] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3300] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3301] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3302] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3303] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3304] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3305] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3306] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3307] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3308] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3309] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3310] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3311] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3312] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3313] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3314] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3315] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3316] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3317] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3318] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3319] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3320] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3321] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3322] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3323] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3324] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3325] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3326] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3327] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[3328] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[3329] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[3330] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3331] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3332] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3333] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3334] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3335] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3336] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3337] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3338] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3339] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3340] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3341] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3342] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3343] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3344] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3345] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3346] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3347] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3348] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3349] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3350] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3351] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3352] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3353] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3354] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3355] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3356] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3357] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3358] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3359] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3360] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3361] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3362] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3363] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3364] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3365] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3366] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3367] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3368] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3369] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3370] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3371] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3372] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3373] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3374] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3375] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[3376] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[3377] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[3378] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3379] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3380] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3381] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3382] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3383] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3384] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3385] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3386] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3387] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3388] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3389] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3390] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3391] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3392] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3393] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3394] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3395] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3396] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3397] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3398] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3399] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3400] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3401] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3402] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3403] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3404] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3405] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3406] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3407] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3408] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3409] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3410] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3411] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3412] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3413] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3414] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3415] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3416] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3417] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3418] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3419] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3420] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3421] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3422] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3423] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[3424] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[3425] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[3426] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3427] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3428] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3429] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3430] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3431] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3432] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3433] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3434] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3435] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3436] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3437] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3438] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3439] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3440] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3441] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3442] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3443] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3444] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3445] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3446] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3447] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3448] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3449] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3450] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3451] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3452] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3453] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3454] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3455] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3456] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3457] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3458] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3459] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3460] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3461] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3462] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3463] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3464] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3465] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3466] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3467] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3468] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3469] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3470] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3471] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[3472] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[3473] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[3474] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3475] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3476] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3477] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3478] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3479] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3480] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3481] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3482] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3483] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3484] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3485] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3486] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3487] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3488] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3489] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3490] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3491] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3492] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3493] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3494] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3495] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3496] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3497] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3498] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3499] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3500] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3501] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3502] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3503] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3504] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3505] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3506] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3507] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3508] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3509] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3510] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3511] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3512] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3513] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3514] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3515] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3516] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3517] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3518] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3519] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[3520] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[3521] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[3522] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3523] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3524] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3525] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3526] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3527] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3528] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3529] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3530] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3531] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3532] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3533] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3534] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3535] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3536] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3537] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3538] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3539] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3540] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3541] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3542] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3543] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3544] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3545] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3546] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3547] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3548] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3549] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3550] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3551] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3552] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3553] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3554] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3555] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3556] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3557] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3558] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3559] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3560] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3561] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3562] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3563] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3564] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3565] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3566] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3567] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[3568] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[3569] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[3570] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3571] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3572] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3573] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3574] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3575] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3576] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3577] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3578] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3579] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3580] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3581] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3582] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3583] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3584] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3585] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3586] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3587] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3588] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3589] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3590] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3591] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3592] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3593] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3594] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3595] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3596] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3597] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3598] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3599] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3600] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3601] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3602] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3603] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3604] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3605] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3606] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3607] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3608] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3609] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3610] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3611] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3612] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3613] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3614] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3615] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[3616] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[3617] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[3618] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3619] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3620] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3621] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3622] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3623] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3624] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3625] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3626] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3627] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3628] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3629] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3630] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3631] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3632] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3633] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3634] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3635] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3636] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3637] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3638] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3639] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3640] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3641] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3642] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3643] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3644] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3645] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3646] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3647] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3648] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3649] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3650] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3651] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3652] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3653] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3654] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3655] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3656] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3657] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3658] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3659] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3660] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3661] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3662] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3663] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[3664] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[3665] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[3666] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3667] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3668] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3669] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3670] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3671] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3672] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3673] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3674] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3675] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3676] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3677] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3678] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3679] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3680] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3681] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3682] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3683] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3684] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3685] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3686] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3687] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3688] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3689] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3690] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3691] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3692] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3693] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3694] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3695] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3696] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3697] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3698] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3699] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3700] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3701] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3702] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3703] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3704] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3705] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3706] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3707] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3708] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3709] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3710] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3711] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[3712] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[3713] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[3714] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3715] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3716] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3717] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3718] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3719] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3720] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3721] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3722] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3723] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3724] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3725] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3726] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3727] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3728] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3729] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3730] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3731] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3732] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3733] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3734] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3735] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3736] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3737] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3738] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3739] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3740] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3741] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3742] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3743] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3744] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3745] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3746] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3747] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3748] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3749] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3750] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3751] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3752] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3753] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3754] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3755] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3756] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3757] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3758] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3759] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[3760] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[3761] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[3762] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3763] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3764] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3765] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3766] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3767] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3768] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3769] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3770] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3771] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3772] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3773] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3774] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3775] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3776] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3777] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3778] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3779] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3780] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3781] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3782] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3783] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3784] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3785] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3786] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3787] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3788] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3789] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3790] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3791] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3792] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3793] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3794] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3795] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3796] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3797] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3798] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3799] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3800] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3801] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3802] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3803] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3804] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3805] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3806] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3807] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[3808] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[3809] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[3810] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3811] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3812] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3813] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3814] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3815] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3816] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3817] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3818] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3819] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3820] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3821] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3822] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3823] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3824] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3825] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3826] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3827] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3828] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3829] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3830] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3831] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3832] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3833] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3834] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3835] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3836] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3837] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3838] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3839] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3840] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3841] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3842] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3843] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3844] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3845] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3846] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3847] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3848] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3849] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3850] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3851] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3852] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[3853] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[3854] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[3855] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[3856] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[3857] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[3858] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3859] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3860] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3861] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3862] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3863] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3864] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3865] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3866] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3867] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3868] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3869] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3870] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3871] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3872] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3873] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3874] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3875] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3876] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3877] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3878] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3879] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3880] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3881] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3882] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3883] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3884] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3885] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3886] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3887] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3888] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3889] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3890] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3891] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3892] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3893] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3894] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3895] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3896] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3897] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3898] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3899] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3900] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3901] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3902] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3903] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[3904] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[3905] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[3906] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3907] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3908] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3909] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3910] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3911] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3912] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3913] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3914] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3915] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3916] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3917] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3918] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3919] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3920] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3921] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3922] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3923] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3924] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3925] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3926] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3927] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3928] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3929] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3930] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3931] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3932] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3933] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3934] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3935] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3936] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3937] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3938] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3939] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3940] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3941] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3942] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3943] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3944] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3945] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3946] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3947] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3948] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3949] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3950] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3951] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[3952] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[3953] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[3954] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3955] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3956] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3957] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3958] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3959] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3960] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3961] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3962] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3963] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3964] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3965] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3966] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3967] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3968] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3969] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3970] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3971] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3972] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3973] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3974] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3975] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3976] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3977] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3978] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3979] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3980] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3981] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3982] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3983] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3984] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3985] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3986] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3987] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3988] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3989] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3990] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3991] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3992] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3993] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3994] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3995] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3996] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[3997] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[3998] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[3999] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[4000] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[4001] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[4002] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4003] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4004] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4005] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4006] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4007] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4008] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4009] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4010] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4011] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4012] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4013] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4014] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4015] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4016] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4017] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4018] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4019] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4020] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4021] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4022] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4023] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4024] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4025] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4026] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4027] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4028] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4029] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4030] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4031] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4032] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4033] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4034] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4035] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4036] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4037] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4038] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4039] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4040] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4041] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4042] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4043] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4044] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4045] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4046] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4047] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[4048] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[4049] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[4050] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4051] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4052] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4053] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4054] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4055] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4056] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4057] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4058] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4059] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4060] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4061] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4062] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4063] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4064] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4065] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4066] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4067] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4068] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4069] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4070] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4071] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4072] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4073] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4074] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4075] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4076] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4077] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4078] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4079] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4080] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4081] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4082] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4083] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4084] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4085] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4086] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4087] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4088] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4089] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4090] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4091] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4092] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4093] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4094] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4095] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[4096] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[4097] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[4098] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4099] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4100] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4101] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4102] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4103] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4104] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4105] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4106] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4107] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4108] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4109] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4110] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4111] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4112] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4113] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4114] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4115] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4116] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4117] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4118] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4119] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4120] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4121] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4122] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4123] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4124] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4125] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4126] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4127] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4128] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4129] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4130] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4131] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4132] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4133] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4134] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4135] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4136] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4137] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4138] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4139] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4140] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4141] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4142] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4143] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[4144] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[4145] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[4146] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4147] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4148] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4149] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4150] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4151] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4152] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4153] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4154] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4155] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4156] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4157] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4158] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4159] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4160] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4161] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4162] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4163] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4164] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4165] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4166] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4167] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4168] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4169] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4170] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4171] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4172] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4173] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4174] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4175] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4176] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4177] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4178] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4179] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4180] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4181] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4182] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4183] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4184] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4185] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4186] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4187] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4188] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4189] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4190] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4191] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[4192] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[4193] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[4194] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4195] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4196] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4197] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4198] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4199] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4200] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4201] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4202] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4203] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4204] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4205] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4206] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4207] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4208] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4209] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4210] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4211] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4212] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4213] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4214] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4215] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4216] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4217] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4218] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4219] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4220] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4221] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4222] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4223] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4224] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4225] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4226] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4227] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4228] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4229] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4230] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4231] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4232] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4233] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4234] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4235] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4236] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4237] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4238] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4239] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[4240] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[4241] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[4242] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4243] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4244] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4245] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4246] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4247] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4248] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4249] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4250] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4251] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4252] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4253] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4254] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4255] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4256] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4257] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4258] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4259] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4260] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4261] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4262] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4263] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4264] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4265] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4266] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4267] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4268] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4269] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4270] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4271] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4272] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4273] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4274] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4275] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4276] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4277] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4278] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4279] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4280] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4281] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4282] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4283] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4284] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4285] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4286] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4287] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[4288] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[4289] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[4290] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4291] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4292] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4293] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4294] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4295] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4296] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4297] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4298] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4299] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4300] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4301] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4302] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4303] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4304] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4305] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4306] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4307] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4308] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4309] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4310] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4311] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4312] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4313] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4314] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4315] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4316] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4317] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4318] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4319] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4320] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4321] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4322] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4323] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4324] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4325] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4326] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4327] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4328] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4329] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4330] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4331] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4332] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4333] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4334] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4335] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[4336] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[4337] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[4338] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4339] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4340] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4341] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4342] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4343] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4344] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4345] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4346] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4347] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4348] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4349] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4350] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4351] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4352] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4353] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4354] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4355] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4356] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4357] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4358] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4359] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4360] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4361] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4362] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4363] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4364] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4365] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4366] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4367] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4368] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4369] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4370] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4371] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4372] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4373] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4374] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4375] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4376] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4377] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4378] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4379] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4380] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4381] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4382] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4383] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[4384] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[4385] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[4386] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4387] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4388] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4389] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4390] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4391] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4392] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4393] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4394] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4395] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4396] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4397] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4398] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4399] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4400] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4401] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4402] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4403] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4404] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4405] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4406] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4407] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4408] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4409] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4410] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4411] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4412] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4413] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4414] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4415] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4416] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4417] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4418] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4419] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4420] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4421] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4422] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4423] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4424] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4425] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4426] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4427] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4428] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4429] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4430] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4431] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[4432] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[4433] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[4434] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4435] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4436] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4437] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4438] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4439] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4440] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4441] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4442] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4443] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4444] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4445] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4446] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4447] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4448] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4449] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4450] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4451] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4452] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4453] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4454] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4455] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4456] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4457] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4458] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4459] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4460] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4461] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4462] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4463] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4464] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4465] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4466] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4467] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4468] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4469] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4470] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4471] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4472] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4473] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4474] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4475] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4476] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4477] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4478] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4479] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[4480] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[4481] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[4482] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4483] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4484] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4485] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4486] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4487] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4488] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4489] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4490] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4491] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4492] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4493] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4494] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4495] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4496] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4497] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4498] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4499] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4500] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4501] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4502] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4503] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4504] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4505] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4506] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4507] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4508] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4509] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4510] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4511] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4512] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4513] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4514] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4515] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4516] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4517] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4518] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4519] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4520] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4521] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4522] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4523] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4524] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4525] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4526] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4527] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[4528] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[4529] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[4530] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4531] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4532] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4533] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4534] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4535] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4536] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4537] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4538] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4539] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4540] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4541] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4542] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4543] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4544] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4545] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4546] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4547] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4548] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4549] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4550] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4551] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4552] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4553] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4554] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4555] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4556] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4557] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4558] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4559] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4560] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4561] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4562] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4563] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4564] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4565] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4566] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4567] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4568] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4569] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4570] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4571] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4572] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4573] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4574] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4575] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[4576] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[4577] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[4578] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4579] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4580] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4581] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4582] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4583] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4584] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4585] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4586] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4587] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4588] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4589] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4590] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4591] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4592] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4593] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4594] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4595] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4596] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4597] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4598] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4599] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4600] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4601] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4602] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4603] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4604] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4605] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4606] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4607] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4608] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4609] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4610] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4611] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4612] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4613] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4614] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4615] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4616] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4617] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4618] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4619] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4620] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[4621] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[4622] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[4623] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[4624] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[4625] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[4626] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4627] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4628] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4629] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4630] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4631] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4632] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4633] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4634] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4635] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4636] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4637] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4638] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4639] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4640] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4641] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4642] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4643] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4644] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4645] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4646] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4647] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4648] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4649] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4650] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4651] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4652] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4653] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4654] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4655] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4656] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4657] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4658] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4659] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4660] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4661] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4662] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4663] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4664] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4665] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4666] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4667] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4668] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4669] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4670] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4671] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[4672] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[4673] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[4674] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4675] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4676] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4677] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4678] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4679] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4680] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4681] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4682] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4683] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4684] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4685] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4686] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4687] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4688] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4689] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4690] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4691] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4692] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4693] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4694] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4695] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4696] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4697] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4698] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4699] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4700] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4701] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4702] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4703] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4704] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4705] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4706] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4707] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4708] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4709] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4710] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4711] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4712] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4713] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4714] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4715] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4716] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4717] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4718] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4719] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[4720] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[4721] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[4722] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4723] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4724] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4725] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4726] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4727] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4728] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4729] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4730] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4731] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4732] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4733] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4734] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4735] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4736] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4737] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4738] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4739] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4740] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4741] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4742] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4743] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4744] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4745] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4746] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4747] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4748] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4749] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4750] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4751] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4752] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4753] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4754] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4755] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4756] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4757] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4758] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4759] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4760] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4761] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4762] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4763] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4764] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4765] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4766] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4767] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[4768] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[4769] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[4770] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4771] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4772] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4773] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4774] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4775] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4776] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4777] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4778] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4779] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4780] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4781] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4782] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4783] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4784] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4785] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4786] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4787] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4788] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4789] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4790] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4791] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4792] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4793] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4794] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4795] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4796] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4797] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4798] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4799] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4800] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4801] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4802] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4803] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4804] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4805] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4806] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4807] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4808] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4809] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4810] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4811] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4812] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4813] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4814] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4815] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[4816] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[4817] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[4818] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4819] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4820] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4821] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4822] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4823] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4824] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4825] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4826] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4827] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4828] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4829] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4830] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4831] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4832] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4833] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4834] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4835] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4836] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4837] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4838] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4839] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4840] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4841] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4842] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4843] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4844] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4845] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4846] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4847] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4848] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4849] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4850] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4851] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4852] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4853] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4854] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4855] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4856] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4857] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4858] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4859] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4860] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4861] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4862] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4863] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[4864] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[4865] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[4866] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4867] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4868] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4869] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4870] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4871] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4872] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4873] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4874] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4875] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4876] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4877] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4878] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4879] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4880] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4881] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4882] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4883] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4884] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4885] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4886] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4887] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4888] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4889] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4890] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4891] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4892] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4893] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4894] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4895] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4896] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4897] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4898] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4899] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4900] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4901] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4902] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4903] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4904] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4905] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4906] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4907] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4908] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4909] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4910] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4911] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[4912] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[4913] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[4914] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4915] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4916] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4917] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4918] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4919] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4920] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4921] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4922] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4923] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4924] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4925] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4926] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4927] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4928] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4929] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4930] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4931] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4932] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4933] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4934] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4935] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4936] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4937] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4938] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4939] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4940] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4941] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4942] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4943] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4944] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4945] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4946] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4947] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4948] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4949] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4950] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4951] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4952] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4953] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4954] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4955] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4956] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4957] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4958] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4959] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[4960] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[4961] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[4962] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4963] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4964] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4965] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4966] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4967] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4968] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4969] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4970] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4971] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4972] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4973] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4974] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4975] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4976] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4977] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4978] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4979] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4980] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4981] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4982] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4983] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4984] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4985] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4986] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4987] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4988] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4989] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4990] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4991] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4992] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4993] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4994] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4995] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4996] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[4997] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[4998] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[4999] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5000] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5001] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5002] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5003] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5004] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5005] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5006] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5007] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[5008] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[5009] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[5010] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5011] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5012] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5013] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5014] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5015] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5016] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5017] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5018] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5019] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5020] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5021] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5022] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5023] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5024] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5025] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5026] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5027] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5028] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5029] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5030] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5031] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5032] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5033] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5034] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5035] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5036] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5037] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5038] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5039] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5040] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5041] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5042] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5043] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5044] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5045] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5046] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5047] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5048] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5049] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5050] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5051] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5052] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5053] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5054] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5055] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[5056] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[5057] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[5058] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5059] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5060] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5061] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5062] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5063] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5064] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5065] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5066] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5067] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5068] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5069] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5070] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5071] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5072] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5073] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5074] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5075] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5076] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5077] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5078] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5079] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5080] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5081] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5082] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5083] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5084] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5085] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5086] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5087] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5088] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5089] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5090] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5091] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5092] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5093] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5094] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5095] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5096] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5097] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5098] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5099] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5100] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5101] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5102] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5103] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[5104] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[5105] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[5106] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5107] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5108] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5109] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5110] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5111] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5112] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5113] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5114] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5115] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5116] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5117] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5118] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5119] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5120] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5121] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5122] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5123] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5124] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5125] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5126] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5127] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5128] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5129] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5130] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5131] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5132] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5133] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5134] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5135] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5136] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5137] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5138] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5139] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5140] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5141] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5142] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5143] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5144] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5145] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5146] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5147] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5148] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5149] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5150] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5151] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[5152] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[5153] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[5154] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5155] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5156] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5157] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5158] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5159] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5160] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5161] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5162] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5163] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5164] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5165] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5166] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5167] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5168] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5169] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5170] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5171] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5172] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5173] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5174] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5175] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5176] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5177] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5178] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5179] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5180] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5181] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5182] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5183] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5184] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5185] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5186] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5187] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5188] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5189] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5190] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5191] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5192] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5193] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5194] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5195] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5196] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5197] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5198] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5199] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[5200] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[5201] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[5202] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5203] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5204] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5205] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5206] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5207] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5208] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5209] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5210] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5211] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5212] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5213] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5214] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5215] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5216] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5217] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5218] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5219] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5220] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5221] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5222] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5223] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5224] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5225] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5226] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5227] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5228] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5229] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5230] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5231] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5232] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5233] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5234] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5235] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5236] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5237] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5238] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5239] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5240] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5241] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5242] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5243] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5244] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5245] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5246] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5247] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[5248] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[5249] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[5250] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5251] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5252] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5253] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5254] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5255] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5256] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5257] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5258] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5259] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5260] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5261] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5262] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5263] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5264] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5265] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5266] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5267] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5268] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5269] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5270] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5271] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5272] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5273] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5274] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5275] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5276] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5277] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5278] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5279] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5280] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5281] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5282] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5283] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5284] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5285] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5286] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5287] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5288] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5289] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5290] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5291] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5292] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5293] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5294] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5295] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[5296] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[5297] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[5298] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5299] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5300] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5301] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5302] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5303] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5304] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5305] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5306] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5307] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5308] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5309] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5310] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5311] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5312] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5313] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5314] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5315] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5316] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5317] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5318] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5319] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5320] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5321] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5322] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5323] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5324] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5325] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5326] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5327] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5328] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5329] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5330] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5331] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5332] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5333] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5334] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5335] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5336] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5337] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5338] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5339] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5340] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5341] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5342] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5343] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[5344] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[5345] = 13'b1_0_0_1_xxxxxxxx_0;
      patterns[5346] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5347] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5348] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5349] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5350] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5351] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5352] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5353] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5354] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5355] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5356] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5357] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5358] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5359] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5360] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5361] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5362] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5363] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5364] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5365] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5366] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5367] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5368] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5369] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5370] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5371] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5372] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5373] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5374] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5375] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5376] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5377] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5378] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5379] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5380] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5381] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5382] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5383] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5384] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5385] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5386] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5387] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5388] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[5389] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[5390] = 13'b0_0_0_1_xxxxxxxx_0;
      patterns[5391] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[5392] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[5393] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[5394] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5395] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5396] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5397] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5398] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5399] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5400] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5401] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5402] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5403] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5404] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5405] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5406] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5407] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5408] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5409] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5410] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5411] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5412] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5413] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5414] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5415] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5416] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5417] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5418] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5419] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5420] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5421] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5422] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5423] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5424] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5425] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5426] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5427] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5428] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5429] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5430] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5431] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5432] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5433] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5434] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5435] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5436] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5437] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5438] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5439] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[5440] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[5441] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[5442] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5443] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5444] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5445] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5446] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5447] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5448] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5449] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5450] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5451] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5452] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5453] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5454] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5455] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5456] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5457] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5458] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5459] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5460] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5461] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5462] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5463] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5464] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5465] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5466] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5467] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5468] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5469] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5470] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5471] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5472] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5473] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5474] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5475] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5476] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5477] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5478] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5479] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5480] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5481] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5482] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5483] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5484] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5485] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5486] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5487] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[5488] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[5489] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[5490] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5491] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5492] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5493] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5494] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5495] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5496] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5497] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5498] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5499] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5500] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5501] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5502] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5503] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5504] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5505] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5506] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5507] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5508] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5509] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5510] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5511] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5512] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5513] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5514] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5515] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5516] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5517] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5518] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5519] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5520] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5521] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5522] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5523] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5524] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5525] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5526] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5527] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5528] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5529] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5530] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5531] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5532] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5533] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5534] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5535] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[5536] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[5537] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[5538] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5539] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5540] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5541] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5542] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5543] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5544] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5545] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5546] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5547] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5548] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5549] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5550] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5551] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5552] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5553] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5554] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5555] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5556] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5557] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5558] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5559] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5560] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5561] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5562] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5563] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5564] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5565] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5566] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5567] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5568] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5569] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5570] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5571] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5572] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5573] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5574] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5575] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5576] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5577] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5578] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5579] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5580] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5581] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5582] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5583] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[5584] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[5585] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[5586] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5587] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5588] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5589] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5590] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5591] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5592] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5593] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5594] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5595] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5596] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5597] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5598] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5599] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5600] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5601] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5602] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5603] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5604] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5605] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5606] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5607] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5608] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5609] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5610] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5611] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5612] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5613] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5614] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5615] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5616] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5617] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5618] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5619] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5620] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5621] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5622] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5623] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5624] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5625] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5626] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5627] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5628] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5629] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5630] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5631] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[5632] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[5633] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[5634] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5635] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5636] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5637] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5638] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5639] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5640] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5641] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5642] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5643] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5644] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5645] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5646] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5647] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5648] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5649] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5650] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5651] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5652] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5653] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5654] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5655] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5656] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5657] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5658] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5659] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5660] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5661] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5662] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5663] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5664] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5665] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5666] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5667] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5668] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5669] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5670] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5671] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5672] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5673] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5674] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5675] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5676] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5677] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5678] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5679] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[5680] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[5681] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[5682] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5683] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5684] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5685] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5686] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5687] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5688] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5689] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5690] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5691] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5692] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5693] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5694] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5695] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5696] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5697] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5698] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5699] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5700] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5701] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5702] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5703] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5704] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5705] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5706] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5707] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5708] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5709] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5710] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5711] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5712] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5713] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5714] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5715] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5716] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5717] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5718] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5719] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5720] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5721] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5722] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5723] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5724] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5725] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5726] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5727] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[5728] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[5729] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[5730] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5731] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5732] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5733] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5734] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5735] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5736] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5737] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5738] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5739] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5740] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5741] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5742] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5743] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5744] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5745] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5746] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5747] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5748] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5749] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5750] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5751] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5752] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5753] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5754] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5755] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5756] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5757] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5758] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5759] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5760] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5761] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5762] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5763] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5764] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5765] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5766] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5767] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5768] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5769] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5770] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5771] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5772] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5773] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5774] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5775] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[5776] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[5777] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[5778] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5779] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5780] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5781] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5782] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5783] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5784] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5785] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5786] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5787] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5788] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5789] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5790] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5791] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5792] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5793] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5794] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5795] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5796] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5797] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5798] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5799] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5800] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5801] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5802] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5803] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5804] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5805] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5806] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5807] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5808] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5809] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5810] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5811] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5812] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5813] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5814] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5815] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5816] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5817] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5818] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5819] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5820] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5821] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5822] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5823] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[5824] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[5825] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[5826] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5827] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5828] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5829] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5830] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5831] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5832] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5833] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5834] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5835] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5836] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5837] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5838] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5839] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5840] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5841] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5842] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5843] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5844] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5845] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5846] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5847] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5848] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5849] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5850] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5851] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5852] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5853] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5854] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5855] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5856] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5857] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5858] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5859] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5860] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5861] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5862] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5863] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5864] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5865] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5866] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5867] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5868] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5869] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5870] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5871] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[5872] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[5873] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[5874] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5875] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5876] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5877] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5878] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5879] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5880] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5881] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5882] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5883] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5884] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5885] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5886] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5887] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5888] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5889] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5890] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5891] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5892] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5893] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5894] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5895] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5896] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5897] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5898] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5899] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5900] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5901] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5902] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5903] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5904] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5905] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5906] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5907] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5908] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5909] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5910] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5911] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5912] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5913] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5914] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5915] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5916] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5917] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5918] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5919] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[5920] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[5921] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[5922] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5923] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5924] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5925] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5926] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5927] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5928] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5929] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5930] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5931] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5932] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5933] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5934] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5935] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5936] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5937] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5938] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5939] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5940] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5941] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5942] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5943] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5944] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5945] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5946] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5947] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5948] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5949] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5950] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5951] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5952] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5953] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5954] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5955] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5956] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5957] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5958] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5959] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5960] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5961] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5962] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5963] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5964] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5965] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5966] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5967] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[5968] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[5969] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[5970] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5971] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5972] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5973] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5974] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5975] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5976] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5977] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5978] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5979] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5980] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5981] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5982] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5983] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5984] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5985] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5986] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5987] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5988] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5989] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5990] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5991] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5992] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5993] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5994] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5995] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5996] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[5997] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[5998] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[5999] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6000] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6001] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6002] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6003] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6004] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6005] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6006] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6007] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6008] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6009] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6010] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6011] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6012] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6013] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6014] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6015] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[6016] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[6017] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[6018] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6019] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6020] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6021] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6022] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6023] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6024] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6025] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6026] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6027] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6028] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6029] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6030] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6031] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6032] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6033] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6034] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6035] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6036] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6037] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6038] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6039] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6040] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6041] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6042] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6043] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6044] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6045] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6046] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6047] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6048] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6049] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6050] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6051] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6052] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6053] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6054] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6055] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6056] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6057] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6058] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6059] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6060] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6061] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6062] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6063] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[6064] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[6065] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[6066] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6067] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6068] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6069] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6070] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6071] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6072] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6073] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6074] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6075] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6076] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6077] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6078] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6079] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6080] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6081] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6082] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6083] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6084] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6085] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6086] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6087] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6088] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6089] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6090] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6091] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6092] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6093] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6094] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6095] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6096] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6097] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6098] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6099] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6100] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6101] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6102] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6103] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6104] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6105] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6106] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6107] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6108] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6109] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6110] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6111] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[6112] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[6113] = 13'b1_0_0_0_xxxxxxxx_0;
      patterns[6114] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6115] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6116] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6117] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6118] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6119] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6120] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6121] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6122] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6123] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6124] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6125] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6126] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6127] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6128] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6129] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6130] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6131] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6132] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6133] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6134] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6135] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6136] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6137] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6138] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6139] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6140] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6141] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6142] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6143] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6144] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6145] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6146] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6147] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6148] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6149] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6150] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6151] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6152] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6153] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6154] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6155] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6156] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6157] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6158] = 13'b0_0_0_0_xxxxxxxx_0;
      patterns[6159] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[6160] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[6161] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[6162] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6163] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6164] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6165] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6166] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6167] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6168] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6169] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6170] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6171] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6172] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6173] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6174] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6175] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6176] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6177] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6178] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6179] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6180] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6181] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6182] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6183] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6184] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6185] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6186] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6187] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6188] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6189] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6190] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6191] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6192] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6193] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6194] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6195] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6196] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6197] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6198] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6199] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6200] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6201] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6202] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6203] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6204] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6205] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6206] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6207] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[6208] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[6209] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[6210] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6211] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6212] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6213] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6214] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6215] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6216] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6217] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6218] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6219] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6220] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6221] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6222] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6223] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6224] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6225] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6226] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6227] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6228] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6229] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6230] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6231] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6232] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6233] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6234] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6235] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6236] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6237] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6238] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6239] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6240] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6241] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6242] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6243] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6244] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6245] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6246] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6247] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6248] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6249] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6250] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6251] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6252] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6253] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6254] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6255] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[6256] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[6257] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[6258] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6259] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6260] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6261] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6262] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6263] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6264] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6265] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6266] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6267] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6268] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6269] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6270] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6271] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6272] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6273] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6274] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6275] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6276] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6277] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6278] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6279] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6280] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6281] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6282] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6283] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6284] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6285] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6286] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6287] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6288] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6289] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6290] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6291] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6292] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6293] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6294] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6295] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6296] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6297] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6298] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6299] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6300] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6301] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6302] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6303] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[6304] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[6305] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[6306] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6307] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6308] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6309] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6310] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6311] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6312] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6313] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6314] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6315] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6316] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6317] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6318] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6319] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6320] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6321] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6322] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6323] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6324] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6325] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6326] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6327] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6328] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6329] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6330] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6331] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6332] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6333] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6334] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6335] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6336] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6337] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6338] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6339] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6340] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6341] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6342] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6343] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6344] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6345] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6346] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6347] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6348] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6349] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6350] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6351] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[6352] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[6353] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[6354] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6355] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6356] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6357] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6358] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6359] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6360] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6361] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6362] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6363] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6364] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6365] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6366] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6367] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6368] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6369] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6370] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6371] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6372] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6373] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6374] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6375] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6376] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6377] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6378] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6379] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6380] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6381] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6382] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6383] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6384] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6385] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6386] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6387] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6388] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6389] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6390] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6391] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6392] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6393] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6394] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6395] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6396] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6397] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6398] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6399] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[6400] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[6401] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[6402] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6403] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6404] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6405] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6406] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6407] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6408] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6409] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6410] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6411] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6412] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6413] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6414] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6415] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6416] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6417] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6418] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6419] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6420] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6421] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6422] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6423] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6424] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6425] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6426] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6427] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6428] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6429] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6430] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6431] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6432] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6433] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6434] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6435] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6436] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6437] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6438] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6439] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6440] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6441] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6442] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6443] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6444] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6445] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6446] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6447] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[6448] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[6449] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[6450] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6451] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6452] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6453] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6454] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6455] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6456] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6457] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6458] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6459] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6460] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6461] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6462] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6463] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6464] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6465] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6466] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6467] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6468] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6469] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6470] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6471] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6472] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6473] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6474] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6475] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6476] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6477] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6478] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6479] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6480] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6481] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6482] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6483] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6484] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6485] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6486] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6487] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6488] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6489] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6490] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6491] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6492] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6493] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6494] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6495] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[6496] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[6497] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[6498] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6499] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6500] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6501] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6502] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6503] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6504] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6505] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6506] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6507] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6508] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6509] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6510] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6511] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6512] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6513] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6514] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6515] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6516] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6517] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6518] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6519] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6520] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6521] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6522] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6523] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6524] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6525] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6526] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6527] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6528] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6529] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6530] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6531] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6532] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6533] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6534] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6535] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6536] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6537] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6538] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6539] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6540] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6541] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6542] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6543] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[6544] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[6545] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[6546] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6547] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6548] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6549] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6550] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6551] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6552] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6553] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6554] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6555] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6556] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6557] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6558] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6559] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6560] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6561] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6562] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6563] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6564] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6565] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6566] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6567] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6568] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6569] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6570] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6571] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6572] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6573] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6574] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6575] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6576] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6577] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6578] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6579] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6580] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6581] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6582] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6583] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6584] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6585] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6586] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6587] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6588] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6589] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6590] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6591] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[6592] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[6593] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[6594] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6595] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6596] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6597] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6598] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6599] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6600] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6601] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6602] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6603] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6604] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6605] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6606] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6607] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6608] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6609] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6610] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6611] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6612] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6613] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6614] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6615] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6616] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6617] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6618] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6619] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6620] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6621] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6622] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6623] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6624] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6625] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6626] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6627] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6628] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6629] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6630] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6631] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6632] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6633] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6634] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6635] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6636] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6637] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6638] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6639] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[6640] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[6641] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[6642] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6643] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6644] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6645] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6646] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6647] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6648] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6649] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6650] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6651] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6652] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6653] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6654] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6655] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6656] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6657] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6658] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6659] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6660] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6661] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6662] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6663] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6664] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6665] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6666] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6667] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6668] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6669] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6670] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6671] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6672] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6673] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6674] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6675] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6676] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6677] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6678] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6679] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6680] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6681] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6682] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6683] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6684] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6685] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6686] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6687] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[6688] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[6689] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[6690] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6691] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6692] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6693] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6694] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6695] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6696] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6697] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6698] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6699] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6700] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6701] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6702] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6703] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6704] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6705] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6706] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6707] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6708] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6709] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6710] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6711] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6712] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6713] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6714] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6715] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6716] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6717] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6718] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6719] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6720] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6721] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6722] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6723] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6724] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6725] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6726] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6727] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6728] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6729] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6730] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6731] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6732] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6733] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6734] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6735] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[6736] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[6737] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[6738] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6739] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6740] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6741] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6742] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6743] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6744] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6745] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6746] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6747] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6748] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6749] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6750] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6751] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6752] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6753] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6754] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6755] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6756] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6757] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6758] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6759] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6760] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6761] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6762] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6763] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6764] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6765] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6766] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6767] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6768] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6769] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6770] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6771] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6772] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6773] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6774] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6775] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6776] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6777] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6778] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6779] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6780] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6781] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6782] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6783] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[6784] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[6785] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[6786] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6787] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6788] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6789] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6790] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6791] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6792] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6793] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6794] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6795] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6796] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6797] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6798] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6799] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6800] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6801] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6802] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6803] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6804] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6805] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6806] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6807] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6808] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6809] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6810] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6811] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6812] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6813] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6814] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6815] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6816] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6817] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6818] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6819] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6820] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6821] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6822] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6823] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6824] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6825] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6826] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6827] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6828] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6829] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6830] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6831] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[6832] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[6833] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[6834] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6835] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6836] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6837] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6838] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6839] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6840] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6841] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6842] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6843] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6844] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6845] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6846] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6847] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6848] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6849] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6850] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6851] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6852] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6853] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6854] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6855] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6856] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6857] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6858] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6859] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6860] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6861] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6862] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6863] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6864] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6865] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6866] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6867] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6868] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6869] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6870] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6871] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6872] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6873] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6874] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6875] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6876] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6877] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6878] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6879] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[6880] = 13'b1_0_1_1_xxxxxxxx_x;
      patterns[6881] = 13'b1_0_0_1_xxxxxxxx_x;
      patterns[6882] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6883] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6884] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6885] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6886] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6887] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6888] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6889] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6890] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6891] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6892] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6893] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6894] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6895] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6896] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6897] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6898] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6899] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6900] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6901] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6902] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6903] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6904] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6905] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6906] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6907] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6908] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6909] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6910] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6911] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6912] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6913] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6914] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6915] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6916] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6917] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6918] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6919] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6920] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6921] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6922] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6923] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6924] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6925] = 13'b0_0_1_1_xxxxxxxx_x;
      patterns[6926] = 13'b0_0_0_1_xxxxxxxx_x;
      patterns[6927] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[6928] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[6929] = 13'b1_0_0_0_10101010_1;
      patterns[6930] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6931] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6932] = 13'b0_0_0_0_10101010_1;
      patterns[6933] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6934] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6935] = 13'b0_0_0_0_10101010_1;
      patterns[6936] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6937] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6938] = 13'b0_0_0_0_10101010_1;
      patterns[6939] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6940] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6941] = 13'b0_0_0_0_10101010_1;
      patterns[6942] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6943] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6944] = 13'b0_0_0_0_10101010_1;
      patterns[6945] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6946] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6947] = 13'b0_0_0_0_10101010_1;
      patterns[6948] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6949] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6950] = 13'b0_0_0_0_10101010_1;
      patterns[6951] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6952] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6953] = 13'b0_0_0_0_10101010_1;
      patterns[6954] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6955] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6956] = 13'b0_0_0_0_10101010_1;
      patterns[6957] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6958] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6959] = 13'b0_0_0_0_10101010_1;
      patterns[6960] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6961] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6962] = 13'b0_0_0_0_10101010_1;
      patterns[6963] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6964] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6965] = 13'b0_0_0_0_10101010_1;
      patterns[6966] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6967] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6968] = 13'b0_0_0_0_10101010_1;
      patterns[6969] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6970] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6971] = 13'b0_0_0_0_10101010_1;
      patterns[6972] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6973] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6974] = 13'b0_0_0_0_10101010_1;
      patterns[6975] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[6976] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[6977] = 13'b1_0_0_0_10101010_1;
      patterns[6978] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6979] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6980] = 13'b0_0_0_0_10101010_1;
      patterns[6981] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6982] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6983] = 13'b0_0_0_0_10101010_1;
      patterns[6984] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6985] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6986] = 13'b0_0_0_0_10101010_1;
      patterns[6987] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6988] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6989] = 13'b0_0_0_0_10101010_1;
      patterns[6990] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6991] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6992] = 13'b0_0_0_0_10101010_1;
      patterns[6993] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6994] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6995] = 13'b0_0_0_0_10101010_1;
      patterns[6996] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[6997] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[6998] = 13'b0_0_0_0_10101010_1;
      patterns[6999] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7000] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7001] = 13'b0_0_0_0_10101010_1;
      patterns[7002] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7003] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7004] = 13'b0_0_0_0_10101010_1;
      patterns[7005] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7006] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7007] = 13'b0_0_0_0_10101010_1;
      patterns[7008] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7009] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7010] = 13'b0_0_0_0_10101010_1;
      patterns[7011] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7012] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7013] = 13'b0_0_0_0_10101010_1;
      patterns[7014] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7015] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7016] = 13'b0_0_0_0_10101010_1;
      patterns[7017] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7018] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7019] = 13'b0_0_0_0_10101010_1;
      patterns[7020] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7021] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7022] = 13'b0_0_0_0_10101010_1;
      patterns[7023] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[7024] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[7025] = 13'b1_0_0_0_10101010_1;
      patterns[7026] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7027] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7028] = 13'b0_0_0_0_10101010_1;
      patterns[7029] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7030] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7031] = 13'b0_0_0_0_10101010_1;
      patterns[7032] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7033] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7034] = 13'b0_0_0_0_10101010_1;
      patterns[7035] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7036] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7037] = 13'b0_0_0_0_10101010_1;
      patterns[7038] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7039] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7040] = 13'b0_0_0_0_10101010_1;
      patterns[7041] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7042] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7043] = 13'b0_0_0_0_10101010_1;
      patterns[7044] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7045] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7046] = 13'b0_0_0_0_10101010_1;
      patterns[7047] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7048] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7049] = 13'b0_0_0_0_10101010_1;
      patterns[7050] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7051] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7052] = 13'b0_0_0_0_10101010_1;
      patterns[7053] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7054] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7055] = 13'b0_0_0_0_10101010_1;
      patterns[7056] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7057] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7058] = 13'b0_0_0_0_10101010_1;
      patterns[7059] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7060] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7061] = 13'b0_0_0_0_10101010_1;
      patterns[7062] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7063] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7064] = 13'b0_0_0_0_10101010_1;
      patterns[7065] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7066] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7067] = 13'b0_0_0_0_10101010_1;
      patterns[7068] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7069] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7070] = 13'b0_0_0_0_10101010_1;
      patterns[7071] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[7072] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[7073] = 13'b1_0_0_0_10101010_1;
      patterns[7074] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7075] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7076] = 13'b0_0_0_0_10101010_1;
      patterns[7077] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7078] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7079] = 13'b0_0_0_0_10101010_1;
      patterns[7080] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7081] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7082] = 13'b0_0_0_0_10101010_1;
      patterns[7083] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7084] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7085] = 13'b0_0_0_0_10101010_1;
      patterns[7086] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7087] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7088] = 13'b0_0_0_0_10101010_1;
      patterns[7089] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7090] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7091] = 13'b0_0_0_0_10101010_1;
      patterns[7092] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7093] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7094] = 13'b0_0_0_0_10101010_1;
      patterns[7095] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7096] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7097] = 13'b0_0_0_0_10101010_1;
      patterns[7098] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7099] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7100] = 13'b0_0_0_0_10101010_1;
      patterns[7101] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7102] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7103] = 13'b0_0_0_0_10101010_1;
      patterns[7104] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7105] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7106] = 13'b0_0_0_0_10101010_1;
      patterns[7107] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7108] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7109] = 13'b0_0_0_0_10101010_1;
      patterns[7110] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7111] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7112] = 13'b0_0_0_0_10101010_1;
      patterns[7113] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7114] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7115] = 13'b0_0_0_0_10101010_1;
      patterns[7116] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7117] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7118] = 13'b0_0_0_0_10101010_1;
      patterns[7119] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[7120] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[7121] = 13'b1_0_0_0_10101010_1;
      patterns[7122] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7123] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7124] = 13'b0_0_0_0_10101010_1;
      patterns[7125] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7126] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7127] = 13'b0_0_0_0_10101010_1;
      patterns[7128] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7129] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7130] = 13'b0_0_0_0_10101010_1;
      patterns[7131] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7132] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7133] = 13'b0_0_0_0_10101010_1;
      patterns[7134] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7135] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7136] = 13'b0_0_0_0_10101010_1;
      patterns[7137] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7138] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7139] = 13'b0_0_0_0_10101010_1;
      patterns[7140] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7141] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7142] = 13'b0_0_0_0_10101010_1;
      patterns[7143] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7144] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7145] = 13'b0_0_0_0_10101010_1;
      patterns[7146] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7147] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7148] = 13'b0_0_0_0_10101010_1;
      patterns[7149] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7150] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7151] = 13'b0_0_0_0_10101010_1;
      patterns[7152] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7153] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7154] = 13'b0_0_0_0_10101010_1;
      patterns[7155] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7156] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7157] = 13'b0_0_0_0_10101010_1;
      patterns[7158] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7159] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7160] = 13'b0_0_0_0_10101010_1;
      patterns[7161] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7162] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7163] = 13'b0_0_0_0_10101010_1;
      patterns[7164] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7165] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7166] = 13'b0_0_0_0_10101010_1;
      patterns[7167] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[7168] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[7169] = 13'b1_0_0_0_10101010_1;
      patterns[7170] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7171] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7172] = 13'b0_0_0_0_10101010_1;
      patterns[7173] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7174] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7175] = 13'b0_0_0_0_10101010_1;
      patterns[7176] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7177] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7178] = 13'b0_0_0_0_10101010_1;
      patterns[7179] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7180] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7181] = 13'b0_0_0_0_10101010_1;
      patterns[7182] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7183] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7184] = 13'b0_0_0_0_10101010_1;
      patterns[7185] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7186] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7187] = 13'b0_0_0_0_10101010_1;
      patterns[7188] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7189] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7190] = 13'b0_0_0_0_10101010_1;
      patterns[7191] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7192] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7193] = 13'b0_0_0_0_10101010_1;
      patterns[7194] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7195] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7196] = 13'b0_0_0_0_10101010_1;
      patterns[7197] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7198] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7199] = 13'b0_0_0_0_10101010_1;
      patterns[7200] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7201] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7202] = 13'b0_0_0_0_10101010_1;
      patterns[7203] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7204] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7205] = 13'b0_0_0_0_10101010_1;
      patterns[7206] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7207] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7208] = 13'b0_0_0_0_10101010_1;
      patterns[7209] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7210] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7211] = 13'b0_0_0_0_10101010_1;
      patterns[7212] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7213] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7214] = 13'b0_0_0_0_10101010_1;
      patterns[7215] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[7216] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[7217] = 13'b1_0_0_0_10101010_1;
      patterns[7218] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7219] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7220] = 13'b0_0_0_0_10101010_1;
      patterns[7221] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7222] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7223] = 13'b0_0_0_0_10101010_1;
      patterns[7224] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7225] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7226] = 13'b0_0_0_0_10101010_1;
      patterns[7227] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7228] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7229] = 13'b0_0_0_0_10101010_1;
      patterns[7230] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7231] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7232] = 13'b0_0_0_0_10101010_1;
      patterns[7233] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7234] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7235] = 13'b0_0_0_0_10101010_1;
      patterns[7236] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7237] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7238] = 13'b0_0_0_0_10101010_1;
      patterns[7239] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7240] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7241] = 13'b0_0_0_0_10101010_1;
      patterns[7242] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7243] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7244] = 13'b0_0_0_0_10101010_1;
      patterns[7245] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7246] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7247] = 13'b0_0_0_0_10101010_1;
      patterns[7248] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7249] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7250] = 13'b0_0_0_0_10101010_1;
      patterns[7251] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7252] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7253] = 13'b0_0_0_0_10101010_1;
      patterns[7254] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7255] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7256] = 13'b0_0_0_0_10101010_1;
      patterns[7257] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7258] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7259] = 13'b0_0_0_0_10101010_1;
      patterns[7260] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7261] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7262] = 13'b0_0_0_0_10101010_1;
      patterns[7263] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[7264] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[7265] = 13'b1_0_0_0_10101010_1;
      patterns[7266] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7267] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7268] = 13'b0_0_0_0_10101010_1;
      patterns[7269] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7270] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7271] = 13'b0_0_0_0_10101010_1;
      patterns[7272] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7273] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7274] = 13'b0_0_0_0_10101010_1;
      patterns[7275] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7276] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7277] = 13'b0_0_0_0_10101010_1;
      patterns[7278] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7279] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7280] = 13'b0_0_0_0_10101010_1;
      patterns[7281] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7282] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7283] = 13'b0_0_0_0_10101010_1;
      patterns[7284] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7285] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7286] = 13'b0_0_0_0_10101010_1;
      patterns[7287] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7288] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7289] = 13'b0_0_0_0_10101010_1;
      patterns[7290] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7291] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7292] = 13'b0_0_0_0_10101010_1;
      patterns[7293] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7294] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7295] = 13'b0_0_0_0_10101010_1;
      patterns[7296] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7297] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7298] = 13'b0_0_0_0_10101010_1;
      patterns[7299] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7300] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7301] = 13'b0_0_0_0_10101010_1;
      patterns[7302] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7303] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7304] = 13'b0_0_0_0_10101010_1;
      patterns[7305] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7306] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7307] = 13'b0_0_0_0_10101010_1;
      patterns[7308] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7309] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7310] = 13'b0_0_0_0_10101010_1;
      patterns[7311] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[7312] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[7313] = 13'b1_0_0_0_10101010_1;
      patterns[7314] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7315] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7316] = 13'b0_0_0_0_10101010_1;
      patterns[7317] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7318] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7319] = 13'b0_0_0_0_10101010_1;
      patterns[7320] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7321] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7322] = 13'b0_0_0_0_10101010_1;
      patterns[7323] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7324] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7325] = 13'b0_0_0_0_10101010_1;
      patterns[7326] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7327] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7328] = 13'b0_0_0_0_10101010_1;
      patterns[7329] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7330] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7331] = 13'b0_0_0_0_10101010_1;
      patterns[7332] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7333] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7334] = 13'b0_0_0_0_10101010_1;
      patterns[7335] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7336] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7337] = 13'b0_0_0_0_10101010_1;
      patterns[7338] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7339] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7340] = 13'b0_0_0_0_10101010_1;
      patterns[7341] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7342] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7343] = 13'b0_0_0_0_10101010_1;
      patterns[7344] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7345] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7346] = 13'b0_0_0_0_10101010_1;
      patterns[7347] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7348] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7349] = 13'b0_0_0_0_10101010_1;
      patterns[7350] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7351] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7352] = 13'b0_0_0_0_10101010_1;
      patterns[7353] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7354] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7355] = 13'b0_0_0_0_10101010_1;
      patterns[7356] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7357] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7358] = 13'b0_0_0_0_10101010_1;
      patterns[7359] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[7360] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[7361] = 13'b1_0_0_0_10101010_1;
      patterns[7362] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7363] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7364] = 13'b0_0_0_0_10101010_1;
      patterns[7365] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7366] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7367] = 13'b0_0_0_0_10101010_1;
      patterns[7368] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7369] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7370] = 13'b0_0_0_0_10101010_1;
      patterns[7371] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7372] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7373] = 13'b0_0_0_0_10101010_1;
      patterns[7374] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7375] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7376] = 13'b0_0_0_0_10101010_1;
      patterns[7377] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7378] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7379] = 13'b0_0_0_0_10101010_1;
      patterns[7380] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7381] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7382] = 13'b0_0_0_0_10101010_1;
      patterns[7383] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7384] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7385] = 13'b0_0_0_0_10101010_1;
      patterns[7386] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7387] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7388] = 13'b0_0_0_0_10101010_1;
      patterns[7389] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7390] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7391] = 13'b0_0_0_0_10101010_1;
      patterns[7392] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7393] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7394] = 13'b0_0_0_0_10101010_1;
      patterns[7395] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7396] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7397] = 13'b0_0_0_0_10101010_1;
      patterns[7398] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7399] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7400] = 13'b0_0_0_0_10101010_1;
      patterns[7401] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7402] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7403] = 13'b0_0_0_0_10101010_1;
      patterns[7404] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7405] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7406] = 13'b0_0_0_0_10101010_1;
      patterns[7407] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[7408] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[7409] = 13'b1_0_0_0_10101010_1;
      patterns[7410] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7411] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7412] = 13'b0_0_0_0_10101010_1;
      patterns[7413] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7414] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7415] = 13'b0_0_0_0_10101010_1;
      patterns[7416] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7417] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7418] = 13'b0_0_0_0_10101010_1;
      patterns[7419] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7420] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7421] = 13'b0_0_0_0_10101010_1;
      patterns[7422] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7423] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7424] = 13'b0_0_0_0_10101010_1;
      patterns[7425] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7426] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7427] = 13'b0_0_0_0_10101010_1;
      patterns[7428] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7429] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7430] = 13'b0_0_0_0_10101010_1;
      patterns[7431] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7432] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7433] = 13'b0_0_0_0_10101010_1;
      patterns[7434] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7435] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7436] = 13'b0_0_0_0_10101010_1;
      patterns[7437] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7438] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7439] = 13'b0_0_0_0_10101010_1;
      patterns[7440] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7441] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7442] = 13'b0_0_0_0_10101010_1;
      patterns[7443] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7444] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7445] = 13'b0_0_0_0_10101010_1;
      patterns[7446] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7447] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7448] = 13'b0_0_0_0_10101010_1;
      patterns[7449] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7450] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7451] = 13'b0_0_0_0_10101010_1;
      patterns[7452] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7453] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7454] = 13'b0_0_0_0_10101010_1;
      patterns[7455] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[7456] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[7457] = 13'b1_0_0_0_10101010_1;
      patterns[7458] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7459] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7460] = 13'b0_0_0_0_10101010_1;
      patterns[7461] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7462] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7463] = 13'b0_0_0_0_10101010_1;
      patterns[7464] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7465] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7466] = 13'b0_0_0_0_10101010_1;
      patterns[7467] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7468] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7469] = 13'b0_0_0_0_10101010_1;
      patterns[7470] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7471] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7472] = 13'b0_0_0_0_10101010_1;
      patterns[7473] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7474] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7475] = 13'b0_0_0_0_10101010_1;
      patterns[7476] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7477] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7478] = 13'b0_0_0_0_10101010_1;
      patterns[7479] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7480] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7481] = 13'b0_0_0_0_10101010_1;
      patterns[7482] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7483] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7484] = 13'b0_0_0_0_10101010_1;
      patterns[7485] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7486] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7487] = 13'b0_0_0_0_10101010_1;
      patterns[7488] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7489] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7490] = 13'b0_0_0_0_10101010_1;
      patterns[7491] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7492] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7493] = 13'b0_0_0_0_10101010_1;
      patterns[7494] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7495] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7496] = 13'b0_0_0_0_10101010_1;
      patterns[7497] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7498] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7499] = 13'b0_0_0_0_10101010_1;
      patterns[7500] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7501] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7502] = 13'b0_0_0_0_10101010_1;
      patterns[7503] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[7504] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[7505] = 13'b1_0_0_0_10101010_1;
      patterns[7506] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7507] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7508] = 13'b0_0_0_0_10101010_1;
      patterns[7509] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7510] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7511] = 13'b0_0_0_0_10101010_1;
      patterns[7512] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7513] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7514] = 13'b0_0_0_0_10101010_1;
      patterns[7515] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7516] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7517] = 13'b0_0_0_0_10101010_1;
      patterns[7518] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7519] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7520] = 13'b0_0_0_0_10101010_1;
      patterns[7521] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7522] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7523] = 13'b0_0_0_0_10101010_1;
      patterns[7524] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7525] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7526] = 13'b0_0_0_0_10101010_1;
      patterns[7527] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7528] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7529] = 13'b0_0_0_0_10101010_1;
      patterns[7530] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7531] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7532] = 13'b0_0_0_0_10101010_1;
      patterns[7533] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7534] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7535] = 13'b0_0_0_0_10101010_1;
      patterns[7536] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7537] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7538] = 13'b0_0_0_0_10101010_1;
      patterns[7539] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7540] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7541] = 13'b0_0_0_0_10101010_1;
      patterns[7542] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7543] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7544] = 13'b0_0_0_0_10101010_1;
      patterns[7545] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7546] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7547] = 13'b0_0_0_0_10101010_1;
      patterns[7548] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7549] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7550] = 13'b0_0_0_0_10101010_1;
      patterns[7551] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[7552] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[7553] = 13'b1_0_0_0_10101010_1;
      patterns[7554] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7555] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7556] = 13'b0_0_0_0_10101010_1;
      patterns[7557] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7558] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7559] = 13'b0_0_0_0_10101010_1;
      patterns[7560] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7561] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7562] = 13'b0_0_0_0_10101010_1;
      patterns[7563] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7564] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7565] = 13'b0_0_0_0_10101010_1;
      patterns[7566] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7567] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7568] = 13'b0_0_0_0_10101010_1;
      patterns[7569] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7570] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7571] = 13'b0_0_0_0_10101010_1;
      patterns[7572] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7573] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7574] = 13'b0_0_0_0_10101010_1;
      patterns[7575] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7576] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7577] = 13'b0_0_0_0_10101010_1;
      patterns[7578] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7579] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7580] = 13'b0_0_0_0_10101010_1;
      patterns[7581] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7582] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7583] = 13'b0_0_0_0_10101010_1;
      patterns[7584] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7585] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7586] = 13'b0_0_0_0_10101010_1;
      patterns[7587] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7588] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7589] = 13'b0_0_0_0_10101010_1;
      patterns[7590] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7591] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7592] = 13'b0_0_0_0_10101010_1;
      patterns[7593] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7594] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7595] = 13'b0_0_0_0_10101010_1;
      patterns[7596] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7597] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7598] = 13'b0_0_0_0_10101010_1;
      patterns[7599] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[7600] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[7601] = 13'b1_0_0_0_10101010_1;
      patterns[7602] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7603] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7604] = 13'b0_0_0_0_10101010_1;
      patterns[7605] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7606] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7607] = 13'b0_0_0_0_10101010_1;
      patterns[7608] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7609] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7610] = 13'b0_0_0_0_10101010_1;
      patterns[7611] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7612] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7613] = 13'b0_0_0_0_10101010_1;
      patterns[7614] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7615] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7616] = 13'b0_0_0_0_10101010_1;
      patterns[7617] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7618] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7619] = 13'b0_0_0_0_10101010_1;
      patterns[7620] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7621] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7622] = 13'b0_0_0_0_10101010_1;
      patterns[7623] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7624] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7625] = 13'b0_0_0_0_10101010_1;
      patterns[7626] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7627] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7628] = 13'b0_0_0_0_10101010_1;
      patterns[7629] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7630] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7631] = 13'b0_0_0_0_10101010_1;
      patterns[7632] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7633] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7634] = 13'b0_0_0_0_10101010_1;
      patterns[7635] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7636] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7637] = 13'b0_0_0_0_10101010_1;
      patterns[7638] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7639] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7640] = 13'b0_0_0_0_10101010_1;
      patterns[7641] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7642] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7643] = 13'b0_0_0_0_10101010_1;
      patterns[7644] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7645] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7646] = 13'b0_0_0_0_10101010_1;
      patterns[7647] = 13'b1_0_0_0_xxxxxxxx_x;
      patterns[7648] = 13'b1_0_1_0_xxxxxxxx_x;
      patterns[7649] = 13'b1_0_0_0_10101010_1;
      patterns[7650] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7651] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7652] = 13'b0_0_0_0_10101010_1;
      patterns[7653] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7654] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7655] = 13'b0_0_0_0_10101010_1;
      patterns[7656] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7657] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7658] = 13'b0_0_0_0_10101010_1;
      patterns[7659] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7660] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7661] = 13'b0_0_0_0_10101010_1;
      patterns[7662] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7663] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7664] = 13'b0_0_0_0_10101010_1;
      patterns[7665] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7666] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7667] = 13'b0_0_0_0_10101010_1;
      patterns[7668] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7669] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7670] = 13'b0_0_0_0_10101010_1;
      patterns[7671] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7672] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7673] = 13'b0_0_0_0_10101010_1;
      patterns[7674] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7675] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7676] = 13'b0_0_0_0_10101010_1;
      patterns[7677] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7678] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7679] = 13'b0_0_0_0_10101010_1;
      patterns[7680] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7681] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7682] = 13'b0_0_0_0_10101010_1;
      patterns[7683] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7684] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7685] = 13'b0_0_0_0_10101010_1;
      patterns[7686] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7687] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7688] = 13'b0_0_0_0_10101010_1;
      patterns[7689] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7690] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7691] = 13'b0_0_0_0_10101010_1;
      patterns[7692] = 13'b0_0_0_0_xxxxxxxx_x;
      patterns[7693] = 13'b0_0_1_0_xxxxxxxx_x;
      patterns[7694] = 13'b0_0_0_0_10101010_1;

      for (i = 0; i < 7695; i = i + 1)
      begin
        en = patterns[i][12];
        CDP = patterns[i][11];
        clk16 = patterns[i][10];
        RX = patterns[i][9];
        #10;
        if (patterns[i][8:1] !== 8'hx)
        begin
          if (DATA !== patterns[i][8:1])
          begin
            $display("%d:DATA: (assertion error). Expected %h, found %h", i, patterns[i][8:1], DATA);
            $finish;
          end
        end
        if (patterns[i][0] !== 1'hx)
        begin
          if (DP !== patterns[i][0])
          begin
            $display("%d:DP: (assertion error). Expected %h, found %h", i, patterns[i][0], DP);
            $finish;
          end
        end
      end

      $display("All tests passed.");
    end
    endmodule
