`timescale 1us/1ns

module ROTATER_tb;
    reg [2:0] OP;
    reg [11:0] AI;
    reg LI;
    reg OE;
    wire [11:0] AO;
    wire LO;

  ROTATER dut (
    .OP(OP),
    .AI(AI),
    .LI(LI),
    .OE(OE),
    .AO(AO),
    .LO(LO)
  );

    reg [28:0] patterns[0:65535];
    integer i;

    initial begin
      OE=1;
      patterns[0] = 29'b0_000000000000_000_0_000000000000;
      patterns[1] = 29'b0_000000000000_001_0_000000000000;
      patterns[2] = 29'b0_000000000000_010_0_000000000000;
      patterns[3] = 29'b0_000000000000_011_0_000000000000;
      patterns[4] = 29'b0_000000000000_100_0_000000000000;
      patterns[5] = 29'b0_000000000000_101_0_000000000000;
      patterns[6] = 29'b0_000000000000_110_0_000000000000;
      patterns[7] = 29'b0_000000000000_111_0_000000000000;
      patterns[8] = 29'b0_000000000001_000_0_000000000001;
      patterns[9] = 29'b0_000000000001_001_0_000001000000;
      patterns[10] = 29'b0_000000000001_010_0_000000000010;
      patterns[11] = 29'b0_000000000001_011_0_000000000100;
      patterns[12] = 29'b0_000000000001_100_1_000000000000;
      patterns[13] = 29'b0_000000000001_101_0_100000000000;
      patterns[14] = 29'b0_000000000001_110_0_000000000001;
      patterns[15] = 29'b0_000000000001_111_0_000000000001;
      patterns[16] = 29'b0_000000000010_000_0_000000000010;
      patterns[17] = 29'b0_000000000010_001_0_000010000000;
      patterns[18] = 29'b0_000000000010_010_0_000000000100;
      patterns[19] = 29'b0_000000000010_011_0_000000001000;
      patterns[20] = 29'b0_000000000010_100_0_000000000001;
      patterns[21] = 29'b0_000000000010_101_1_000000000000;
      patterns[22] = 29'b0_000000000010_110_0_000000000010;
      patterns[23] = 29'b0_000000000010_111_0_000000000010;
      patterns[24] = 29'b0_000000000011_000_0_000000000011;
      patterns[25] = 29'b0_000000000011_001_0_000011000000;
      patterns[26] = 29'b0_000000000011_010_0_000000000110;
      patterns[27] = 29'b0_000000000011_011_0_000000001100;
      patterns[28] = 29'b0_000000000011_100_1_000000000001;
      patterns[29] = 29'b0_000000000011_101_1_100000000000;
      patterns[30] = 29'b0_000000000011_110_0_000000000011;
      patterns[31] = 29'b0_000000000011_111_0_000000000011;
      patterns[32] = 29'b0_000000000100_000_0_000000000100;
      patterns[33] = 29'b0_000000000100_001_0_000100000000;
      patterns[34] = 29'b0_000000000100_010_0_000000001000;
      patterns[35] = 29'b0_000000000100_011_0_000000010000;
      patterns[36] = 29'b0_000000000100_100_0_000000000010;
      patterns[37] = 29'b0_000000000100_101_0_000000000001;
      patterns[38] = 29'b0_000000000100_110_0_000000000100;
      patterns[39] = 29'b0_000000000100_111_0_000000000100;
      patterns[40] = 29'b0_000000000101_000_0_000000000101;
      patterns[41] = 29'b0_000000000101_001_0_000101000000;
      patterns[42] = 29'b0_000000000101_010_0_000000001010;
      patterns[43] = 29'b0_000000000101_011_0_000000010100;
      patterns[44] = 29'b0_000000000101_100_1_000000000010;
      patterns[45] = 29'b0_000000000101_101_0_100000000001;
      patterns[46] = 29'b0_000000000101_110_0_000000000101;
      patterns[47] = 29'b0_000000000101_111_0_000000000101;
      patterns[48] = 29'b0_000000000110_000_0_000000000110;
      patterns[49] = 29'b0_000000000110_001_0_000110000000;
      patterns[50] = 29'b0_000000000110_010_0_000000001100;
      patterns[51] = 29'b0_000000000110_011_0_000000011000;
      patterns[52] = 29'b0_000000000110_100_0_000000000011;
      patterns[53] = 29'b0_000000000110_101_1_000000000001;
      patterns[54] = 29'b0_000000000110_110_0_000000000110;
      patterns[55] = 29'b0_000000000110_111_0_000000000110;
      patterns[56] = 29'b0_000000000111_000_0_000000000111;
      patterns[57] = 29'b0_000000000111_001_0_000111000000;
      patterns[58] = 29'b0_000000000111_010_0_000000001110;
      patterns[59] = 29'b0_000000000111_011_0_000000011100;
      patterns[60] = 29'b0_000000000111_100_1_000000000011;
      patterns[61] = 29'b0_000000000111_101_1_100000000001;
      patterns[62] = 29'b0_000000000111_110_0_000000000111;
      patterns[63] = 29'b0_000000000111_111_0_000000000111;
      patterns[64] = 29'b0_000000001000_000_0_000000001000;
      patterns[65] = 29'b0_000000001000_001_0_001000000000;
      patterns[66] = 29'b0_000000001000_010_0_000000010000;
      patterns[67] = 29'b0_000000001000_011_0_000000100000;
      patterns[68] = 29'b0_000000001000_100_0_000000000100;
      patterns[69] = 29'b0_000000001000_101_0_000000000010;
      patterns[70] = 29'b0_000000001000_110_0_000000001000;
      patterns[71] = 29'b0_000000001000_111_0_000000001000;
      patterns[72] = 29'b0_000000001001_000_0_000000001001;
      patterns[73] = 29'b0_000000001001_001_0_001001000000;
      patterns[74] = 29'b0_000000001001_010_0_000000010010;
      patterns[75] = 29'b0_000000001001_011_0_000000100100;
      patterns[76] = 29'b0_000000001001_100_1_000000000100;
      patterns[77] = 29'b0_000000001001_101_0_100000000010;
      patterns[78] = 29'b0_000000001001_110_0_000000001001;
      patterns[79] = 29'b0_000000001001_111_0_000000001001;
      patterns[80] = 29'b0_000000001010_000_0_000000001010;
      patterns[81] = 29'b0_000000001010_001_0_001010000000;
      patterns[82] = 29'b0_000000001010_010_0_000000010100;
      patterns[83] = 29'b0_000000001010_011_0_000000101000;
      patterns[84] = 29'b0_000000001010_100_0_000000000101;
      patterns[85] = 29'b0_000000001010_101_1_000000000010;
      patterns[86] = 29'b0_000000001010_110_0_000000001010;
      patterns[87] = 29'b0_000000001010_111_0_000000001010;
      patterns[88] = 29'b0_000000001011_000_0_000000001011;
      patterns[89] = 29'b0_000000001011_001_0_001011000000;
      patterns[90] = 29'b0_000000001011_010_0_000000010110;
      patterns[91] = 29'b0_000000001011_011_0_000000101100;
      patterns[92] = 29'b0_000000001011_100_1_000000000101;
      patterns[93] = 29'b0_000000001011_101_1_100000000010;
      patterns[94] = 29'b0_000000001011_110_0_000000001011;
      patterns[95] = 29'b0_000000001011_111_0_000000001011;
      patterns[96] = 29'b0_000000001100_000_0_000000001100;
      patterns[97] = 29'b0_000000001100_001_0_001100000000;
      patterns[98] = 29'b0_000000001100_010_0_000000011000;
      patterns[99] = 29'b0_000000001100_011_0_000000110000;
      patterns[100] = 29'b0_000000001100_100_0_000000000110;
      patterns[101] = 29'b0_000000001100_101_0_000000000011;
      patterns[102] = 29'b0_000000001100_110_0_000000001100;
      patterns[103] = 29'b0_000000001100_111_0_000000001100;
      patterns[104] = 29'b0_000000001101_000_0_000000001101;
      patterns[105] = 29'b0_000000001101_001_0_001101000000;
      patterns[106] = 29'b0_000000001101_010_0_000000011010;
      patterns[107] = 29'b0_000000001101_011_0_000000110100;
      patterns[108] = 29'b0_000000001101_100_1_000000000110;
      patterns[109] = 29'b0_000000001101_101_0_100000000011;
      patterns[110] = 29'b0_000000001101_110_0_000000001101;
      patterns[111] = 29'b0_000000001101_111_0_000000001101;
      patterns[112] = 29'b0_000000001110_000_0_000000001110;
      patterns[113] = 29'b0_000000001110_001_0_001110000000;
      patterns[114] = 29'b0_000000001110_010_0_000000011100;
      patterns[115] = 29'b0_000000001110_011_0_000000111000;
      patterns[116] = 29'b0_000000001110_100_0_000000000111;
      patterns[117] = 29'b0_000000001110_101_1_000000000011;
      patterns[118] = 29'b0_000000001110_110_0_000000001110;
      patterns[119] = 29'b0_000000001110_111_0_000000001110;
      patterns[120] = 29'b0_000000001111_000_0_000000001111;
      patterns[121] = 29'b0_000000001111_001_0_001111000000;
      patterns[122] = 29'b0_000000001111_010_0_000000011110;
      patterns[123] = 29'b0_000000001111_011_0_000000111100;
      patterns[124] = 29'b0_000000001111_100_1_000000000111;
      patterns[125] = 29'b0_000000001111_101_1_100000000011;
      patterns[126] = 29'b0_000000001111_110_0_000000001111;
      patterns[127] = 29'b0_000000001111_111_0_000000001111;
      patterns[128] = 29'b0_000000010000_000_0_000000010000;
      patterns[129] = 29'b0_000000010000_001_0_010000000000;
      patterns[130] = 29'b0_000000010000_010_0_000000100000;
      patterns[131] = 29'b0_000000010000_011_0_000001000000;
      patterns[132] = 29'b0_000000010000_100_0_000000001000;
      patterns[133] = 29'b0_000000010000_101_0_000000000100;
      patterns[134] = 29'b0_000000010000_110_0_000000010000;
      patterns[135] = 29'b0_000000010000_111_0_000000010000;
      patterns[136] = 29'b0_000000010001_000_0_000000010001;
      patterns[137] = 29'b0_000000010001_001_0_010001000000;
      patterns[138] = 29'b0_000000010001_010_0_000000100010;
      patterns[139] = 29'b0_000000010001_011_0_000001000100;
      patterns[140] = 29'b0_000000010001_100_1_000000001000;
      patterns[141] = 29'b0_000000010001_101_0_100000000100;
      patterns[142] = 29'b0_000000010001_110_0_000000010001;
      patterns[143] = 29'b0_000000010001_111_0_000000010001;
      patterns[144] = 29'b0_000000010010_000_0_000000010010;
      patterns[145] = 29'b0_000000010010_001_0_010010000000;
      patterns[146] = 29'b0_000000010010_010_0_000000100100;
      patterns[147] = 29'b0_000000010010_011_0_000001001000;
      patterns[148] = 29'b0_000000010010_100_0_000000001001;
      patterns[149] = 29'b0_000000010010_101_1_000000000100;
      patterns[150] = 29'b0_000000010010_110_0_000000010010;
      patterns[151] = 29'b0_000000010010_111_0_000000010010;
      patterns[152] = 29'b0_000000010011_000_0_000000010011;
      patterns[153] = 29'b0_000000010011_001_0_010011000000;
      patterns[154] = 29'b0_000000010011_010_0_000000100110;
      patterns[155] = 29'b0_000000010011_011_0_000001001100;
      patterns[156] = 29'b0_000000010011_100_1_000000001001;
      patterns[157] = 29'b0_000000010011_101_1_100000000100;
      patterns[158] = 29'b0_000000010011_110_0_000000010011;
      patterns[159] = 29'b0_000000010011_111_0_000000010011;
      patterns[160] = 29'b0_000000010100_000_0_000000010100;
      patterns[161] = 29'b0_000000010100_001_0_010100000000;
      patterns[162] = 29'b0_000000010100_010_0_000000101000;
      patterns[163] = 29'b0_000000010100_011_0_000001010000;
      patterns[164] = 29'b0_000000010100_100_0_000000001010;
      patterns[165] = 29'b0_000000010100_101_0_000000000101;
      patterns[166] = 29'b0_000000010100_110_0_000000010100;
      patterns[167] = 29'b0_000000010100_111_0_000000010100;
      patterns[168] = 29'b0_000000010101_000_0_000000010101;
      patterns[169] = 29'b0_000000010101_001_0_010101000000;
      patterns[170] = 29'b0_000000010101_010_0_000000101010;
      patterns[171] = 29'b0_000000010101_011_0_000001010100;
      patterns[172] = 29'b0_000000010101_100_1_000000001010;
      patterns[173] = 29'b0_000000010101_101_0_100000000101;
      patterns[174] = 29'b0_000000010101_110_0_000000010101;
      patterns[175] = 29'b0_000000010101_111_0_000000010101;
      patterns[176] = 29'b0_000000010110_000_0_000000010110;
      patterns[177] = 29'b0_000000010110_001_0_010110000000;
      patterns[178] = 29'b0_000000010110_010_0_000000101100;
      patterns[179] = 29'b0_000000010110_011_0_000001011000;
      patterns[180] = 29'b0_000000010110_100_0_000000001011;
      patterns[181] = 29'b0_000000010110_101_1_000000000101;
      patterns[182] = 29'b0_000000010110_110_0_000000010110;
      patterns[183] = 29'b0_000000010110_111_0_000000010110;
      patterns[184] = 29'b0_000000010111_000_0_000000010111;
      patterns[185] = 29'b0_000000010111_001_0_010111000000;
      patterns[186] = 29'b0_000000010111_010_0_000000101110;
      patterns[187] = 29'b0_000000010111_011_0_000001011100;
      patterns[188] = 29'b0_000000010111_100_1_000000001011;
      patterns[189] = 29'b0_000000010111_101_1_100000000101;
      patterns[190] = 29'b0_000000010111_110_0_000000010111;
      patterns[191] = 29'b0_000000010111_111_0_000000010111;
      patterns[192] = 29'b0_000000011000_000_0_000000011000;
      patterns[193] = 29'b0_000000011000_001_0_011000000000;
      patterns[194] = 29'b0_000000011000_010_0_000000110000;
      patterns[195] = 29'b0_000000011000_011_0_000001100000;
      patterns[196] = 29'b0_000000011000_100_0_000000001100;
      patterns[197] = 29'b0_000000011000_101_0_000000000110;
      patterns[198] = 29'b0_000000011000_110_0_000000011000;
      patterns[199] = 29'b0_000000011000_111_0_000000011000;
      patterns[200] = 29'b0_000000011001_000_0_000000011001;
      patterns[201] = 29'b0_000000011001_001_0_011001000000;
      patterns[202] = 29'b0_000000011001_010_0_000000110010;
      patterns[203] = 29'b0_000000011001_011_0_000001100100;
      patterns[204] = 29'b0_000000011001_100_1_000000001100;
      patterns[205] = 29'b0_000000011001_101_0_100000000110;
      patterns[206] = 29'b0_000000011001_110_0_000000011001;
      patterns[207] = 29'b0_000000011001_111_0_000000011001;
      patterns[208] = 29'b0_000000011010_000_0_000000011010;
      patterns[209] = 29'b0_000000011010_001_0_011010000000;
      patterns[210] = 29'b0_000000011010_010_0_000000110100;
      patterns[211] = 29'b0_000000011010_011_0_000001101000;
      patterns[212] = 29'b0_000000011010_100_0_000000001101;
      patterns[213] = 29'b0_000000011010_101_1_000000000110;
      patterns[214] = 29'b0_000000011010_110_0_000000011010;
      patterns[215] = 29'b0_000000011010_111_0_000000011010;
      patterns[216] = 29'b0_000000011011_000_0_000000011011;
      patterns[217] = 29'b0_000000011011_001_0_011011000000;
      patterns[218] = 29'b0_000000011011_010_0_000000110110;
      patterns[219] = 29'b0_000000011011_011_0_000001101100;
      patterns[220] = 29'b0_000000011011_100_1_000000001101;
      patterns[221] = 29'b0_000000011011_101_1_100000000110;
      patterns[222] = 29'b0_000000011011_110_0_000000011011;
      patterns[223] = 29'b0_000000011011_111_0_000000011011;
      patterns[224] = 29'b0_000000011100_000_0_000000011100;
      patterns[225] = 29'b0_000000011100_001_0_011100000000;
      patterns[226] = 29'b0_000000011100_010_0_000000111000;
      patterns[227] = 29'b0_000000011100_011_0_000001110000;
      patterns[228] = 29'b0_000000011100_100_0_000000001110;
      patterns[229] = 29'b0_000000011100_101_0_000000000111;
      patterns[230] = 29'b0_000000011100_110_0_000000011100;
      patterns[231] = 29'b0_000000011100_111_0_000000011100;
      patterns[232] = 29'b0_000000011101_000_0_000000011101;
      patterns[233] = 29'b0_000000011101_001_0_011101000000;
      patterns[234] = 29'b0_000000011101_010_0_000000111010;
      patterns[235] = 29'b0_000000011101_011_0_000001110100;
      patterns[236] = 29'b0_000000011101_100_1_000000001110;
      patterns[237] = 29'b0_000000011101_101_0_100000000111;
      patterns[238] = 29'b0_000000011101_110_0_000000011101;
      patterns[239] = 29'b0_000000011101_111_0_000000011101;
      patterns[240] = 29'b0_000000011110_000_0_000000011110;
      patterns[241] = 29'b0_000000011110_001_0_011110000000;
      patterns[242] = 29'b0_000000011110_010_0_000000111100;
      patterns[243] = 29'b0_000000011110_011_0_000001111000;
      patterns[244] = 29'b0_000000011110_100_0_000000001111;
      patterns[245] = 29'b0_000000011110_101_1_000000000111;
      patterns[246] = 29'b0_000000011110_110_0_000000011110;
      patterns[247] = 29'b0_000000011110_111_0_000000011110;
      patterns[248] = 29'b0_000000011111_000_0_000000011111;
      patterns[249] = 29'b0_000000011111_001_0_011111000000;
      patterns[250] = 29'b0_000000011111_010_0_000000111110;
      patterns[251] = 29'b0_000000011111_011_0_000001111100;
      patterns[252] = 29'b0_000000011111_100_1_000000001111;
      patterns[253] = 29'b0_000000011111_101_1_100000000111;
      patterns[254] = 29'b0_000000011111_110_0_000000011111;
      patterns[255] = 29'b0_000000011111_111_0_000000011111;
      patterns[256] = 29'b0_000000100000_000_0_000000100000;
      patterns[257] = 29'b0_000000100000_001_0_100000000000;
      patterns[258] = 29'b0_000000100000_010_0_000001000000;
      patterns[259] = 29'b0_000000100000_011_0_000010000000;
      patterns[260] = 29'b0_000000100000_100_0_000000010000;
      patterns[261] = 29'b0_000000100000_101_0_000000001000;
      patterns[262] = 29'b0_000000100000_110_0_000000100000;
      patterns[263] = 29'b0_000000100000_111_0_000000100000;
      patterns[264] = 29'b0_000000100001_000_0_000000100001;
      patterns[265] = 29'b0_000000100001_001_0_100001000000;
      patterns[266] = 29'b0_000000100001_010_0_000001000010;
      patterns[267] = 29'b0_000000100001_011_0_000010000100;
      patterns[268] = 29'b0_000000100001_100_1_000000010000;
      patterns[269] = 29'b0_000000100001_101_0_100000001000;
      patterns[270] = 29'b0_000000100001_110_0_000000100001;
      patterns[271] = 29'b0_000000100001_111_0_000000100001;
      patterns[272] = 29'b0_000000100010_000_0_000000100010;
      patterns[273] = 29'b0_000000100010_001_0_100010000000;
      patterns[274] = 29'b0_000000100010_010_0_000001000100;
      patterns[275] = 29'b0_000000100010_011_0_000010001000;
      patterns[276] = 29'b0_000000100010_100_0_000000010001;
      patterns[277] = 29'b0_000000100010_101_1_000000001000;
      patterns[278] = 29'b0_000000100010_110_0_000000100010;
      patterns[279] = 29'b0_000000100010_111_0_000000100010;
      patterns[280] = 29'b0_000000100011_000_0_000000100011;
      patterns[281] = 29'b0_000000100011_001_0_100011000000;
      patterns[282] = 29'b0_000000100011_010_0_000001000110;
      patterns[283] = 29'b0_000000100011_011_0_000010001100;
      patterns[284] = 29'b0_000000100011_100_1_000000010001;
      patterns[285] = 29'b0_000000100011_101_1_100000001000;
      patterns[286] = 29'b0_000000100011_110_0_000000100011;
      patterns[287] = 29'b0_000000100011_111_0_000000100011;
      patterns[288] = 29'b0_000000100100_000_0_000000100100;
      patterns[289] = 29'b0_000000100100_001_0_100100000000;
      patterns[290] = 29'b0_000000100100_010_0_000001001000;
      patterns[291] = 29'b0_000000100100_011_0_000010010000;
      patterns[292] = 29'b0_000000100100_100_0_000000010010;
      patterns[293] = 29'b0_000000100100_101_0_000000001001;
      patterns[294] = 29'b0_000000100100_110_0_000000100100;
      patterns[295] = 29'b0_000000100100_111_0_000000100100;
      patterns[296] = 29'b0_000000100101_000_0_000000100101;
      patterns[297] = 29'b0_000000100101_001_0_100101000000;
      patterns[298] = 29'b0_000000100101_010_0_000001001010;
      patterns[299] = 29'b0_000000100101_011_0_000010010100;
      patterns[300] = 29'b0_000000100101_100_1_000000010010;
      patterns[301] = 29'b0_000000100101_101_0_100000001001;
      patterns[302] = 29'b0_000000100101_110_0_000000100101;
      patterns[303] = 29'b0_000000100101_111_0_000000100101;
      patterns[304] = 29'b0_000000100110_000_0_000000100110;
      patterns[305] = 29'b0_000000100110_001_0_100110000000;
      patterns[306] = 29'b0_000000100110_010_0_000001001100;
      patterns[307] = 29'b0_000000100110_011_0_000010011000;
      patterns[308] = 29'b0_000000100110_100_0_000000010011;
      patterns[309] = 29'b0_000000100110_101_1_000000001001;
      patterns[310] = 29'b0_000000100110_110_0_000000100110;
      patterns[311] = 29'b0_000000100110_111_0_000000100110;
      patterns[312] = 29'b0_000000100111_000_0_000000100111;
      patterns[313] = 29'b0_000000100111_001_0_100111000000;
      patterns[314] = 29'b0_000000100111_010_0_000001001110;
      patterns[315] = 29'b0_000000100111_011_0_000010011100;
      patterns[316] = 29'b0_000000100111_100_1_000000010011;
      patterns[317] = 29'b0_000000100111_101_1_100000001001;
      patterns[318] = 29'b0_000000100111_110_0_000000100111;
      patterns[319] = 29'b0_000000100111_111_0_000000100111;
      patterns[320] = 29'b0_000000101000_000_0_000000101000;
      patterns[321] = 29'b0_000000101000_001_0_101000000000;
      patterns[322] = 29'b0_000000101000_010_0_000001010000;
      patterns[323] = 29'b0_000000101000_011_0_000010100000;
      patterns[324] = 29'b0_000000101000_100_0_000000010100;
      patterns[325] = 29'b0_000000101000_101_0_000000001010;
      patterns[326] = 29'b0_000000101000_110_0_000000101000;
      patterns[327] = 29'b0_000000101000_111_0_000000101000;
      patterns[328] = 29'b0_000000101001_000_0_000000101001;
      patterns[329] = 29'b0_000000101001_001_0_101001000000;
      patterns[330] = 29'b0_000000101001_010_0_000001010010;
      patterns[331] = 29'b0_000000101001_011_0_000010100100;
      patterns[332] = 29'b0_000000101001_100_1_000000010100;
      patterns[333] = 29'b0_000000101001_101_0_100000001010;
      patterns[334] = 29'b0_000000101001_110_0_000000101001;
      patterns[335] = 29'b0_000000101001_111_0_000000101001;
      patterns[336] = 29'b0_000000101010_000_0_000000101010;
      patterns[337] = 29'b0_000000101010_001_0_101010000000;
      patterns[338] = 29'b0_000000101010_010_0_000001010100;
      patterns[339] = 29'b0_000000101010_011_0_000010101000;
      patterns[340] = 29'b0_000000101010_100_0_000000010101;
      patterns[341] = 29'b0_000000101010_101_1_000000001010;
      patterns[342] = 29'b0_000000101010_110_0_000000101010;
      patterns[343] = 29'b0_000000101010_111_0_000000101010;
      patterns[344] = 29'b0_000000101011_000_0_000000101011;
      patterns[345] = 29'b0_000000101011_001_0_101011000000;
      patterns[346] = 29'b0_000000101011_010_0_000001010110;
      patterns[347] = 29'b0_000000101011_011_0_000010101100;
      patterns[348] = 29'b0_000000101011_100_1_000000010101;
      patterns[349] = 29'b0_000000101011_101_1_100000001010;
      patterns[350] = 29'b0_000000101011_110_0_000000101011;
      patterns[351] = 29'b0_000000101011_111_0_000000101011;
      patterns[352] = 29'b0_000000101100_000_0_000000101100;
      patterns[353] = 29'b0_000000101100_001_0_101100000000;
      patterns[354] = 29'b0_000000101100_010_0_000001011000;
      patterns[355] = 29'b0_000000101100_011_0_000010110000;
      patterns[356] = 29'b0_000000101100_100_0_000000010110;
      patterns[357] = 29'b0_000000101100_101_0_000000001011;
      patterns[358] = 29'b0_000000101100_110_0_000000101100;
      patterns[359] = 29'b0_000000101100_111_0_000000101100;
      patterns[360] = 29'b0_000000101101_000_0_000000101101;
      patterns[361] = 29'b0_000000101101_001_0_101101000000;
      patterns[362] = 29'b0_000000101101_010_0_000001011010;
      patterns[363] = 29'b0_000000101101_011_0_000010110100;
      patterns[364] = 29'b0_000000101101_100_1_000000010110;
      patterns[365] = 29'b0_000000101101_101_0_100000001011;
      patterns[366] = 29'b0_000000101101_110_0_000000101101;
      patterns[367] = 29'b0_000000101101_111_0_000000101101;
      patterns[368] = 29'b0_000000101110_000_0_000000101110;
      patterns[369] = 29'b0_000000101110_001_0_101110000000;
      patterns[370] = 29'b0_000000101110_010_0_000001011100;
      patterns[371] = 29'b0_000000101110_011_0_000010111000;
      patterns[372] = 29'b0_000000101110_100_0_000000010111;
      patterns[373] = 29'b0_000000101110_101_1_000000001011;
      patterns[374] = 29'b0_000000101110_110_0_000000101110;
      patterns[375] = 29'b0_000000101110_111_0_000000101110;
      patterns[376] = 29'b0_000000101111_000_0_000000101111;
      patterns[377] = 29'b0_000000101111_001_0_101111000000;
      patterns[378] = 29'b0_000000101111_010_0_000001011110;
      patterns[379] = 29'b0_000000101111_011_0_000010111100;
      patterns[380] = 29'b0_000000101111_100_1_000000010111;
      patterns[381] = 29'b0_000000101111_101_1_100000001011;
      patterns[382] = 29'b0_000000101111_110_0_000000101111;
      patterns[383] = 29'b0_000000101111_111_0_000000101111;
      patterns[384] = 29'b0_000000110000_000_0_000000110000;
      patterns[385] = 29'b0_000000110000_001_0_110000000000;
      patterns[386] = 29'b0_000000110000_010_0_000001100000;
      patterns[387] = 29'b0_000000110000_011_0_000011000000;
      patterns[388] = 29'b0_000000110000_100_0_000000011000;
      patterns[389] = 29'b0_000000110000_101_0_000000001100;
      patterns[390] = 29'b0_000000110000_110_0_000000110000;
      patterns[391] = 29'b0_000000110000_111_0_000000110000;
      patterns[392] = 29'b0_000000110001_000_0_000000110001;
      patterns[393] = 29'b0_000000110001_001_0_110001000000;
      patterns[394] = 29'b0_000000110001_010_0_000001100010;
      patterns[395] = 29'b0_000000110001_011_0_000011000100;
      patterns[396] = 29'b0_000000110001_100_1_000000011000;
      patterns[397] = 29'b0_000000110001_101_0_100000001100;
      patterns[398] = 29'b0_000000110001_110_0_000000110001;
      patterns[399] = 29'b0_000000110001_111_0_000000110001;
      patterns[400] = 29'b0_000000110010_000_0_000000110010;
      patterns[401] = 29'b0_000000110010_001_0_110010000000;
      patterns[402] = 29'b0_000000110010_010_0_000001100100;
      patterns[403] = 29'b0_000000110010_011_0_000011001000;
      patterns[404] = 29'b0_000000110010_100_0_000000011001;
      patterns[405] = 29'b0_000000110010_101_1_000000001100;
      patterns[406] = 29'b0_000000110010_110_0_000000110010;
      patterns[407] = 29'b0_000000110010_111_0_000000110010;
      patterns[408] = 29'b0_000000110011_000_0_000000110011;
      patterns[409] = 29'b0_000000110011_001_0_110011000000;
      patterns[410] = 29'b0_000000110011_010_0_000001100110;
      patterns[411] = 29'b0_000000110011_011_0_000011001100;
      patterns[412] = 29'b0_000000110011_100_1_000000011001;
      patterns[413] = 29'b0_000000110011_101_1_100000001100;
      patterns[414] = 29'b0_000000110011_110_0_000000110011;
      patterns[415] = 29'b0_000000110011_111_0_000000110011;
      patterns[416] = 29'b0_000000110100_000_0_000000110100;
      patterns[417] = 29'b0_000000110100_001_0_110100000000;
      patterns[418] = 29'b0_000000110100_010_0_000001101000;
      patterns[419] = 29'b0_000000110100_011_0_000011010000;
      patterns[420] = 29'b0_000000110100_100_0_000000011010;
      patterns[421] = 29'b0_000000110100_101_0_000000001101;
      patterns[422] = 29'b0_000000110100_110_0_000000110100;
      patterns[423] = 29'b0_000000110100_111_0_000000110100;
      patterns[424] = 29'b0_000000110101_000_0_000000110101;
      patterns[425] = 29'b0_000000110101_001_0_110101000000;
      patterns[426] = 29'b0_000000110101_010_0_000001101010;
      patterns[427] = 29'b0_000000110101_011_0_000011010100;
      patterns[428] = 29'b0_000000110101_100_1_000000011010;
      patterns[429] = 29'b0_000000110101_101_0_100000001101;
      patterns[430] = 29'b0_000000110101_110_0_000000110101;
      patterns[431] = 29'b0_000000110101_111_0_000000110101;
      patterns[432] = 29'b0_000000110110_000_0_000000110110;
      patterns[433] = 29'b0_000000110110_001_0_110110000000;
      patterns[434] = 29'b0_000000110110_010_0_000001101100;
      patterns[435] = 29'b0_000000110110_011_0_000011011000;
      patterns[436] = 29'b0_000000110110_100_0_000000011011;
      patterns[437] = 29'b0_000000110110_101_1_000000001101;
      patterns[438] = 29'b0_000000110110_110_0_000000110110;
      patterns[439] = 29'b0_000000110110_111_0_000000110110;
      patterns[440] = 29'b0_000000110111_000_0_000000110111;
      patterns[441] = 29'b0_000000110111_001_0_110111000000;
      patterns[442] = 29'b0_000000110111_010_0_000001101110;
      patterns[443] = 29'b0_000000110111_011_0_000011011100;
      patterns[444] = 29'b0_000000110111_100_1_000000011011;
      patterns[445] = 29'b0_000000110111_101_1_100000001101;
      patterns[446] = 29'b0_000000110111_110_0_000000110111;
      patterns[447] = 29'b0_000000110111_111_0_000000110111;
      patterns[448] = 29'b0_000000111000_000_0_000000111000;
      patterns[449] = 29'b0_000000111000_001_0_111000000000;
      patterns[450] = 29'b0_000000111000_010_0_000001110000;
      patterns[451] = 29'b0_000000111000_011_0_000011100000;
      patterns[452] = 29'b0_000000111000_100_0_000000011100;
      patterns[453] = 29'b0_000000111000_101_0_000000001110;
      patterns[454] = 29'b0_000000111000_110_0_000000111000;
      patterns[455] = 29'b0_000000111000_111_0_000000111000;
      patterns[456] = 29'b0_000000111001_000_0_000000111001;
      patterns[457] = 29'b0_000000111001_001_0_111001000000;
      patterns[458] = 29'b0_000000111001_010_0_000001110010;
      patterns[459] = 29'b0_000000111001_011_0_000011100100;
      patterns[460] = 29'b0_000000111001_100_1_000000011100;
      patterns[461] = 29'b0_000000111001_101_0_100000001110;
      patterns[462] = 29'b0_000000111001_110_0_000000111001;
      patterns[463] = 29'b0_000000111001_111_0_000000111001;
      patterns[464] = 29'b0_000000111010_000_0_000000111010;
      patterns[465] = 29'b0_000000111010_001_0_111010000000;
      patterns[466] = 29'b0_000000111010_010_0_000001110100;
      patterns[467] = 29'b0_000000111010_011_0_000011101000;
      patterns[468] = 29'b0_000000111010_100_0_000000011101;
      patterns[469] = 29'b0_000000111010_101_1_000000001110;
      patterns[470] = 29'b0_000000111010_110_0_000000111010;
      patterns[471] = 29'b0_000000111010_111_0_000000111010;
      patterns[472] = 29'b0_000000111011_000_0_000000111011;
      patterns[473] = 29'b0_000000111011_001_0_111011000000;
      patterns[474] = 29'b0_000000111011_010_0_000001110110;
      patterns[475] = 29'b0_000000111011_011_0_000011101100;
      patterns[476] = 29'b0_000000111011_100_1_000000011101;
      patterns[477] = 29'b0_000000111011_101_1_100000001110;
      patterns[478] = 29'b0_000000111011_110_0_000000111011;
      patterns[479] = 29'b0_000000111011_111_0_000000111011;
      patterns[480] = 29'b0_000000111100_000_0_000000111100;
      patterns[481] = 29'b0_000000111100_001_0_111100000000;
      patterns[482] = 29'b0_000000111100_010_0_000001111000;
      patterns[483] = 29'b0_000000111100_011_0_000011110000;
      patterns[484] = 29'b0_000000111100_100_0_000000011110;
      patterns[485] = 29'b0_000000111100_101_0_000000001111;
      patterns[486] = 29'b0_000000111100_110_0_000000111100;
      patterns[487] = 29'b0_000000111100_111_0_000000111100;
      patterns[488] = 29'b0_000000111101_000_0_000000111101;
      patterns[489] = 29'b0_000000111101_001_0_111101000000;
      patterns[490] = 29'b0_000000111101_010_0_000001111010;
      patterns[491] = 29'b0_000000111101_011_0_000011110100;
      patterns[492] = 29'b0_000000111101_100_1_000000011110;
      patterns[493] = 29'b0_000000111101_101_0_100000001111;
      patterns[494] = 29'b0_000000111101_110_0_000000111101;
      patterns[495] = 29'b0_000000111101_111_0_000000111101;
      patterns[496] = 29'b0_000000111110_000_0_000000111110;
      patterns[497] = 29'b0_000000111110_001_0_111110000000;
      patterns[498] = 29'b0_000000111110_010_0_000001111100;
      patterns[499] = 29'b0_000000111110_011_0_000011111000;
      patterns[500] = 29'b0_000000111110_100_0_000000011111;
      patterns[501] = 29'b0_000000111110_101_1_000000001111;
      patterns[502] = 29'b0_000000111110_110_0_000000111110;
      patterns[503] = 29'b0_000000111110_111_0_000000111110;
      patterns[504] = 29'b0_000000111111_000_0_000000111111;
      patterns[505] = 29'b0_000000111111_001_0_111111000000;
      patterns[506] = 29'b0_000000111111_010_0_000001111110;
      patterns[507] = 29'b0_000000111111_011_0_000011111100;
      patterns[508] = 29'b0_000000111111_100_1_000000011111;
      patterns[509] = 29'b0_000000111111_101_1_100000001111;
      patterns[510] = 29'b0_000000111111_110_0_000000111111;
      patterns[511] = 29'b0_000000111111_111_0_000000111111;
      patterns[512] = 29'b0_000001000000_000_0_000001000000;
      patterns[513] = 29'b0_000001000000_001_0_000000000001;
      patterns[514] = 29'b0_000001000000_010_0_000010000000;
      patterns[515] = 29'b0_000001000000_011_0_000100000000;
      patterns[516] = 29'b0_000001000000_100_0_000000100000;
      patterns[517] = 29'b0_000001000000_101_0_000000010000;
      patterns[518] = 29'b0_000001000000_110_0_000001000000;
      patterns[519] = 29'b0_000001000000_111_0_000001000000;
      patterns[520] = 29'b0_000001000001_000_0_000001000001;
      patterns[521] = 29'b0_000001000001_001_0_000001000001;
      patterns[522] = 29'b0_000001000001_010_0_000010000010;
      patterns[523] = 29'b0_000001000001_011_0_000100000100;
      patterns[524] = 29'b0_000001000001_100_1_000000100000;
      patterns[525] = 29'b0_000001000001_101_0_100000010000;
      patterns[526] = 29'b0_000001000001_110_0_000001000001;
      patterns[527] = 29'b0_000001000001_111_0_000001000001;
      patterns[528] = 29'b0_000001000010_000_0_000001000010;
      patterns[529] = 29'b0_000001000010_001_0_000010000001;
      patterns[530] = 29'b0_000001000010_010_0_000010000100;
      patterns[531] = 29'b0_000001000010_011_0_000100001000;
      patterns[532] = 29'b0_000001000010_100_0_000000100001;
      patterns[533] = 29'b0_000001000010_101_1_000000010000;
      patterns[534] = 29'b0_000001000010_110_0_000001000010;
      patterns[535] = 29'b0_000001000010_111_0_000001000010;
      patterns[536] = 29'b0_000001000011_000_0_000001000011;
      patterns[537] = 29'b0_000001000011_001_0_000011000001;
      patterns[538] = 29'b0_000001000011_010_0_000010000110;
      patterns[539] = 29'b0_000001000011_011_0_000100001100;
      patterns[540] = 29'b0_000001000011_100_1_000000100001;
      patterns[541] = 29'b0_000001000011_101_1_100000010000;
      patterns[542] = 29'b0_000001000011_110_0_000001000011;
      patterns[543] = 29'b0_000001000011_111_0_000001000011;
      patterns[544] = 29'b0_000001000100_000_0_000001000100;
      patterns[545] = 29'b0_000001000100_001_0_000100000001;
      patterns[546] = 29'b0_000001000100_010_0_000010001000;
      patterns[547] = 29'b0_000001000100_011_0_000100010000;
      patterns[548] = 29'b0_000001000100_100_0_000000100010;
      patterns[549] = 29'b0_000001000100_101_0_000000010001;
      patterns[550] = 29'b0_000001000100_110_0_000001000100;
      patterns[551] = 29'b0_000001000100_111_0_000001000100;
      patterns[552] = 29'b0_000001000101_000_0_000001000101;
      patterns[553] = 29'b0_000001000101_001_0_000101000001;
      patterns[554] = 29'b0_000001000101_010_0_000010001010;
      patterns[555] = 29'b0_000001000101_011_0_000100010100;
      patterns[556] = 29'b0_000001000101_100_1_000000100010;
      patterns[557] = 29'b0_000001000101_101_0_100000010001;
      patterns[558] = 29'b0_000001000101_110_0_000001000101;
      patterns[559] = 29'b0_000001000101_111_0_000001000101;
      patterns[560] = 29'b0_000001000110_000_0_000001000110;
      patterns[561] = 29'b0_000001000110_001_0_000110000001;
      patterns[562] = 29'b0_000001000110_010_0_000010001100;
      patterns[563] = 29'b0_000001000110_011_0_000100011000;
      patterns[564] = 29'b0_000001000110_100_0_000000100011;
      patterns[565] = 29'b0_000001000110_101_1_000000010001;
      patterns[566] = 29'b0_000001000110_110_0_000001000110;
      patterns[567] = 29'b0_000001000110_111_0_000001000110;
      patterns[568] = 29'b0_000001000111_000_0_000001000111;
      patterns[569] = 29'b0_000001000111_001_0_000111000001;
      patterns[570] = 29'b0_000001000111_010_0_000010001110;
      patterns[571] = 29'b0_000001000111_011_0_000100011100;
      patterns[572] = 29'b0_000001000111_100_1_000000100011;
      patterns[573] = 29'b0_000001000111_101_1_100000010001;
      patterns[574] = 29'b0_000001000111_110_0_000001000111;
      patterns[575] = 29'b0_000001000111_111_0_000001000111;
      patterns[576] = 29'b0_000001001000_000_0_000001001000;
      patterns[577] = 29'b0_000001001000_001_0_001000000001;
      patterns[578] = 29'b0_000001001000_010_0_000010010000;
      patterns[579] = 29'b0_000001001000_011_0_000100100000;
      patterns[580] = 29'b0_000001001000_100_0_000000100100;
      patterns[581] = 29'b0_000001001000_101_0_000000010010;
      patterns[582] = 29'b0_000001001000_110_0_000001001000;
      patterns[583] = 29'b0_000001001000_111_0_000001001000;
      patterns[584] = 29'b0_000001001001_000_0_000001001001;
      patterns[585] = 29'b0_000001001001_001_0_001001000001;
      patterns[586] = 29'b0_000001001001_010_0_000010010010;
      patterns[587] = 29'b0_000001001001_011_0_000100100100;
      patterns[588] = 29'b0_000001001001_100_1_000000100100;
      patterns[589] = 29'b0_000001001001_101_0_100000010010;
      patterns[590] = 29'b0_000001001001_110_0_000001001001;
      patterns[591] = 29'b0_000001001001_111_0_000001001001;
      patterns[592] = 29'b0_000001001010_000_0_000001001010;
      patterns[593] = 29'b0_000001001010_001_0_001010000001;
      patterns[594] = 29'b0_000001001010_010_0_000010010100;
      patterns[595] = 29'b0_000001001010_011_0_000100101000;
      patterns[596] = 29'b0_000001001010_100_0_000000100101;
      patterns[597] = 29'b0_000001001010_101_1_000000010010;
      patterns[598] = 29'b0_000001001010_110_0_000001001010;
      patterns[599] = 29'b0_000001001010_111_0_000001001010;
      patterns[600] = 29'b0_000001001011_000_0_000001001011;
      patterns[601] = 29'b0_000001001011_001_0_001011000001;
      patterns[602] = 29'b0_000001001011_010_0_000010010110;
      patterns[603] = 29'b0_000001001011_011_0_000100101100;
      patterns[604] = 29'b0_000001001011_100_1_000000100101;
      patterns[605] = 29'b0_000001001011_101_1_100000010010;
      patterns[606] = 29'b0_000001001011_110_0_000001001011;
      patterns[607] = 29'b0_000001001011_111_0_000001001011;
      patterns[608] = 29'b0_000001001100_000_0_000001001100;
      patterns[609] = 29'b0_000001001100_001_0_001100000001;
      patterns[610] = 29'b0_000001001100_010_0_000010011000;
      patterns[611] = 29'b0_000001001100_011_0_000100110000;
      patterns[612] = 29'b0_000001001100_100_0_000000100110;
      patterns[613] = 29'b0_000001001100_101_0_000000010011;
      patterns[614] = 29'b0_000001001100_110_0_000001001100;
      patterns[615] = 29'b0_000001001100_111_0_000001001100;
      patterns[616] = 29'b0_000001001101_000_0_000001001101;
      patterns[617] = 29'b0_000001001101_001_0_001101000001;
      patterns[618] = 29'b0_000001001101_010_0_000010011010;
      patterns[619] = 29'b0_000001001101_011_0_000100110100;
      patterns[620] = 29'b0_000001001101_100_1_000000100110;
      patterns[621] = 29'b0_000001001101_101_0_100000010011;
      patterns[622] = 29'b0_000001001101_110_0_000001001101;
      patterns[623] = 29'b0_000001001101_111_0_000001001101;
      patterns[624] = 29'b0_000001001110_000_0_000001001110;
      patterns[625] = 29'b0_000001001110_001_0_001110000001;
      patterns[626] = 29'b0_000001001110_010_0_000010011100;
      patterns[627] = 29'b0_000001001110_011_0_000100111000;
      patterns[628] = 29'b0_000001001110_100_0_000000100111;
      patterns[629] = 29'b0_000001001110_101_1_000000010011;
      patterns[630] = 29'b0_000001001110_110_0_000001001110;
      patterns[631] = 29'b0_000001001110_111_0_000001001110;
      patterns[632] = 29'b0_000001001111_000_0_000001001111;
      patterns[633] = 29'b0_000001001111_001_0_001111000001;
      patterns[634] = 29'b0_000001001111_010_0_000010011110;
      patterns[635] = 29'b0_000001001111_011_0_000100111100;
      patterns[636] = 29'b0_000001001111_100_1_000000100111;
      patterns[637] = 29'b0_000001001111_101_1_100000010011;
      patterns[638] = 29'b0_000001001111_110_0_000001001111;
      patterns[639] = 29'b0_000001001111_111_0_000001001111;
      patterns[640] = 29'b0_000001010000_000_0_000001010000;
      patterns[641] = 29'b0_000001010000_001_0_010000000001;
      patterns[642] = 29'b0_000001010000_010_0_000010100000;
      patterns[643] = 29'b0_000001010000_011_0_000101000000;
      patterns[644] = 29'b0_000001010000_100_0_000000101000;
      patterns[645] = 29'b0_000001010000_101_0_000000010100;
      patterns[646] = 29'b0_000001010000_110_0_000001010000;
      patterns[647] = 29'b0_000001010000_111_0_000001010000;
      patterns[648] = 29'b0_000001010001_000_0_000001010001;
      patterns[649] = 29'b0_000001010001_001_0_010001000001;
      patterns[650] = 29'b0_000001010001_010_0_000010100010;
      patterns[651] = 29'b0_000001010001_011_0_000101000100;
      patterns[652] = 29'b0_000001010001_100_1_000000101000;
      patterns[653] = 29'b0_000001010001_101_0_100000010100;
      patterns[654] = 29'b0_000001010001_110_0_000001010001;
      patterns[655] = 29'b0_000001010001_111_0_000001010001;
      patterns[656] = 29'b0_000001010010_000_0_000001010010;
      patterns[657] = 29'b0_000001010010_001_0_010010000001;
      patterns[658] = 29'b0_000001010010_010_0_000010100100;
      patterns[659] = 29'b0_000001010010_011_0_000101001000;
      patterns[660] = 29'b0_000001010010_100_0_000000101001;
      patterns[661] = 29'b0_000001010010_101_1_000000010100;
      patterns[662] = 29'b0_000001010010_110_0_000001010010;
      patterns[663] = 29'b0_000001010010_111_0_000001010010;
      patterns[664] = 29'b0_000001010011_000_0_000001010011;
      patterns[665] = 29'b0_000001010011_001_0_010011000001;
      patterns[666] = 29'b0_000001010011_010_0_000010100110;
      patterns[667] = 29'b0_000001010011_011_0_000101001100;
      patterns[668] = 29'b0_000001010011_100_1_000000101001;
      patterns[669] = 29'b0_000001010011_101_1_100000010100;
      patterns[670] = 29'b0_000001010011_110_0_000001010011;
      patterns[671] = 29'b0_000001010011_111_0_000001010011;
      patterns[672] = 29'b0_000001010100_000_0_000001010100;
      patterns[673] = 29'b0_000001010100_001_0_010100000001;
      patterns[674] = 29'b0_000001010100_010_0_000010101000;
      patterns[675] = 29'b0_000001010100_011_0_000101010000;
      patterns[676] = 29'b0_000001010100_100_0_000000101010;
      patterns[677] = 29'b0_000001010100_101_0_000000010101;
      patterns[678] = 29'b0_000001010100_110_0_000001010100;
      patterns[679] = 29'b0_000001010100_111_0_000001010100;
      patterns[680] = 29'b0_000001010101_000_0_000001010101;
      patterns[681] = 29'b0_000001010101_001_0_010101000001;
      patterns[682] = 29'b0_000001010101_010_0_000010101010;
      patterns[683] = 29'b0_000001010101_011_0_000101010100;
      patterns[684] = 29'b0_000001010101_100_1_000000101010;
      patterns[685] = 29'b0_000001010101_101_0_100000010101;
      patterns[686] = 29'b0_000001010101_110_0_000001010101;
      patterns[687] = 29'b0_000001010101_111_0_000001010101;
      patterns[688] = 29'b0_000001010110_000_0_000001010110;
      patterns[689] = 29'b0_000001010110_001_0_010110000001;
      patterns[690] = 29'b0_000001010110_010_0_000010101100;
      patterns[691] = 29'b0_000001010110_011_0_000101011000;
      patterns[692] = 29'b0_000001010110_100_0_000000101011;
      patterns[693] = 29'b0_000001010110_101_1_000000010101;
      patterns[694] = 29'b0_000001010110_110_0_000001010110;
      patterns[695] = 29'b0_000001010110_111_0_000001010110;
      patterns[696] = 29'b0_000001010111_000_0_000001010111;
      patterns[697] = 29'b0_000001010111_001_0_010111000001;
      patterns[698] = 29'b0_000001010111_010_0_000010101110;
      patterns[699] = 29'b0_000001010111_011_0_000101011100;
      patterns[700] = 29'b0_000001010111_100_1_000000101011;
      patterns[701] = 29'b0_000001010111_101_1_100000010101;
      patterns[702] = 29'b0_000001010111_110_0_000001010111;
      patterns[703] = 29'b0_000001010111_111_0_000001010111;
      patterns[704] = 29'b0_000001011000_000_0_000001011000;
      patterns[705] = 29'b0_000001011000_001_0_011000000001;
      patterns[706] = 29'b0_000001011000_010_0_000010110000;
      patterns[707] = 29'b0_000001011000_011_0_000101100000;
      patterns[708] = 29'b0_000001011000_100_0_000000101100;
      patterns[709] = 29'b0_000001011000_101_0_000000010110;
      patterns[710] = 29'b0_000001011000_110_0_000001011000;
      patterns[711] = 29'b0_000001011000_111_0_000001011000;
      patterns[712] = 29'b0_000001011001_000_0_000001011001;
      patterns[713] = 29'b0_000001011001_001_0_011001000001;
      patterns[714] = 29'b0_000001011001_010_0_000010110010;
      patterns[715] = 29'b0_000001011001_011_0_000101100100;
      patterns[716] = 29'b0_000001011001_100_1_000000101100;
      patterns[717] = 29'b0_000001011001_101_0_100000010110;
      patterns[718] = 29'b0_000001011001_110_0_000001011001;
      patterns[719] = 29'b0_000001011001_111_0_000001011001;
      patterns[720] = 29'b0_000001011010_000_0_000001011010;
      patterns[721] = 29'b0_000001011010_001_0_011010000001;
      patterns[722] = 29'b0_000001011010_010_0_000010110100;
      patterns[723] = 29'b0_000001011010_011_0_000101101000;
      patterns[724] = 29'b0_000001011010_100_0_000000101101;
      patterns[725] = 29'b0_000001011010_101_1_000000010110;
      patterns[726] = 29'b0_000001011010_110_0_000001011010;
      patterns[727] = 29'b0_000001011010_111_0_000001011010;
      patterns[728] = 29'b0_000001011011_000_0_000001011011;
      patterns[729] = 29'b0_000001011011_001_0_011011000001;
      patterns[730] = 29'b0_000001011011_010_0_000010110110;
      patterns[731] = 29'b0_000001011011_011_0_000101101100;
      patterns[732] = 29'b0_000001011011_100_1_000000101101;
      patterns[733] = 29'b0_000001011011_101_1_100000010110;
      patterns[734] = 29'b0_000001011011_110_0_000001011011;
      patterns[735] = 29'b0_000001011011_111_0_000001011011;
      patterns[736] = 29'b0_000001011100_000_0_000001011100;
      patterns[737] = 29'b0_000001011100_001_0_011100000001;
      patterns[738] = 29'b0_000001011100_010_0_000010111000;
      patterns[739] = 29'b0_000001011100_011_0_000101110000;
      patterns[740] = 29'b0_000001011100_100_0_000000101110;
      patterns[741] = 29'b0_000001011100_101_0_000000010111;
      patterns[742] = 29'b0_000001011100_110_0_000001011100;
      patterns[743] = 29'b0_000001011100_111_0_000001011100;
      patterns[744] = 29'b0_000001011101_000_0_000001011101;
      patterns[745] = 29'b0_000001011101_001_0_011101000001;
      patterns[746] = 29'b0_000001011101_010_0_000010111010;
      patterns[747] = 29'b0_000001011101_011_0_000101110100;
      patterns[748] = 29'b0_000001011101_100_1_000000101110;
      patterns[749] = 29'b0_000001011101_101_0_100000010111;
      patterns[750] = 29'b0_000001011101_110_0_000001011101;
      patterns[751] = 29'b0_000001011101_111_0_000001011101;
      patterns[752] = 29'b0_000001011110_000_0_000001011110;
      patterns[753] = 29'b0_000001011110_001_0_011110000001;
      patterns[754] = 29'b0_000001011110_010_0_000010111100;
      patterns[755] = 29'b0_000001011110_011_0_000101111000;
      patterns[756] = 29'b0_000001011110_100_0_000000101111;
      patterns[757] = 29'b0_000001011110_101_1_000000010111;
      patterns[758] = 29'b0_000001011110_110_0_000001011110;
      patterns[759] = 29'b0_000001011110_111_0_000001011110;
      patterns[760] = 29'b0_000001011111_000_0_000001011111;
      patterns[761] = 29'b0_000001011111_001_0_011111000001;
      patterns[762] = 29'b0_000001011111_010_0_000010111110;
      patterns[763] = 29'b0_000001011111_011_0_000101111100;
      patterns[764] = 29'b0_000001011111_100_1_000000101111;
      patterns[765] = 29'b0_000001011111_101_1_100000010111;
      patterns[766] = 29'b0_000001011111_110_0_000001011111;
      patterns[767] = 29'b0_000001011111_111_0_000001011111;
      patterns[768] = 29'b0_000001100000_000_0_000001100000;
      patterns[769] = 29'b0_000001100000_001_0_100000000001;
      patterns[770] = 29'b0_000001100000_010_0_000011000000;
      patterns[771] = 29'b0_000001100000_011_0_000110000000;
      patterns[772] = 29'b0_000001100000_100_0_000000110000;
      patterns[773] = 29'b0_000001100000_101_0_000000011000;
      patterns[774] = 29'b0_000001100000_110_0_000001100000;
      patterns[775] = 29'b0_000001100000_111_0_000001100000;
      patterns[776] = 29'b0_000001100001_000_0_000001100001;
      patterns[777] = 29'b0_000001100001_001_0_100001000001;
      patterns[778] = 29'b0_000001100001_010_0_000011000010;
      patterns[779] = 29'b0_000001100001_011_0_000110000100;
      patterns[780] = 29'b0_000001100001_100_1_000000110000;
      patterns[781] = 29'b0_000001100001_101_0_100000011000;
      patterns[782] = 29'b0_000001100001_110_0_000001100001;
      patterns[783] = 29'b0_000001100001_111_0_000001100001;
      patterns[784] = 29'b0_000001100010_000_0_000001100010;
      patterns[785] = 29'b0_000001100010_001_0_100010000001;
      patterns[786] = 29'b0_000001100010_010_0_000011000100;
      patterns[787] = 29'b0_000001100010_011_0_000110001000;
      patterns[788] = 29'b0_000001100010_100_0_000000110001;
      patterns[789] = 29'b0_000001100010_101_1_000000011000;
      patterns[790] = 29'b0_000001100010_110_0_000001100010;
      patterns[791] = 29'b0_000001100010_111_0_000001100010;
      patterns[792] = 29'b0_000001100011_000_0_000001100011;
      patterns[793] = 29'b0_000001100011_001_0_100011000001;
      patterns[794] = 29'b0_000001100011_010_0_000011000110;
      patterns[795] = 29'b0_000001100011_011_0_000110001100;
      patterns[796] = 29'b0_000001100011_100_1_000000110001;
      patterns[797] = 29'b0_000001100011_101_1_100000011000;
      patterns[798] = 29'b0_000001100011_110_0_000001100011;
      patterns[799] = 29'b0_000001100011_111_0_000001100011;
      patterns[800] = 29'b0_000001100100_000_0_000001100100;
      patterns[801] = 29'b0_000001100100_001_0_100100000001;
      patterns[802] = 29'b0_000001100100_010_0_000011001000;
      patterns[803] = 29'b0_000001100100_011_0_000110010000;
      patterns[804] = 29'b0_000001100100_100_0_000000110010;
      patterns[805] = 29'b0_000001100100_101_0_000000011001;
      patterns[806] = 29'b0_000001100100_110_0_000001100100;
      patterns[807] = 29'b0_000001100100_111_0_000001100100;
      patterns[808] = 29'b0_000001100101_000_0_000001100101;
      patterns[809] = 29'b0_000001100101_001_0_100101000001;
      patterns[810] = 29'b0_000001100101_010_0_000011001010;
      patterns[811] = 29'b0_000001100101_011_0_000110010100;
      patterns[812] = 29'b0_000001100101_100_1_000000110010;
      patterns[813] = 29'b0_000001100101_101_0_100000011001;
      patterns[814] = 29'b0_000001100101_110_0_000001100101;
      patterns[815] = 29'b0_000001100101_111_0_000001100101;
      patterns[816] = 29'b0_000001100110_000_0_000001100110;
      patterns[817] = 29'b0_000001100110_001_0_100110000001;
      patterns[818] = 29'b0_000001100110_010_0_000011001100;
      patterns[819] = 29'b0_000001100110_011_0_000110011000;
      patterns[820] = 29'b0_000001100110_100_0_000000110011;
      patterns[821] = 29'b0_000001100110_101_1_000000011001;
      patterns[822] = 29'b0_000001100110_110_0_000001100110;
      patterns[823] = 29'b0_000001100110_111_0_000001100110;
      patterns[824] = 29'b0_000001100111_000_0_000001100111;
      patterns[825] = 29'b0_000001100111_001_0_100111000001;
      patterns[826] = 29'b0_000001100111_010_0_000011001110;
      patterns[827] = 29'b0_000001100111_011_0_000110011100;
      patterns[828] = 29'b0_000001100111_100_1_000000110011;
      patterns[829] = 29'b0_000001100111_101_1_100000011001;
      patterns[830] = 29'b0_000001100111_110_0_000001100111;
      patterns[831] = 29'b0_000001100111_111_0_000001100111;
      patterns[832] = 29'b0_000001101000_000_0_000001101000;
      patterns[833] = 29'b0_000001101000_001_0_101000000001;
      patterns[834] = 29'b0_000001101000_010_0_000011010000;
      patterns[835] = 29'b0_000001101000_011_0_000110100000;
      patterns[836] = 29'b0_000001101000_100_0_000000110100;
      patterns[837] = 29'b0_000001101000_101_0_000000011010;
      patterns[838] = 29'b0_000001101000_110_0_000001101000;
      patterns[839] = 29'b0_000001101000_111_0_000001101000;
      patterns[840] = 29'b0_000001101001_000_0_000001101001;
      patterns[841] = 29'b0_000001101001_001_0_101001000001;
      patterns[842] = 29'b0_000001101001_010_0_000011010010;
      patterns[843] = 29'b0_000001101001_011_0_000110100100;
      patterns[844] = 29'b0_000001101001_100_1_000000110100;
      patterns[845] = 29'b0_000001101001_101_0_100000011010;
      patterns[846] = 29'b0_000001101001_110_0_000001101001;
      patterns[847] = 29'b0_000001101001_111_0_000001101001;
      patterns[848] = 29'b0_000001101010_000_0_000001101010;
      patterns[849] = 29'b0_000001101010_001_0_101010000001;
      patterns[850] = 29'b0_000001101010_010_0_000011010100;
      patterns[851] = 29'b0_000001101010_011_0_000110101000;
      patterns[852] = 29'b0_000001101010_100_0_000000110101;
      patterns[853] = 29'b0_000001101010_101_1_000000011010;
      patterns[854] = 29'b0_000001101010_110_0_000001101010;
      patterns[855] = 29'b0_000001101010_111_0_000001101010;
      patterns[856] = 29'b0_000001101011_000_0_000001101011;
      patterns[857] = 29'b0_000001101011_001_0_101011000001;
      patterns[858] = 29'b0_000001101011_010_0_000011010110;
      patterns[859] = 29'b0_000001101011_011_0_000110101100;
      patterns[860] = 29'b0_000001101011_100_1_000000110101;
      patterns[861] = 29'b0_000001101011_101_1_100000011010;
      patterns[862] = 29'b0_000001101011_110_0_000001101011;
      patterns[863] = 29'b0_000001101011_111_0_000001101011;
      patterns[864] = 29'b0_000001101100_000_0_000001101100;
      patterns[865] = 29'b0_000001101100_001_0_101100000001;
      patterns[866] = 29'b0_000001101100_010_0_000011011000;
      patterns[867] = 29'b0_000001101100_011_0_000110110000;
      patterns[868] = 29'b0_000001101100_100_0_000000110110;
      patterns[869] = 29'b0_000001101100_101_0_000000011011;
      patterns[870] = 29'b0_000001101100_110_0_000001101100;
      patterns[871] = 29'b0_000001101100_111_0_000001101100;
      patterns[872] = 29'b0_000001101101_000_0_000001101101;
      patterns[873] = 29'b0_000001101101_001_0_101101000001;
      patterns[874] = 29'b0_000001101101_010_0_000011011010;
      patterns[875] = 29'b0_000001101101_011_0_000110110100;
      patterns[876] = 29'b0_000001101101_100_1_000000110110;
      patterns[877] = 29'b0_000001101101_101_0_100000011011;
      patterns[878] = 29'b0_000001101101_110_0_000001101101;
      patterns[879] = 29'b0_000001101101_111_0_000001101101;
      patterns[880] = 29'b0_000001101110_000_0_000001101110;
      patterns[881] = 29'b0_000001101110_001_0_101110000001;
      patterns[882] = 29'b0_000001101110_010_0_000011011100;
      patterns[883] = 29'b0_000001101110_011_0_000110111000;
      patterns[884] = 29'b0_000001101110_100_0_000000110111;
      patterns[885] = 29'b0_000001101110_101_1_000000011011;
      patterns[886] = 29'b0_000001101110_110_0_000001101110;
      patterns[887] = 29'b0_000001101110_111_0_000001101110;
      patterns[888] = 29'b0_000001101111_000_0_000001101111;
      patterns[889] = 29'b0_000001101111_001_0_101111000001;
      patterns[890] = 29'b0_000001101111_010_0_000011011110;
      patterns[891] = 29'b0_000001101111_011_0_000110111100;
      patterns[892] = 29'b0_000001101111_100_1_000000110111;
      patterns[893] = 29'b0_000001101111_101_1_100000011011;
      patterns[894] = 29'b0_000001101111_110_0_000001101111;
      patterns[895] = 29'b0_000001101111_111_0_000001101111;
      patterns[896] = 29'b0_000001110000_000_0_000001110000;
      patterns[897] = 29'b0_000001110000_001_0_110000000001;
      patterns[898] = 29'b0_000001110000_010_0_000011100000;
      patterns[899] = 29'b0_000001110000_011_0_000111000000;
      patterns[900] = 29'b0_000001110000_100_0_000000111000;
      patterns[901] = 29'b0_000001110000_101_0_000000011100;
      patterns[902] = 29'b0_000001110000_110_0_000001110000;
      patterns[903] = 29'b0_000001110000_111_0_000001110000;
      patterns[904] = 29'b0_000001110001_000_0_000001110001;
      patterns[905] = 29'b0_000001110001_001_0_110001000001;
      patterns[906] = 29'b0_000001110001_010_0_000011100010;
      patterns[907] = 29'b0_000001110001_011_0_000111000100;
      patterns[908] = 29'b0_000001110001_100_1_000000111000;
      patterns[909] = 29'b0_000001110001_101_0_100000011100;
      patterns[910] = 29'b0_000001110001_110_0_000001110001;
      patterns[911] = 29'b0_000001110001_111_0_000001110001;
      patterns[912] = 29'b0_000001110010_000_0_000001110010;
      patterns[913] = 29'b0_000001110010_001_0_110010000001;
      patterns[914] = 29'b0_000001110010_010_0_000011100100;
      patterns[915] = 29'b0_000001110010_011_0_000111001000;
      patterns[916] = 29'b0_000001110010_100_0_000000111001;
      patterns[917] = 29'b0_000001110010_101_1_000000011100;
      patterns[918] = 29'b0_000001110010_110_0_000001110010;
      patterns[919] = 29'b0_000001110010_111_0_000001110010;
      patterns[920] = 29'b0_000001110011_000_0_000001110011;
      patterns[921] = 29'b0_000001110011_001_0_110011000001;
      patterns[922] = 29'b0_000001110011_010_0_000011100110;
      patterns[923] = 29'b0_000001110011_011_0_000111001100;
      patterns[924] = 29'b0_000001110011_100_1_000000111001;
      patterns[925] = 29'b0_000001110011_101_1_100000011100;
      patterns[926] = 29'b0_000001110011_110_0_000001110011;
      patterns[927] = 29'b0_000001110011_111_0_000001110011;
      patterns[928] = 29'b0_000001110100_000_0_000001110100;
      patterns[929] = 29'b0_000001110100_001_0_110100000001;
      patterns[930] = 29'b0_000001110100_010_0_000011101000;
      patterns[931] = 29'b0_000001110100_011_0_000111010000;
      patterns[932] = 29'b0_000001110100_100_0_000000111010;
      patterns[933] = 29'b0_000001110100_101_0_000000011101;
      patterns[934] = 29'b0_000001110100_110_0_000001110100;
      patterns[935] = 29'b0_000001110100_111_0_000001110100;
      patterns[936] = 29'b0_000001110101_000_0_000001110101;
      patterns[937] = 29'b0_000001110101_001_0_110101000001;
      patterns[938] = 29'b0_000001110101_010_0_000011101010;
      patterns[939] = 29'b0_000001110101_011_0_000111010100;
      patterns[940] = 29'b0_000001110101_100_1_000000111010;
      patterns[941] = 29'b0_000001110101_101_0_100000011101;
      patterns[942] = 29'b0_000001110101_110_0_000001110101;
      patterns[943] = 29'b0_000001110101_111_0_000001110101;
      patterns[944] = 29'b0_000001110110_000_0_000001110110;
      patterns[945] = 29'b0_000001110110_001_0_110110000001;
      patterns[946] = 29'b0_000001110110_010_0_000011101100;
      patterns[947] = 29'b0_000001110110_011_0_000111011000;
      patterns[948] = 29'b0_000001110110_100_0_000000111011;
      patterns[949] = 29'b0_000001110110_101_1_000000011101;
      patterns[950] = 29'b0_000001110110_110_0_000001110110;
      patterns[951] = 29'b0_000001110110_111_0_000001110110;
      patterns[952] = 29'b0_000001110111_000_0_000001110111;
      patterns[953] = 29'b0_000001110111_001_0_110111000001;
      patterns[954] = 29'b0_000001110111_010_0_000011101110;
      patterns[955] = 29'b0_000001110111_011_0_000111011100;
      patterns[956] = 29'b0_000001110111_100_1_000000111011;
      patterns[957] = 29'b0_000001110111_101_1_100000011101;
      patterns[958] = 29'b0_000001110111_110_0_000001110111;
      patterns[959] = 29'b0_000001110111_111_0_000001110111;
      patterns[960] = 29'b0_000001111000_000_0_000001111000;
      patterns[961] = 29'b0_000001111000_001_0_111000000001;
      patterns[962] = 29'b0_000001111000_010_0_000011110000;
      patterns[963] = 29'b0_000001111000_011_0_000111100000;
      patterns[964] = 29'b0_000001111000_100_0_000000111100;
      patterns[965] = 29'b0_000001111000_101_0_000000011110;
      patterns[966] = 29'b0_000001111000_110_0_000001111000;
      patterns[967] = 29'b0_000001111000_111_0_000001111000;
      patterns[968] = 29'b0_000001111001_000_0_000001111001;
      patterns[969] = 29'b0_000001111001_001_0_111001000001;
      patterns[970] = 29'b0_000001111001_010_0_000011110010;
      patterns[971] = 29'b0_000001111001_011_0_000111100100;
      patterns[972] = 29'b0_000001111001_100_1_000000111100;
      patterns[973] = 29'b0_000001111001_101_0_100000011110;
      patterns[974] = 29'b0_000001111001_110_0_000001111001;
      patterns[975] = 29'b0_000001111001_111_0_000001111001;
      patterns[976] = 29'b0_000001111010_000_0_000001111010;
      patterns[977] = 29'b0_000001111010_001_0_111010000001;
      patterns[978] = 29'b0_000001111010_010_0_000011110100;
      patterns[979] = 29'b0_000001111010_011_0_000111101000;
      patterns[980] = 29'b0_000001111010_100_0_000000111101;
      patterns[981] = 29'b0_000001111010_101_1_000000011110;
      patterns[982] = 29'b0_000001111010_110_0_000001111010;
      patterns[983] = 29'b0_000001111010_111_0_000001111010;
      patterns[984] = 29'b0_000001111011_000_0_000001111011;
      patterns[985] = 29'b0_000001111011_001_0_111011000001;
      patterns[986] = 29'b0_000001111011_010_0_000011110110;
      patterns[987] = 29'b0_000001111011_011_0_000111101100;
      patterns[988] = 29'b0_000001111011_100_1_000000111101;
      patterns[989] = 29'b0_000001111011_101_1_100000011110;
      patterns[990] = 29'b0_000001111011_110_0_000001111011;
      patterns[991] = 29'b0_000001111011_111_0_000001111011;
      patterns[992] = 29'b0_000001111100_000_0_000001111100;
      patterns[993] = 29'b0_000001111100_001_0_111100000001;
      patterns[994] = 29'b0_000001111100_010_0_000011111000;
      patterns[995] = 29'b0_000001111100_011_0_000111110000;
      patterns[996] = 29'b0_000001111100_100_0_000000111110;
      patterns[997] = 29'b0_000001111100_101_0_000000011111;
      patterns[998] = 29'b0_000001111100_110_0_000001111100;
      patterns[999] = 29'b0_000001111100_111_0_000001111100;
      patterns[1000] = 29'b0_000001111101_000_0_000001111101;
      patterns[1001] = 29'b0_000001111101_001_0_111101000001;
      patterns[1002] = 29'b0_000001111101_010_0_000011111010;
      patterns[1003] = 29'b0_000001111101_011_0_000111110100;
      patterns[1004] = 29'b0_000001111101_100_1_000000111110;
      patterns[1005] = 29'b0_000001111101_101_0_100000011111;
      patterns[1006] = 29'b0_000001111101_110_0_000001111101;
      patterns[1007] = 29'b0_000001111101_111_0_000001111101;
      patterns[1008] = 29'b0_000001111110_000_0_000001111110;
      patterns[1009] = 29'b0_000001111110_001_0_111110000001;
      patterns[1010] = 29'b0_000001111110_010_0_000011111100;
      patterns[1011] = 29'b0_000001111110_011_0_000111111000;
      patterns[1012] = 29'b0_000001111110_100_0_000000111111;
      patterns[1013] = 29'b0_000001111110_101_1_000000011111;
      patterns[1014] = 29'b0_000001111110_110_0_000001111110;
      patterns[1015] = 29'b0_000001111110_111_0_000001111110;
      patterns[1016] = 29'b0_000001111111_000_0_000001111111;
      patterns[1017] = 29'b0_000001111111_001_0_111111000001;
      patterns[1018] = 29'b0_000001111111_010_0_000011111110;
      patterns[1019] = 29'b0_000001111111_011_0_000111111100;
      patterns[1020] = 29'b0_000001111111_100_1_000000111111;
      patterns[1021] = 29'b0_000001111111_101_1_100000011111;
      patterns[1022] = 29'b0_000001111111_110_0_000001111111;
      patterns[1023] = 29'b0_000001111111_111_0_000001111111;
      patterns[1024] = 29'b0_000010000000_000_0_000010000000;
      patterns[1025] = 29'b0_000010000000_001_0_000000000010;
      patterns[1026] = 29'b0_000010000000_010_0_000100000000;
      patterns[1027] = 29'b0_000010000000_011_0_001000000000;
      patterns[1028] = 29'b0_000010000000_100_0_000001000000;
      patterns[1029] = 29'b0_000010000000_101_0_000000100000;
      patterns[1030] = 29'b0_000010000000_110_0_000010000000;
      patterns[1031] = 29'b0_000010000000_111_0_000010000000;
      patterns[1032] = 29'b0_000010000001_000_0_000010000001;
      patterns[1033] = 29'b0_000010000001_001_0_000001000010;
      patterns[1034] = 29'b0_000010000001_010_0_000100000010;
      patterns[1035] = 29'b0_000010000001_011_0_001000000100;
      patterns[1036] = 29'b0_000010000001_100_1_000001000000;
      patterns[1037] = 29'b0_000010000001_101_0_100000100000;
      patterns[1038] = 29'b0_000010000001_110_0_000010000001;
      patterns[1039] = 29'b0_000010000001_111_0_000010000001;
      patterns[1040] = 29'b0_000010000010_000_0_000010000010;
      patterns[1041] = 29'b0_000010000010_001_0_000010000010;
      patterns[1042] = 29'b0_000010000010_010_0_000100000100;
      patterns[1043] = 29'b0_000010000010_011_0_001000001000;
      patterns[1044] = 29'b0_000010000010_100_0_000001000001;
      patterns[1045] = 29'b0_000010000010_101_1_000000100000;
      patterns[1046] = 29'b0_000010000010_110_0_000010000010;
      patterns[1047] = 29'b0_000010000010_111_0_000010000010;
      patterns[1048] = 29'b0_000010000011_000_0_000010000011;
      patterns[1049] = 29'b0_000010000011_001_0_000011000010;
      patterns[1050] = 29'b0_000010000011_010_0_000100000110;
      patterns[1051] = 29'b0_000010000011_011_0_001000001100;
      patterns[1052] = 29'b0_000010000011_100_1_000001000001;
      patterns[1053] = 29'b0_000010000011_101_1_100000100000;
      patterns[1054] = 29'b0_000010000011_110_0_000010000011;
      patterns[1055] = 29'b0_000010000011_111_0_000010000011;
      patterns[1056] = 29'b0_000010000100_000_0_000010000100;
      patterns[1057] = 29'b0_000010000100_001_0_000100000010;
      patterns[1058] = 29'b0_000010000100_010_0_000100001000;
      patterns[1059] = 29'b0_000010000100_011_0_001000010000;
      patterns[1060] = 29'b0_000010000100_100_0_000001000010;
      patterns[1061] = 29'b0_000010000100_101_0_000000100001;
      patterns[1062] = 29'b0_000010000100_110_0_000010000100;
      patterns[1063] = 29'b0_000010000100_111_0_000010000100;
      patterns[1064] = 29'b0_000010000101_000_0_000010000101;
      patterns[1065] = 29'b0_000010000101_001_0_000101000010;
      patterns[1066] = 29'b0_000010000101_010_0_000100001010;
      patterns[1067] = 29'b0_000010000101_011_0_001000010100;
      patterns[1068] = 29'b0_000010000101_100_1_000001000010;
      patterns[1069] = 29'b0_000010000101_101_0_100000100001;
      patterns[1070] = 29'b0_000010000101_110_0_000010000101;
      patterns[1071] = 29'b0_000010000101_111_0_000010000101;
      patterns[1072] = 29'b0_000010000110_000_0_000010000110;
      patterns[1073] = 29'b0_000010000110_001_0_000110000010;
      patterns[1074] = 29'b0_000010000110_010_0_000100001100;
      patterns[1075] = 29'b0_000010000110_011_0_001000011000;
      patterns[1076] = 29'b0_000010000110_100_0_000001000011;
      patterns[1077] = 29'b0_000010000110_101_1_000000100001;
      patterns[1078] = 29'b0_000010000110_110_0_000010000110;
      patterns[1079] = 29'b0_000010000110_111_0_000010000110;
      patterns[1080] = 29'b0_000010000111_000_0_000010000111;
      patterns[1081] = 29'b0_000010000111_001_0_000111000010;
      patterns[1082] = 29'b0_000010000111_010_0_000100001110;
      patterns[1083] = 29'b0_000010000111_011_0_001000011100;
      patterns[1084] = 29'b0_000010000111_100_1_000001000011;
      patterns[1085] = 29'b0_000010000111_101_1_100000100001;
      patterns[1086] = 29'b0_000010000111_110_0_000010000111;
      patterns[1087] = 29'b0_000010000111_111_0_000010000111;
      patterns[1088] = 29'b0_000010001000_000_0_000010001000;
      patterns[1089] = 29'b0_000010001000_001_0_001000000010;
      patterns[1090] = 29'b0_000010001000_010_0_000100010000;
      patterns[1091] = 29'b0_000010001000_011_0_001000100000;
      patterns[1092] = 29'b0_000010001000_100_0_000001000100;
      patterns[1093] = 29'b0_000010001000_101_0_000000100010;
      patterns[1094] = 29'b0_000010001000_110_0_000010001000;
      patterns[1095] = 29'b0_000010001000_111_0_000010001000;
      patterns[1096] = 29'b0_000010001001_000_0_000010001001;
      patterns[1097] = 29'b0_000010001001_001_0_001001000010;
      patterns[1098] = 29'b0_000010001001_010_0_000100010010;
      patterns[1099] = 29'b0_000010001001_011_0_001000100100;
      patterns[1100] = 29'b0_000010001001_100_1_000001000100;
      patterns[1101] = 29'b0_000010001001_101_0_100000100010;
      patterns[1102] = 29'b0_000010001001_110_0_000010001001;
      patterns[1103] = 29'b0_000010001001_111_0_000010001001;
      patterns[1104] = 29'b0_000010001010_000_0_000010001010;
      patterns[1105] = 29'b0_000010001010_001_0_001010000010;
      patterns[1106] = 29'b0_000010001010_010_0_000100010100;
      patterns[1107] = 29'b0_000010001010_011_0_001000101000;
      patterns[1108] = 29'b0_000010001010_100_0_000001000101;
      patterns[1109] = 29'b0_000010001010_101_1_000000100010;
      patterns[1110] = 29'b0_000010001010_110_0_000010001010;
      patterns[1111] = 29'b0_000010001010_111_0_000010001010;
      patterns[1112] = 29'b0_000010001011_000_0_000010001011;
      patterns[1113] = 29'b0_000010001011_001_0_001011000010;
      patterns[1114] = 29'b0_000010001011_010_0_000100010110;
      patterns[1115] = 29'b0_000010001011_011_0_001000101100;
      patterns[1116] = 29'b0_000010001011_100_1_000001000101;
      patterns[1117] = 29'b0_000010001011_101_1_100000100010;
      patterns[1118] = 29'b0_000010001011_110_0_000010001011;
      patterns[1119] = 29'b0_000010001011_111_0_000010001011;
      patterns[1120] = 29'b0_000010001100_000_0_000010001100;
      patterns[1121] = 29'b0_000010001100_001_0_001100000010;
      patterns[1122] = 29'b0_000010001100_010_0_000100011000;
      patterns[1123] = 29'b0_000010001100_011_0_001000110000;
      patterns[1124] = 29'b0_000010001100_100_0_000001000110;
      patterns[1125] = 29'b0_000010001100_101_0_000000100011;
      patterns[1126] = 29'b0_000010001100_110_0_000010001100;
      patterns[1127] = 29'b0_000010001100_111_0_000010001100;
      patterns[1128] = 29'b0_000010001101_000_0_000010001101;
      patterns[1129] = 29'b0_000010001101_001_0_001101000010;
      patterns[1130] = 29'b0_000010001101_010_0_000100011010;
      patterns[1131] = 29'b0_000010001101_011_0_001000110100;
      patterns[1132] = 29'b0_000010001101_100_1_000001000110;
      patterns[1133] = 29'b0_000010001101_101_0_100000100011;
      patterns[1134] = 29'b0_000010001101_110_0_000010001101;
      patterns[1135] = 29'b0_000010001101_111_0_000010001101;
      patterns[1136] = 29'b0_000010001110_000_0_000010001110;
      patterns[1137] = 29'b0_000010001110_001_0_001110000010;
      patterns[1138] = 29'b0_000010001110_010_0_000100011100;
      patterns[1139] = 29'b0_000010001110_011_0_001000111000;
      patterns[1140] = 29'b0_000010001110_100_0_000001000111;
      patterns[1141] = 29'b0_000010001110_101_1_000000100011;
      patterns[1142] = 29'b0_000010001110_110_0_000010001110;
      patterns[1143] = 29'b0_000010001110_111_0_000010001110;
      patterns[1144] = 29'b0_000010001111_000_0_000010001111;
      patterns[1145] = 29'b0_000010001111_001_0_001111000010;
      patterns[1146] = 29'b0_000010001111_010_0_000100011110;
      patterns[1147] = 29'b0_000010001111_011_0_001000111100;
      patterns[1148] = 29'b0_000010001111_100_1_000001000111;
      patterns[1149] = 29'b0_000010001111_101_1_100000100011;
      patterns[1150] = 29'b0_000010001111_110_0_000010001111;
      patterns[1151] = 29'b0_000010001111_111_0_000010001111;
      patterns[1152] = 29'b0_000010010000_000_0_000010010000;
      patterns[1153] = 29'b0_000010010000_001_0_010000000010;
      patterns[1154] = 29'b0_000010010000_010_0_000100100000;
      patterns[1155] = 29'b0_000010010000_011_0_001001000000;
      patterns[1156] = 29'b0_000010010000_100_0_000001001000;
      patterns[1157] = 29'b0_000010010000_101_0_000000100100;
      patterns[1158] = 29'b0_000010010000_110_0_000010010000;
      patterns[1159] = 29'b0_000010010000_111_0_000010010000;
      patterns[1160] = 29'b0_000010010001_000_0_000010010001;
      patterns[1161] = 29'b0_000010010001_001_0_010001000010;
      patterns[1162] = 29'b0_000010010001_010_0_000100100010;
      patterns[1163] = 29'b0_000010010001_011_0_001001000100;
      patterns[1164] = 29'b0_000010010001_100_1_000001001000;
      patterns[1165] = 29'b0_000010010001_101_0_100000100100;
      patterns[1166] = 29'b0_000010010001_110_0_000010010001;
      patterns[1167] = 29'b0_000010010001_111_0_000010010001;
      patterns[1168] = 29'b0_000010010010_000_0_000010010010;
      patterns[1169] = 29'b0_000010010010_001_0_010010000010;
      patterns[1170] = 29'b0_000010010010_010_0_000100100100;
      patterns[1171] = 29'b0_000010010010_011_0_001001001000;
      patterns[1172] = 29'b0_000010010010_100_0_000001001001;
      patterns[1173] = 29'b0_000010010010_101_1_000000100100;
      patterns[1174] = 29'b0_000010010010_110_0_000010010010;
      patterns[1175] = 29'b0_000010010010_111_0_000010010010;
      patterns[1176] = 29'b0_000010010011_000_0_000010010011;
      patterns[1177] = 29'b0_000010010011_001_0_010011000010;
      patterns[1178] = 29'b0_000010010011_010_0_000100100110;
      patterns[1179] = 29'b0_000010010011_011_0_001001001100;
      patterns[1180] = 29'b0_000010010011_100_1_000001001001;
      patterns[1181] = 29'b0_000010010011_101_1_100000100100;
      patterns[1182] = 29'b0_000010010011_110_0_000010010011;
      patterns[1183] = 29'b0_000010010011_111_0_000010010011;
      patterns[1184] = 29'b0_000010010100_000_0_000010010100;
      patterns[1185] = 29'b0_000010010100_001_0_010100000010;
      patterns[1186] = 29'b0_000010010100_010_0_000100101000;
      patterns[1187] = 29'b0_000010010100_011_0_001001010000;
      patterns[1188] = 29'b0_000010010100_100_0_000001001010;
      patterns[1189] = 29'b0_000010010100_101_0_000000100101;
      patterns[1190] = 29'b0_000010010100_110_0_000010010100;
      patterns[1191] = 29'b0_000010010100_111_0_000010010100;
      patterns[1192] = 29'b0_000010010101_000_0_000010010101;
      patterns[1193] = 29'b0_000010010101_001_0_010101000010;
      patterns[1194] = 29'b0_000010010101_010_0_000100101010;
      patterns[1195] = 29'b0_000010010101_011_0_001001010100;
      patterns[1196] = 29'b0_000010010101_100_1_000001001010;
      patterns[1197] = 29'b0_000010010101_101_0_100000100101;
      patterns[1198] = 29'b0_000010010101_110_0_000010010101;
      patterns[1199] = 29'b0_000010010101_111_0_000010010101;
      patterns[1200] = 29'b0_000010010110_000_0_000010010110;
      patterns[1201] = 29'b0_000010010110_001_0_010110000010;
      patterns[1202] = 29'b0_000010010110_010_0_000100101100;
      patterns[1203] = 29'b0_000010010110_011_0_001001011000;
      patterns[1204] = 29'b0_000010010110_100_0_000001001011;
      patterns[1205] = 29'b0_000010010110_101_1_000000100101;
      patterns[1206] = 29'b0_000010010110_110_0_000010010110;
      patterns[1207] = 29'b0_000010010110_111_0_000010010110;
      patterns[1208] = 29'b0_000010010111_000_0_000010010111;
      patterns[1209] = 29'b0_000010010111_001_0_010111000010;
      patterns[1210] = 29'b0_000010010111_010_0_000100101110;
      patterns[1211] = 29'b0_000010010111_011_0_001001011100;
      patterns[1212] = 29'b0_000010010111_100_1_000001001011;
      patterns[1213] = 29'b0_000010010111_101_1_100000100101;
      patterns[1214] = 29'b0_000010010111_110_0_000010010111;
      patterns[1215] = 29'b0_000010010111_111_0_000010010111;
      patterns[1216] = 29'b0_000010011000_000_0_000010011000;
      patterns[1217] = 29'b0_000010011000_001_0_011000000010;
      patterns[1218] = 29'b0_000010011000_010_0_000100110000;
      patterns[1219] = 29'b0_000010011000_011_0_001001100000;
      patterns[1220] = 29'b0_000010011000_100_0_000001001100;
      patterns[1221] = 29'b0_000010011000_101_0_000000100110;
      patterns[1222] = 29'b0_000010011000_110_0_000010011000;
      patterns[1223] = 29'b0_000010011000_111_0_000010011000;
      patterns[1224] = 29'b0_000010011001_000_0_000010011001;
      patterns[1225] = 29'b0_000010011001_001_0_011001000010;
      patterns[1226] = 29'b0_000010011001_010_0_000100110010;
      patterns[1227] = 29'b0_000010011001_011_0_001001100100;
      patterns[1228] = 29'b0_000010011001_100_1_000001001100;
      patterns[1229] = 29'b0_000010011001_101_0_100000100110;
      patterns[1230] = 29'b0_000010011001_110_0_000010011001;
      patterns[1231] = 29'b0_000010011001_111_0_000010011001;
      patterns[1232] = 29'b0_000010011010_000_0_000010011010;
      patterns[1233] = 29'b0_000010011010_001_0_011010000010;
      patterns[1234] = 29'b0_000010011010_010_0_000100110100;
      patterns[1235] = 29'b0_000010011010_011_0_001001101000;
      patterns[1236] = 29'b0_000010011010_100_0_000001001101;
      patterns[1237] = 29'b0_000010011010_101_1_000000100110;
      patterns[1238] = 29'b0_000010011010_110_0_000010011010;
      patterns[1239] = 29'b0_000010011010_111_0_000010011010;
      patterns[1240] = 29'b0_000010011011_000_0_000010011011;
      patterns[1241] = 29'b0_000010011011_001_0_011011000010;
      patterns[1242] = 29'b0_000010011011_010_0_000100110110;
      patterns[1243] = 29'b0_000010011011_011_0_001001101100;
      patterns[1244] = 29'b0_000010011011_100_1_000001001101;
      patterns[1245] = 29'b0_000010011011_101_1_100000100110;
      patterns[1246] = 29'b0_000010011011_110_0_000010011011;
      patterns[1247] = 29'b0_000010011011_111_0_000010011011;
      patterns[1248] = 29'b0_000010011100_000_0_000010011100;
      patterns[1249] = 29'b0_000010011100_001_0_011100000010;
      patterns[1250] = 29'b0_000010011100_010_0_000100111000;
      patterns[1251] = 29'b0_000010011100_011_0_001001110000;
      patterns[1252] = 29'b0_000010011100_100_0_000001001110;
      patterns[1253] = 29'b0_000010011100_101_0_000000100111;
      patterns[1254] = 29'b0_000010011100_110_0_000010011100;
      patterns[1255] = 29'b0_000010011100_111_0_000010011100;
      patterns[1256] = 29'b0_000010011101_000_0_000010011101;
      patterns[1257] = 29'b0_000010011101_001_0_011101000010;
      patterns[1258] = 29'b0_000010011101_010_0_000100111010;
      patterns[1259] = 29'b0_000010011101_011_0_001001110100;
      patterns[1260] = 29'b0_000010011101_100_1_000001001110;
      patterns[1261] = 29'b0_000010011101_101_0_100000100111;
      patterns[1262] = 29'b0_000010011101_110_0_000010011101;
      patterns[1263] = 29'b0_000010011101_111_0_000010011101;
      patterns[1264] = 29'b0_000010011110_000_0_000010011110;
      patterns[1265] = 29'b0_000010011110_001_0_011110000010;
      patterns[1266] = 29'b0_000010011110_010_0_000100111100;
      patterns[1267] = 29'b0_000010011110_011_0_001001111000;
      patterns[1268] = 29'b0_000010011110_100_0_000001001111;
      patterns[1269] = 29'b0_000010011110_101_1_000000100111;
      patterns[1270] = 29'b0_000010011110_110_0_000010011110;
      patterns[1271] = 29'b0_000010011110_111_0_000010011110;
      patterns[1272] = 29'b0_000010011111_000_0_000010011111;
      patterns[1273] = 29'b0_000010011111_001_0_011111000010;
      patterns[1274] = 29'b0_000010011111_010_0_000100111110;
      patterns[1275] = 29'b0_000010011111_011_0_001001111100;
      patterns[1276] = 29'b0_000010011111_100_1_000001001111;
      patterns[1277] = 29'b0_000010011111_101_1_100000100111;
      patterns[1278] = 29'b0_000010011111_110_0_000010011111;
      patterns[1279] = 29'b0_000010011111_111_0_000010011111;
      patterns[1280] = 29'b0_000010100000_000_0_000010100000;
      patterns[1281] = 29'b0_000010100000_001_0_100000000010;
      patterns[1282] = 29'b0_000010100000_010_0_000101000000;
      patterns[1283] = 29'b0_000010100000_011_0_001010000000;
      patterns[1284] = 29'b0_000010100000_100_0_000001010000;
      patterns[1285] = 29'b0_000010100000_101_0_000000101000;
      patterns[1286] = 29'b0_000010100000_110_0_000010100000;
      patterns[1287] = 29'b0_000010100000_111_0_000010100000;
      patterns[1288] = 29'b0_000010100001_000_0_000010100001;
      patterns[1289] = 29'b0_000010100001_001_0_100001000010;
      patterns[1290] = 29'b0_000010100001_010_0_000101000010;
      patterns[1291] = 29'b0_000010100001_011_0_001010000100;
      patterns[1292] = 29'b0_000010100001_100_1_000001010000;
      patterns[1293] = 29'b0_000010100001_101_0_100000101000;
      patterns[1294] = 29'b0_000010100001_110_0_000010100001;
      patterns[1295] = 29'b0_000010100001_111_0_000010100001;
      patterns[1296] = 29'b0_000010100010_000_0_000010100010;
      patterns[1297] = 29'b0_000010100010_001_0_100010000010;
      patterns[1298] = 29'b0_000010100010_010_0_000101000100;
      patterns[1299] = 29'b0_000010100010_011_0_001010001000;
      patterns[1300] = 29'b0_000010100010_100_0_000001010001;
      patterns[1301] = 29'b0_000010100010_101_1_000000101000;
      patterns[1302] = 29'b0_000010100010_110_0_000010100010;
      patterns[1303] = 29'b0_000010100010_111_0_000010100010;
      patterns[1304] = 29'b0_000010100011_000_0_000010100011;
      patterns[1305] = 29'b0_000010100011_001_0_100011000010;
      patterns[1306] = 29'b0_000010100011_010_0_000101000110;
      patterns[1307] = 29'b0_000010100011_011_0_001010001100;
      patterns[1308] = 29'b0_000010100011_100_1_000001010001;
      patterns[1309] = 29'b0_000010100011_101_1_100000101000;
      patterns[1310] = 29'b0_000010100011_110_0_000010100011;
      patterns[1311] = 29'b0_000010100011_111_0_000010100011;
      patterns[1312] = 29'b0_000010100100_000_0_000010100100;
      patterns[1313] = 29'b0_000010100100_001_0_100100000010;
      patterns[1314] = 29'b0_000010100100_010_0_000101001000;
      patterns[1315] = 29'b0_000010100100_011_0_001010010000;
      patterns[1316] = 29'b0_000010100100_100_0_000001010010;
      patterns[1317] = 29'b0_000010100100_101_0_000000101001;
      patterns[1318] = 29'b0_000010100100_110_0_000010100100;
      patterns[1319] = 29'b0_000010100100_111_0_000010100100;
      patterns[1320] = 29'b0_000010100101_000_0_000010100101;
      patterns[1321] = 29'b0_000010100101_001_0_100101000010;
      patterns[1322] = 29'b0_000010100101_010_0_000101001010;
      patterns[1323] = 29'b0_000010100101_011_0_001010010100;
      patterns[1324] = 29'b0_000010100101_100_1_000001010010;
      patterns[1325] = 29'b0_000010100101_101_0_100000101001;
      patterns[1326] = 29'b0_000010100101_110_0_000010100101;
      patterns[1327] = 29'b0_000010100101_111_0_000010100101;
      patterns[1328] = 29'b0_000010100110_000_0_000010100110;
      patterns[1329] = 29'b0_000010100110_001_0_100110000010;
      patterns[1330] = 29'b0_000010100110_010_0_000101001100;
      patterns[1331] = 29'b0_000010100110_011_0_001010011000;
      patterns[1332] = 29'b0_000010100110_100_0_000001010011;
      patterns[1333] = 29'b0_000010100110_101_1_000000101001;
      patterns[1334] = 29'b0_000010100110_110_0_000010100110;
      patterns[1335] = 29'b0_000010100110_111_0_000010100110;
      patterns[1336] = 29'b0_000010100111_000_0_000010100111;
      patterns[1337] = 29'b0_000010100111_001_0_100111000010;
      patterns[1338] = 29'b0_000010100111_010_0_000101001110;
      patterns[1339] = 29'b0_000010100111_011_0_001010011100;
      patterns[1340] = 29'b0_000010100111_100_1_000001010011;
      patterns[1341] = 29'b0_000010100111_101_1_100000101001;
      patterns[1342] = 29'b0_000010100111_110_0_000010100111;
      patterns[1343] = 29'b0_000010100111_111_0_000010100111;
      patterns[1344] = 29'b0_000010101000_000_0_000010101000;
      patterns[1345] = 29'b0_000010101000_001_0_101000000010;
      patterns[1346] = 29'b0_000010101000_010_0_000101010000;
      patterns[1347] = 29'b0_000010101000_011_0_001010100000;
      patterns[1348] = 29'b0_000010101000_100_0_000001010100;
      patterns[1349] = 29'b0_000010101000_101_0_000000101010;
      patterns[1350] = 29'b0_000010101000_110_0_000010101000;
      patterns[1351] = 29'b0_000010101000_111_0_000010101000;
      patterns[1352] = 29'b0_000010101001_000_0_000010101001;
      patterns[1353] = 29'b0_000010101001_001_0_101001000010;
      patterns[1354] = 29'b0_000010101001_010_0_000101010010;
      patterns[1355] = 29'b0_000010101001_011_0_001010100100;
      patterns[1356] = 29'b0_000010101001_100_1_000001010100;
      patterns[1357] = 29'b0_000010101001_101_0_100000101010;
      patterns[1358] = 29'b0_000010101001_110_0_000010101001;
      patterns[1359] = 29'b0_000010101001_111_0_000010101001;
      patterns[1360] = 29'b0_000010101010_000_0_000010101010;
      patterns[1361] = 29'b0_000010101010_001_0_101010000010;
      patterns[1362] = 29'b0_000010101010_010_0_000101010100;
      patterns[1363] = 29'b0_000010101010_011_0_001010101000;
      patterns[1364] = 29'b0_000010101010_100_0_000001010101;
      patterns[1365] = 29'b0_000010101010_101_1_000000101010;
      patterns[1366] = 29'b0_000010101010_110_0_000010101010;
      patterns[1367] = 29'b0_000010101010_111_0_000010101010;
      patterns[1368] = 29'b0_000010101011_000_0_000010101011;
      patterns[1369] = 29'b0_000010101011_001_0_101011000010;
      patterns[1370] = 29'b0_000010101011_010_0_000101010110;
      patterns[1371] = 29'b0_000010101011_011_0_001010101100;
      patterns[1372] = 29'b0_000010101011_100_1_000001010101;
      patterns[1373] = 29'b0_000010101011_101_1_100000101010;
      patterns[1374] = 29'b0_000010101011_110_0_000010101011;
      patterns[1375] = 29'b0_000010101011_111_0_000010101011;
      patterns[1376] = 29'b0_000010101100_000_0_000010101100;
      patterns[1377] = 29'b0_000010101100_001_0_101100000010;
      patterns[1378] = 29'b0_000010101100_010_0_000101011000;
      patterns[1379] = 29'b0_000010101100_011_0_001010110000;
      patterns[1380] = 29'b0_000010101100_100_0_000001010110;
      patterns[1381] = 29'b0_000010101100_101_0_000000101011;
      patterns[1382] = 29'b0_000010101100_110_0_000010101100;
      patterns[1383] = 29'b0_000010101100_111_0_000010101100;
      patterns[1384] = 29'b0_000010101101_000_0_000010101101;
      patterns[1385] = 29'b0_000010101101_001_0_101101000010;
      patterns[1386] = 29'b0_000010101101_010_0_000101011010;
      patterns[1387] = 29'b0_000010101101_011_0_001010110100;
      patterns[1388] = 29'b0_000010101101_100_1_000001010110;
      patterns[1389] = 29'b0_000010101101_101_0_100000101011;
      patterns[1390] = 29'b0_000010101101_110_0_000010101101;
      patterns[1391] = 29'b0_000010101101_111_0_000010101101;
      patterns[1392] = 29'b0_000010101110_000_0_000010101110;
      patterns[1393] = 29'b0_000010101110_001_0_101110000010;
      patterns[1394] = 29'b0_000010101110_010_0_000101011100;
      patterns[1395] = 29'b0_000010101110_011_0_001010111000;
      patterns[1396] = 29'b0_000010101110_100_0_000001010111;
      patterns[1397] = 29'b0_000010101110_101_1_000000101011;
      patterns[1398] = 29'b0_000010101110_110_0_000010101110;
      patterns[1399] = 29'b0_000010101110_111_0_000010101110;
      patterns[1400] = 29'b0_000010101111_000_0_000010101111;
      patterns[1401] = 29'b0_000010101111_001_0_101111000010;
      patterns[1402] = 29'b0_000010101111_010_0_000101011110;
      patterns[1403] = 29'b0_000010101111_011_0_001010111100;
      patterns[1404] = 29'b0_000010101111_100_1_000001010111;
      patterns[1405] = 29'b0_000010101111_101_1_100000101011;
      patterns[1406] = 29'b0_000010101111_110_0_000010101111;
      patterns[1407] = 29'b0_000010101111_111_0_000010101111;
      patterns[1408] = 29'b0_000010110000_000_0_000010110000;
      patterns[1409] = 29'b0_000010110000_001_0_110000000010;
      patterns[1410] = 29'b0_000010110000_010_0_000101100000;
      patterns[1411] = 29'b0_000010110000_011_0_001011000000;
      patterns[1412] = 29'b0_000010110000_100_0_000001011000;
      patterns[1413] = 29'b0_000010110000_101_0_000000101100;
      patterns[1414] = 29'b0_000010110000_110_0_000010110000;
      patterns[1415] = 29'b0_000010110000_111_0_000010110000;
      patterns[1416] = 29'b0_000010110001_000_0_000010110001;
      patterns[1417] = 29'b0_000010110001_001_0_110001000010;
      patterns[1418] = 29'b0_000010110001_010_0_000101100010;
      patterns[1419] = 29'b0_000010110001_011_0_001011000100;
      patterns[1420] = 29'b0_000010110001_100_1_000001011000;
      patterns[1421] = 29'b0_000010110001_101_0_100000101100;
      patterns[1422] = 29'b0_000010110001_110_0_000010110001;
      patterns[1423] = 29'b0_000010110001_111_0_000010110001;
      patterns[1424] = 29'b0_000010110010_000_0_000010110010;
      patterns[1425] = 29'b0_000010110010_001_0_110010000010;
      patterns[1426] = 29'b0_000010110010_010_0_000101100100;
      patterns[1427] = 29'b0_000010110010_011_0_001011001000;
      patterns[1428] = 29'b0_000010110010_100_0_000001011001;
      patterns[1429] = 29'b0_000010110010_101_1_000000101100;
      patterns[1430] = 29'b0_000010110010_110_0_000010110010;
      patterns[1431] = 29'b0_000010110010_111_0_000010110010;
      patterns[1432] = 29'b0_000010110011_000_0_000010110011;
      patterns[1433] = 29'b0_000010110011_001_0_110011000010;
      patterns[1434] = 29'b0_000010110011_010_0_000101100110;
      patterns[1435] = 29'b0_000010110011_011_0_001011001100;
      patterns[1436] = 29'b0_000010110011_100_1_000001011001;
      patterns[1437] = 29'b0_000010110011_101_1_100000101100;
      patterns[1438] = 29'b0_000010110011_110_0_000010110011;
      patterns[1439] = 29'b0_000010110011_111_0_000010110011;
      patterns[1440] = 29'b0_000010110100_000_0_000010110100;
      patterns[1441] = 29'b0_000010110100_001_0_110100000010;
      patterns[1442] = 29'b0_000010110100_010_0_000101101000;
      patterns[1443] = 29'b0_000010110100_011_0_001011010000;
      patterns[1444] = 29'b0_000010110100_100_0_000001011010;
      patterns[1445] = 29'b0_000010110100_101_0_000000101101;
      patterns[1446] = 29'b0_000010110100_110_0_000010110100;
      patterns[1447] = 29'b0_000010110100_111_0_000010110100;
      patterns[1448] = 29'b0_000010110101_000_0_000010110101;
      patterns[1449] = 29'b0_000010110101_001_0_110101000010;
      patterns[1450] = 29'b0_000010110101_010_0_000101101010;
      patterns[1451] = 29'b0_000010110101_011_0_001011010100;
      patterns[1452] = 29'b0_000010110101_100_1_000001011010;
      patterns[1453] = 29'b0_000010110101_101_0_100000101101;
      patterns[1454] = 29'b0_000010110101_110_0_000010110101;
      patterns[1455] = 29'b0_000010110101_111_0_000010110101;
      patterns[1456] = 29'b0_000010110110_000_0_000010110110;
      patterns[1457] = 29'b0_000010110110_001_0_110110000010;
      patterns[1458] = 29'b0_000010110110_010_0_000101101100;
      patterns[1459] = 29'b0_000010110110_011_0_001011011000;
      patterns[1460] = 29'b0_000010110110_100_0_000001011011;
      patterns[1461] = 29'b0_000010110110_101_1_000000101101;
      patterns[1462] = 29'b0_000010110110_110_0_000010110110;
      patterns[1463] = 29'b0_000010110110_111_0_000010110110;
      patterns[1464] = 29'b0_000010110111_000_0_000010110111;
      patterns[1465] = 29'b0_000010110111_001_0_110111000010;
      patterns[1466] = 29'b0_000010110111_010_0_000101101110;
      patterns[1467] = 29'b0_000010110111_011_0_001011011100;
      patterns[1468] = 29'b0_000010110111_100_1_000001011011;
      patterns[1469] = 29'b0_000010110111_101_1_100000101101;
      patterns[1470] = 29'b0_000010110111_110_0_000010110111;
      patterns[1471] = 29'b0_000010110111_111_0_000010110111;
      patterns[1472] = 29'b0_000010111000_000_0_000010111000;
      patterns[1473] = 29'b0_000010111000_001_0_111000000010;
      patterns[1474] = 29'b0_000010111000_010_0_000101110000;
      patterns[1475] = 29'b0_000010111000_011_0_001011100000;
      patterns[1476] = 29'b0_000010111000_100_0_000001011100;
      patterns[1477] = 29'b0_000010111000_101_0_000000101110;
      patterns[1478] = 29'b0_000010111000_110_0_000010111000;
      patterns[1479] = 29'b0_000010111000_111_0_000010111000;
      patterns[1480] = 29'b0_000010111001_000_0_000010111001;
      patterns[1481] = 29'b0_000010111001_001_0_111001000010;
      patterns[1482] = 29'b0_000010111001_010_0_000101110010;
      patterns[1483] = 29'b0_000010111001_011_0_001011100100;
      patterns[1484] = 29'b0_000010111001_100_1_000001011100;
      patterns[1485] = 29'b0_000010111001_101_0_100000101110;
      patterns[1486] = 29'b0_000010111001_110_0_000010111001;
      patterns[1487] = 29'b0_000010111001_111_0_000010111001;
      patterns[1488] = 29'b0_000010111010_000_0_000010111010;
      patterns[1489] = 29'b0_000010111010_001_0_111010000010;
      patterns[1490] = 29'b0_000010111010_010_0_000101110100;
      patterns[1491] = 29'b0_000010111010_011_0_001011101000;
      patterns[1492] = 29'b0_000010111010_100_0_000001011101;
      patterns[1493] = 29'b0_000010111010_101_1_000000101110;
      patterns[1494] = 29'b0_000010111010_110_0_000010111010;
      patterns[1495] = 29'b0_000010111010_111_0_000010111010;
      patterns[1496] = 29'b0_000010111011_000_0_000010111011;
      patterns[1497] = 29'b0_000010111011_001_0_111011000010;
      patterns[1498] = 29'b0_000010111011_010_0_000101110110;
      patterns[1499] = 29'b0_000010111011_011_0_001011101100;
      patterns[1500] = 29'b0_000010111011_100_1_000001011101;
      patterns[1501] = 29'b0_000010111011_101_1_100000101110;
      patterns[1502] = 29'b0_000010111011_110_0_000010111011;
      patterns[1503] = 29'b0_000010111011_111_0_000010111011;
      patterns[1504] = 29'b0_000010111100_000_0_000010111100;
      patterns[1505] = 29'b0_000010111100_001_0_111100000010;
      patterns[1506] = 29'b0_000010111100_010_0_000101111000;
      patterns[1507] = 29'b0_000010111100_011_0_001011110000;
      patterns[1508] = 29'b0_000010111100_100_0_000001011110;
      patterns[1509] = 29'b0_000010111100_101_0_000000101111;
      patterns[1510] = 29'b0_000010111100_110_0_000010111100;
      patterns[1511] = 29'b0_000010111100_111_0_000010111100;
      patterns[1512] = 29'b0_000010111101_000_0_000010111101;
      patterns[1513] = 29'b0_000010111101_001_0_111101000010;
      patterns[1514] = 29'b0_000010111101_010_0_000101111010;
      patterns[1515] = 29'b0_000010111101_011_0_001011110100;
      patterns[1516] = 29'b0_000010111101_100_1_000001011110;
      patterns[1517] = 29'b0_000010111101_101_0_100000101111;
      patterns[1518] = 29'b0_000010111101_110_0_000010111101;
      patterns[1519] = 29'b0_000010111101_111_0_000010111101;
      patterns[1520] = 29'b0_000010111110_000_0_000010111110;
      patterns[1521] = 29'b0_000010111110_001_0_111110000010;
      patterns[1522] = 29'b0_000010111110_010_0_000101111100;
      patterns[1523] = 29'b0_000010111110_011_0_001011111000;
      patterns[1524] = 29'b0_000010111110_100_0_000001011111;
      patterns[1525] = 29'b0_000010111110_101_1_000000101111;
      patterns[1526] = 29'b0_000010111110_110_0_000010111110;
      patterns[1527] = 29'b0_000010111110_111_0_000010111110;
      patterns[1528] = 29'b0_000010111111_000_0_000010111111;
      patterns[1529] = 29'b0_000010111111_001_0_111111000010;
      patterns[1530] = 29'b0_000010111111_010_0_000101111110;
      patterns[1531] = 29'b0_000010111111_011_0_001011111100;
      patterns[1532] = 29'b0_000010111111_100_1_000001011111;
      patterns[1533] = 29'b0_000010111111_101_1_100000101111;
      patterns[1534] = 29'b0_000010111111_110_0_000010111111;
      patterns[1535] = 29'b0_000010111111_111_0_000010111111;
      patterns[1536] = 29'b0_000011000000_000_0_000011000000;
      patterns[1537] = 29'b0_000011000000_001_0_000000000011;
      patterns[1538] = 29'b0_000011000000_010_0_000110000000;
      patterns[1539] = 29'b0_000011000000_011_0_001100000000;
      patterns[1540] = 29'b0_000011000000_100_0_000001100000;
      patterns[1541] = 29'b0_000011000000_101_0_000000110000;
      patterns[1542] = 29'b0_000011000000_110_0_000011000000;
      patterns[1543] = 29'b0_000011000000_111_0_000011000000;
      patterns[1544] = 29'b0_000011000001_000_0_000011000001;
      patterns[1545] = 29'b0_000011000001_001_0_000001000011;
      patterns[1546] = 29'b0_000011000001_010_0_000110000010;
      patterns[1547] = 29'b0_000011000001_011_0_001100000100;
      patterns[1548] = 29'b0_000011000001_100_1_000001100000;
      patterns[1549] = 29'b0_000011000001_101_0_100000110000;
      patterns[1550] = 29'b0_000011000001_110_0_000011000001;
      patterns[1551] = 29'b0_000011000001_111_0_000011000001;
      patterns[1552] = 29'b0_000011000010_000_0_000011000010;
      patterns[1553] = 29'b0_000011000010_001_0_000010000011;
      patterns[1554] = 29'b0_000011000010_010_0_000110000100;
      patterns[1555] = 29'b0_000011000010_011_0_001100001000;
      patterns[1556] = 29'b0_000011000010_100_0_000001100001;
      patterns[1557] = 29'b0_000011000010_101_1_000000110000;
      patterns[1558] = 29'b0_000011000010_110_0_000011000010;
      patterns[1559] = 29'b0_000011000010_111_0_000011000010;
      patterns[1560] = 29'b0_000011000011_000_0_000011000011;
      patterns[1561] = 29'b0_000011000011_001_0_000011000011;
      patterns[1562] = 29'b0_000011000011_010_0_000110000110;
      patterns[1563] = 29'b0_000011000011_011_0_001100001100;
      patterns[1564] = 29'b0_000011000011_100_1_000001100001;
      patterns[1565] = 29'b0_000011000011_101_1_100000110000;
      patterns[1566] = 29'b0_000011000011_110_0_000011000011;
      patterns[1567] = 29'b0_000011000011_111_0_000011000011;
      patterns[1568] = 29'b0_000011000100_000_0_000011000100;
      patterns[1569] = 29'b0_000011000100_001_0_000100000011;
      patterns[1570] = 29'b0_000011000100_010_0_000110001000;
      patterns[1571] = 29'b0_000011000100_011_0_001100010000;
      patterns[1572] = 29'b0_000011000100_100_0_000001100010;
      patterns[1573] = 29'b0_000011000100_101_0_000000110001;
      patterns[1574] = 29'b0_000011000100_110_0_000011000100;
      patterns[1575] = 29'b0_000011000100_111_0_000011000100;
      patterns[1576] = 29'b0_000011000101_000_0_000011000101;
      patterns[1577] = 29'b0_000011000101_001_0_000101000011;
      patterns[1578] = 29'b0_000011000101_010_0_000110001010;
      patterns[1579] = 29'b0_000011000101_011_0_001100010100;
      patterns[1580] = 29'b0_000011000101_100_1_000001100010;
      patterns[1581] = 29'b0_000011000101_101_0_100000110001;
      patterns[1582] = 29'b0_000011000101_110_0_000011000101;
      patterns[1583] = 29'b0_000011000101_111_0_000011000101;
      patterns[1584] = 29'b0_000011000110_000_0_000011000110;
      patterns[1585] = 29'b0_000011000110_001_0_000110000011;
      patterns[1586] = 29'b0_000011000110_010_0_000110001100;
      patterns[1587] = 29'b0_000011000110_011_0_001100011000;
      patterns[1588] = 29'b0_000011000110_100_0_000001100011;
      patterns[1589] = 29'b0_000011000110_101_1_000000110001;
      patterns[1590] = 29'b0_000011000110_110_0_000011000110;
      patterns[1591] = 29'b0_000011000110_111_0_000011000110;
      patterns[1592] = 29'b0_000011000111_000_0_000011000111;
      patterns[1593] = 29'b0_000011000111_001_0_000111000011;
      patterns[1594] = 29'b0_000011000111_010_0_000110001110;
      patterns[1595] = 29'b0_000011000111_011_0_001100011100;
      patterns[1596] = 29'b0_000011000111_100_1_000001100011;
      patterns[1597] = 29'b0_000011000111_101_1_100000110001;
      patterns[1598] = 29'b0_000011000111_110_0_000011000111;
      patterns[1599] = 29'b0_000011000111_111_0_000011000111;
      patterns[1600] = 29'b0_000011001000_000_0_000011001000;
      patterns[1601] = 29'b0_000011001000_001_0_001000000011;
      patterns[1602] = 29'b0_000011001000_010_0_000110010000;
      patterns[1603] = 29'b0_000011001000_011_0_001100100000;
      patterns[1604] = 29'b0_000011001000_100_0_000001100100;
      patterns[1605] = 29'b0_000011001000_101_0_000000110010;
      patterns[1606] = 29'b0_000011001000_110_0_000011001000;
      patterns[1607] = 29'b0_000011001000_111_0_000011001000;
      patterns[1608] = 29'b0_000011001001_000_0_000011001001;
      patterns[1609] = 29'b0_000011001001_001_0_001001000011;
      patterns[1610] = 29'b0_000011001001_010_0_000110010010;
      patterns[1611] = 29'b0_000011001001_011_0_001100100100;
      patterns[1612] = 29'b0_000011001001_100_1_000001100100;
      patterns[1613] = 29'b0_000011001001_101_0_100000110010;
      patterns[1614] = 29'b0_000011001001_110_0_000011001001;
      patterns[1615] = 29'b0_000011001001_111_0_000011001001;
      patterns[1616] = 29'b0_000011001010_000_0_000011001010;
      patterns[1617] = 29'b0_000011001010_001_0_001010000011;
      patterns[1618] = 29'b0_000011001010_010_0_000110010100;
      patterns[1619] = 29'b0_000011001010_011_0_001100101000;
      patterns[1620] = 29'b0_000011001010_100_0_000001100101;
      patterns[1621] = 29'b0_000011001010_101_1_000000110010;
      patterns[1622] = 29'b0_000011001010_110_0_000011001010;
      patterns[1623] = 29'b0_000011001010_111_0_000011001010;
      patterns[1624] = 29'b0_000011001011_000_0_000011001011;
      patterns[1625] = 29'b0_000011001011_001_0_001011000011;
      patterns[1626] = 29'b0_000011001011_010_0_000110010110;
      patterns[1627] = 29'b0_000011001011_011_0_001100101100;
      patterns[1628] = 29'b0_000011001011_100_1_000001100101;
      patterns[1629] = 29'b0_000011001011_101_1_100000110010;
      patterns[1630] = 29'b0_000011001011_110_0_000011001011;
      patterns[1631] = 29'b0_000011001011_111_0_000011001011;
      patterns[1632] = 29'b0_000011001100_000_0_000011001100;
      patterns[1633] = 29'b0_000011001100_001_0_001100000011;
      patterns[1634] = 29'b0_000011001100_010_0_000110011000;
      patterns[1635] = 29'b0_000011001100_011_0_001100110000;
      patterns[1636] = 29'b0_000011001100_100_0_000001100110;
      patterns[1637] = 29'b0_000011001100_101_0_000000110011;
      patterns[1638] = 29'b0_000011001100_110_0_000011001100;
      patterns[1639] = 29'b0_000011001100_111_0_000011001100;
      patterns[1640] = 29'b0_000011001101_000_0_000011001101;
      patterns[1641] = 29'b0_000011001101_001_0_001101000011;
      patterns[1642] = 29'b0_000011001101_010_0_000110011010;
      patterns[1643] = 29'b0_000011001101_011_0_001100110100;
      patterns[1644] = 29'b0_000011001101_100_1_000001100110;
      patterns[1645] = 29'b0_000011001101_101_0_100000110011;
      patterns[1646] = 29'b0_000011001101_110_0_000011001101;
      patterns[1647] = 29'b0_000011001101_111_0_000011001101;
      patterns[1648] = 29'b0_000011001110_000_0_000011001110;
      patterns[1649] = 29'b0_000011001110_001_0_001110000011;
      patterns[1650] = 29'b0_000011001110_010_0_000110011100;
      patterns[1651] = 29'b0_000011001110_011_0_001100111000;
      patterns[1652] = 29'b0_000011001110_100_0_000001100111;
      patterns[1653] = 29'b0_000011001110_101_1_000000110011;
      patterns[1654] = 29'b0_000011001110_110_0_000011001110;
      patterns[1655] = 29'b0_000011001110_111_0_000011001110;
      patterns[1656] = 29'b0_000011001111_000_0_000011001111;
      patterns[1657] = 29'b0_000011001111_001_0_001111000011;
      patterns[1658] = 29'b0_000011001111_010_0_000110011110;
      patterns[1659] = 29'b0_000011001111_011_0_001100111100;
      patterns[1660] = 29'b0_000011001111_100_1_000001100111;
      patterns[1661] = 29'b0_000011001111_101_1_100000110011;
      patterns[1662] = 29'b0_000011001111_110_0_000011001111;
      patterns[1663] = 29'b0_000011001111_111_0_000011001111;
      patterns[1664] = 29'b0_000011010000_000_0_000011010000;
      patterns[1665] = 29'b0_000011010000_001_0_010000000011;
      patterns[1666] = 29'b0_000011010000_010_0_000110100000;
      patterns[1667] = 29'b0_000011010000_011_0_001101000000;
      patterns[1668] = 29'b0_000011010000_100_0_000001101000;
      patterns[1669] = 29'b0_000011010000_101_0_000000110100;
      patterns[1670] = 29'b0_000011010000_110_0_000011010000;
      patterns[1671] = 29'b0_000011010000_111_0_000011010000;
      patterns[1672] = 29'b0_000011010001_000_0_000011010001;
      patterns[1673] = 29'b0_000011010001_001_0_010001000011;
      patterns[1674] = 29'b0_000011010001_010_0_000110100010;
      patterns[1675] = 29'b0_000011010001_011_0_001101000100;
      patterns[1676] = 29'b0_000011010001_100_1_000001101000;
      patterns[1677] = 29'b0_000011010001_101_0_100000110100;
      patterns[1678] = 29'b0_000011010001_110_0_000011010001;
      patterns[1679] = 29'b0_000011010001_111_0_000011010001;
      patterns[1680] = 29'b0_000011010010_000_0_000011010010;
      patterns[1681] = 29'b0_000011010010_001_0_010010000011;
      patterns[1682] = 29'b0_000011010010_010_0_000110100100;
      patterns[1683] = 29'b0_000011010010_011_0_001101001000;
      patterns[1684] = 29'b0_000011010010_100_0_000001101001;
      patterns[1685] = 29'b0_000011010010_101_1_000000110100;
      patterns[1686] = 29'b0_000011010010_110_0_000011010010;
      patterns[1687] = 29'b0_000011010010_111_0_000011010010;
      patterns[1688] = 29'b0_000011010011_000_0_000011010011;
      patterns[1689] = 29'b0_000011010011_001_0_010011000011;
      patterns[1690] = 29'b0_000011010011_010_0_000110100110;
      patterns[1691] = 29'b0_000011010011_011_0_001101001100;
      patterns[1692] = 29'b0_000011010011_100_1_000001101001;
      patterns[1693] = 29'b0_000011010011_101_1_100000110100;
      patterns[1694] = 29'b0_000011010011_110_0_000011010011;
      patterns[1695] = 29'b0_000011010011_111_0_000011010011;
      patterns[1696] = 29'b0_000011010100_000_0_000011010100;
      patterns[1697] = 29'b0_000011010100_001_0_010100000011;
      patterns[1698] = 29'b0_000011010100_010_0_000110101000;
      patterns[1699] = 29'b0_000011010100_011_0_001101010000;
      patterns[1700] = 29'b0_000011010100_100_0_000001101010;
      patterns[1701] = 29'b0_000011010100_101_0_000000110101;
      patterns[1702] = 29'b0_000011010100_110_0_000011010100;
      patterns[1703] = 29'b0_000011010100_111_0_000011010100;
      patterns[1704] = 29'b0_000011010101_000_0_000011010101;
      patterns[1705] = 29'b0_000011010101_001_0_010101000011;
      patterns[1706] = 29'b0_000011010101_010_0_000110101010;
      patterns[1707] = 29'b0_000011010101_011_0_001101010100;
      patterns[1708] = 29'b0_000011010101_100_1_000001101010;
      patterns[1709] = 29'b0_000011010101_101_0_100000110101;
      patterns[1710] = 29'b0_000011010101_110_0_000011010101;
      patterns[1711] = 29'b0_000011010101_111_0_000011010101;
      patterns[1712] = 29'b0_000011010110_000_0_000011010110;
      patterns[1713] = 29'b0_000011010110_001_0_010110000011;
      patterns[1714] = 29'b0_000011010110_010_0_000110101100;
      patterns[1715] = 29'b0_000011010110_011_0_001101011000;
      patterns[1716] = 29'b0_000011010110_100_0_000001101011;
      patterns[1717] = 29'b0_000011010110_101_1_000000110101;
      patterns[1718] = 29'b0_000011010110_110_0_000011010110;
      patterns[1719] = 29'b0_000011010110_111_0_000011010110;
      patterns[1720] = 29'b0_000011010111_000_0_000011010111;
      patterns[1721] = 29'b0_000011010111_001_0_010111000011;
      patterns[1722] = 29'b0_000011010111_010_0_000110101110;
      patterns[1723] = 29'b0_000011010111_011_0_001101011100;
      patterns[1724] = 29'b0_000011010111_100_1_000001101011;
      patterns[1725] = 29'b0_000011010111_101_1_100000110101;
      patterns[1726] = 29'b0_000011010111_110_0_000011010111;
      patterns[1727] = 29'b0_000011010111_111_0_000011010111;
      patterns[1728] = 29'b0_000011011000_000_0_000011011000;
      patterns[1729] = 29'b0_000011011000_001_0_011000000011;
      patterns[1730] = 29'b0_000011011000_010_0_000110110000;
      patterns[1731] = 29'b0_000011011000_011_0_001101100000;
      patterns[1732] = 29'b0_000011011000_100_0_000001101100;
      patterns[1733] = 29'b0_000011011000_101_0_000000110110;
      patterns[1734] = 29'b0_000011011000_110_0_000011011000;
      patterns[1735] = 29'b0_000011011000_111_0_000011011000;
      patterns[1736] = 29'b0_000011011001_000_0_000011011001;
      patterns[1737] = 29'b0_000011011001_001_0_011001000011;
      patterns[1738] = 29'b0_000011011001_010_0_000110110010;
      patterns[1739] = 29'b0_000011011001_011_0_001101100100;
      patterns[1740] = 29'b0_000011011001_100_1_000001101100;
      patterns[1741] = 29'b0_000011011001_101_0_100000110110;
      patterns[1742] = 29'b0_000011011001_110_0_000011011001;
      patterns[1743] = 29'b0_000011011001_111_0_000011011001;
      patterns[1744] = 29'b0_000011011010_000_0_000011011010;
      patterns[1745] = 29'b0_000011011010_001_0_011010000011;
      patterns[1746] = 29'b0_000011011010_010_0_000110110100;
      patterns[1747] = 29'b0_000011011010_011_0_001101101000;
      patterns[1748] = 29'b0_000011011010_100_0_000001101101;
      patterns[1749] = 29'b0_000011011010_101_1_000000110110;
      patterns[1750] = 29'b0_000011011010_110_0_000011011010;
      patterns[1751] = 29'b0_000011011010_111_0_000011011010;
      patterns[1752] = 29'b0_000011011011_000_0_000011011011;
      patterns[1753] = 29'b0_000011011011_001_0_011011000011;
      patterns[1754] = 29'b0_000011011011_010_0_000110110110;
      patterns[1755] = 29'b0_000011011011_011_0_001101101100;
      patterns[1756] = 29'b0_000011011011_100_1_000001101101;
      patterns[1757] = 29'b0_000011011011_101_1_100000110110;
      patterns[1758] = 29'b0_000011011011_110_0_000011011011;
      patterns[1759] = 29'b0_000011011011_111_0_000011011011;
      patterns[1760] = 29'b0_000011011100_000_0_000011011100;
      patterns[1761] = 29'b0_000011011100_001_0_011100000011;
      patterns[1762] = 29'b0_000011011100_010_0_000110111000;
      patterns[1763] = 29'b0_000011011100_011_0_001101110000;
      patterns[1764] = 29'b0_000011011100_100_0_000001101110;
      patterns[1765] = 29'b0_000011011100_101_0_000000110111;
      patterns[1766] = 29'b0_000011011100_110_0_000011011100;
      patterns[1767] = 29'b0_000011011100_111_0_000011011100;
      patterns[1768] = 29'b0_000011011101_000_0_000011011101;
      patterns[1769] = 29'b0_000011011101_001_0_011101000011;
      patterns[1770] = 29'b0_000011011101_010_0_000110111010;
      patterns[1771] = 29'b0_000011011101_011_0_001101110100;
      patterns[1772] = 29'b0_000011011101_100_1_000001101110;
      patterns[1773] = 29'b0_000011011101_101_0_100000110111;
      patterns[1774] = 29'b0_000011011101_110_0_000011011101;
      patterns[1775] = 29'b0_000011011101_111_0_000011011101;
      patterns[1776] = 29'b0_000011011110_000_0_000011011110;
      patterns[1777] = 29'b0_000011011110_001_0_011110000011;
      patterns[1778] = 29'b0_000011011110_010_0_000110111100;
      patterns[1779] = 29'b0_000011011110_011_0_001101111000;
      patterns[1780] = 29'b0_000011011110_100_0_000001101111;
      patterns[1781] = 29'b0_000011011110_101_1_000000110111;
      patterns[1782] = 29'b0_000011011110_110_0_000011011110;
      patterns[1783] = 29'b0_000011011110_111_0_000011011110;
      patterns[1784] = 29'b0_000011011111_000_0_000011011111;
      patterns[1785] = 29'b0_000011011111_001_0_011111000011;
      patterns[1786] = 29'b0_000011011111_010_0_000110111110;
      patterns[1787] = 29'b0_000011011111_011_0_001101111100;
      patterns[1788] = 29'b0_000011011111_100_1_000001101111;
      patterns[1789] = 29'b0_000011011111_101_1_100000110111;
      patterns[1790] = 29'b0_000011011111_110_0_000011011111;
      patterns[1791] = 29'b0_000011011111_111_0_000011011111;
      patterns[1792] = 29'b0_000011100000_000_0_000011100000;
      patterns[1793] = 29'b0_000011100000_001_0_100000000011;
      patterns[1794] = 29'b0_000011100000_010_0_000111000000;
      patterns[1795] = 29'b0_000011100000_011_0_001110000000;
      patterns[1796] = 29'b0_000011100000_100_0_000001110000;
      patterns[1797] = 29'b0_000011100000_101_0_000000111000;
      patterns[1798] = 29'b0_000011100000_110_0_000011100000;
      patterns[1799] = 29'b0_000011100000_111_0_000011100000;
      patterns[1800] = 29'b0_000011100001_000_0_000011100001;
      patterns[1801] = 29'b0_000011100001_001_0_100001000011;
      patterns[1802] = 29'b0_000011100001_010_0_000111000010;
      patterns[1803] = 29'b0_000011100001_011_0_001110000100;
      patterns[1804] = 29'b0_000011100001_100_1_000001110000;
      patterns[1805] = 29'b0_000011100001_101_0_100000111000;
      patterns[1806] = 29'b0_000011100001_110_0_000011100001;
      patterns[1807] = 29'b0_000011100001_111_0_000011100001;
      patterns[1808] = 29'b0_000011100010_000_0_000011100010;
      patterns[1809] = 29'b0_000011100010_001_0_100010000011;
      patterns[1810] = 29'b0_000011100010_010_0_000111000100;
      patterns[1811] = 29'b0_000011100010_011_0_001110001000;
      patterns[1812] = 29'b0_000011100010_100_0_000001110001;
      patterns[1813] = 29'b0_000011100010_101_1_000000111000;
      patterns[1814] = 29'b0_000011100010_110_0_000011100010;
      patterns[1815] = 29'b0_000011100010_111_0_000011100010;
      patterns[1816] = 29'b0_000011100011_000_0_000011100011;
      patterns[1817] = 29'b0_000011100011_001_0_100011000011;
      patterns[1818] = 29'b0_000011100011_010_0_000111000110;
      patterns[1819] = 29'b0_000011100011_011_0_001110001100;
      patterns[1820] = 29'b0_000011100011_100_1_000001110001;
      patterns[1821] = 29'b0_000011100011_101_1_100000111000;
      patterns[1822] = 29'b0_000011100011_110_0_000011100011;
      patterns[1823] = 29'b0_000011100011_111_0_000011100011;
      patterns[1824] = 29'b0_000011100100_000_0_000011100100;
      patterns[1825] = 29'b0_000011100100_001_0_100100000011;
      patterns[1826] = 29'b0_000011100100_010_0_000111001000;
      patterns[1827] = 29'b0_000011100100_011_0_001110010000;
      patterns[1828] = 29'b0_000011100100_100_0_000001110010;
      patterns[1829] = 29'b0_000011100100_101_0_000000111001;
      patterns[1830] = 29'b0_000011100100_110_0_000011100100;
      patterns[1831] = 29'b0_000011100100_111_0_000011100100;
      patterns[1832] = 29'b0_000011100101_000_0_000011100101;
      patterns[1833] = 29'b0_000011100101_001_0_100101000011;
      patterns[1834] = 29'b0_000011100101_010_0_000111001010;
      patterns[1835] = 29'b0_000011100101_011_0_001110010100;
      patterns[1836] = 29'b0_000011100101_100_1_000001110010;
      patterns[1837] = 29'b0_000011100101_101_0_100000111001;
      patterns[1838] = 29'b0_000011100101_110_0_000011100101;
      patterns[1839] = 29'b0_000011100101_111_0_000011100101;
      patterns[1840] = 29'b0_000011100110_000_0_000011100110;
      patterns[1841] = 29'b0_000011100110_001_0_100110000011;
      patterns[1842] = 29'b0_000011100110_010_0_000111001100;
      patterns[1843] = 29'b0_000011100110_011_0_001110011000;
      patterns[1844] = 29'b0_000011100110_100_0_000001110011;
      patterns[1845] = 29'b0_000011100110_101_1_000000111001;
      patterns[1846] = 29'b0_000011100110_110_0_000011100110;
      patterns[1847] = 29'b0_000011100110_111_0_000011100110;
      patterns[1848] = 29'b0_000011100111_000_0_000011100111;
      patterns[1849] = 29'b0_000011100111_001_0_100111000011;
      patterns[1850] = 29'b0_000011100111_010_0_000111001110;
      patterns[1851] = 29'b0_000011100111_011_0_001110011100;
      patterns[1852] = 29'b0_000011100111_100_1_000001110011;
      patterns[1853] = 29'b0_000011100111_101_1_100000111001;
      patterns[1854] = 29'b0_000011100111_110_0_000011100111;
      patterns[1855] = 29'b0_000011100111_111_0_000011100111;
      patterns[1856] = 29'b0_000011101000_000_0_000011101000;
      patterns[1857] = 29'b0_000011101000_001_0_101000000011;
      patterns[1858] = 29'b0_000011101000_010_0_000111010000;
      patterns[1859] = 29'b0_000011101000_011_0_001110100000;
      patterns[1860] = 29'b0_000011101000_100_0_000001110100;
      patterns[1861] = 29'b0_000011101000_101_0_000000111010;
      patterns[1862] = 29'b0_000011101000_110_0_000011101000;
      patterns[1863] = 29'b0_000011101000_111_0_000011101000;
      patterns[1864] = 29'b0_000011101001_000_0_000011101001;
      patterns[1865] = 29'b0_000011101001_001_0_101001000011;
      patterns[1866] = 29'b0_000011101001_010_0_000111010010;
      patterns[1867] = 29'b0_000011101001_011_0_001110100100;
      patterns[1868] = 29'b0_000011101001_100_1_000001110100;
      patterns[1869] = 29'b0_000011101001_101_0_100000111010;
      patterns[1870] = 29'b0_000011101001_110_0_000011101001;
      patterns[1871] = 29'b0_000011101001_111_0_000011101001;
      patterns[1872] = 29'b0_000011101010_000_0_000011101010;
      patterns[1873] = 29'b0_000011101010_001_0_101010000011;
      patterns[1874] = 29'b0_000011101010_010_0_000111010100;
      patterns[1875] = 29'b0_000011101010_011_0_001110101000;
      patterns[1876] = 29'b0_000011101010_100_0_000001110101;
      patterns[1877] = 29'b0_000011101010_101_1_000000111010;
      patterns[1878] = 29'b0_000011101010_110_0_000011101010;
      patterns[1879] = 29'b0_000011101010_111_0_000011101010;
      patterns[1880] = 29'b0_000011101011_000_0_000011101011;
      patterns[1881] = 29'b0_000011101011_001_0_101011000011;
      patterns[1882] = 29'b0_000011101011_010_0_000111010110;
      patterns[1883] = 29'b0_000011101011_011_0_001110101100;
      patterns[1884] = 29'b0_000011101011_100_1_000001110101;
      patterns[1885] = 29'b0_000011101011_101_1_100000111010;
      patterns[1886] = 29'b0_000011101011_110_0_000011101011;
      patterns[1887] = 29'b0_000011101011_111_0_000011101011;
      patterns[1888] = 29'b0_000011101100_000_0_000011101100;
      patterns[1889] = 29'b0_000011101100_001_0_101100000011;
      patterns[1890] = 29'b0_000011101100_010_0_000111011000;
      patterns[1891] = 29'b0_000011101100_011_0_001110110000;
      patterns[1892] = 29'b0_000011101100_100_0_000001110110;
      patterns[1893] = 29'b0_000011101100_101_0_000000111011;
      patterns[1894] = 29'b0_000011101100_110_0_000011101100;
      patterns[1895] = 29'b0_000011101100_111_0_000011101100;
      patterns[1896] = 29'b0_000011101101_000_0_000011101101;
      patterns[1897] = 29'b0_000011101101_001_0_101101000011;
      patterns[1898] = 29'b0_000011101101_010_0_000111011010;
      patterns[1899] = 29'b0_000011101101_011_0_001110110100;
      patterns[1900] = 29'b0_000011101101_100_1_000001110110;
      patterns[1901] = 29'b0_000011101101_101_0_100000111011;
      patterns[1902] = 29'b0_000011101101_110_0_000011101101;
      patterns[1903] = 29'b0_000011101101_111_0_000011101101;
      patterns[1904] = 29'b0_000011101110_000_0_000011101110;
      patterns[1905] = 29'b0_000011101110_001_0_101110000011;
      patterns[1906] = 29'b0_000011101110_010_0_000111011100;
      patterns[1907] = 29'b0_000011101110_011_0_001110111000;
      patterns[1908] = 29'b0_000011101110_100_0_000001110111;
      patterns[1909] = 29'b0_000011101110_101_1_000000111011;
      patterns[1910] = 29'b0_000011101110_110_0_000011101110;
      patterns[1911] = 29'b0_000011101110_111_0_000011101110;
      patterns[1912] = 29'b0_000011101111_000_0_000011101111;
      patterns[1913] = 29'b0_000011101111_001_0_101111000011;
      patterns[1914] = 29'b0_000011101111_010_0_000111011110;
      patterns[1915] = 29'b0_000011101111_011_0_001110111100;
      patterns[1916] = 29'b0_000011101111_100_1_000001110111;
      patterns[1917] = 29'b0_000011101111_101_1_100000111011;
      patterns[1918] = 29'b0_000011101111_110_0_000011101111;
      patterns[1919] = 29'b0_000011101111_111_0_000011101111;
      patterns[1920] = 29'b0_000011110000_000_0_000011110000;
      patterns[1921] = 29'b0_000011110000_001_0_110000000011;
      patterns[1922] = 29'b0_000011110000_010_0_000111100000;
      patterns[1923] = 29'b0_000011110000_011_0_001111000000;
      patterns[1924] = 29'b0_000011110000_100_0_000001111000;
      patterns[1925] = 29'b0_000011110000_101_0_000000111100;
      patterns[1926] = 29'b0_000011110000_110_0_000011110000;
      patterns[1927] = 29'b0_000011110000_111_0_000011110000;
      patterns[1928] = 29'b0_000011110001_000_0_000011110001;
      patterns[1929] = 29'b0_000011110001_001_0_110001000011;
      patterns[1930] = 29'b0_000011110001_010_0_000111100010;
      patterns[1931] = 29'b0_000011110001_011_0_001111000100;
      patterns[1932] = 29'b0_000011110001_100_1_000001111000;
      patterns[1933] = 29'b0_000011110001_101_0_100000111100;
      patterns[1934] = 29'b0_000011110001_110_0_000011110001;
      patterns[1935] = 29'b0_000011110001_111_0_000011110001;
      patterns[1936] = 29'b0_000011110010_000_0_000011110010;
      patterns[1937] = 29'b0_000011110010_001_0_110010000011;
      patterns[1938] = 29'b0_000011110010_010_0_000111100100;
      patterns[1939] = 29'b0_000011110010_011_0_001111001000;
      patterns[1940] = 29'b0_000011110010_100_0_000001111001;
      patterns[1941] = 29'b0_000011110010_101_1_000000111100;
      patterns[1942] = 29'b0_000011110010_110_0_000011110010;
      patterns[1943] = 29'b0_000011110010_111_0_000011110010;
      patterns[1944] = 29'b0_000011110011_000_0_000011110011;
      patterns[1945] = 29'b0_000011110011_001_0_110011000011;
      patterns[1946] = 29'b0_000011110011_010_0_000111100110;
      patterns[1947] = 29'b0_000011110011_011_0_001111001100;
      patterns[1948] = 29'b0_000011110011_100_1_000001111001;
      patterns[1949] = 29'b0_000011110011_101_1_100000111100;
      patterns[1950] = 29'b0_000011110011_110_0_000011110011;
      patterns[1951] = 29'b0_000011110011_111_0_000011110011;
      patterns[1952] = 29'b0_000011110100_000_0_000011110100;
      patterns[1953] = 29'b0_000011110100_001_0_110100000011;
      patterns[1954] = 29'b0_000011110100_010_0_000111101000;
      patterns[1955] = 29'b0_000011110100_011_0_001111010000;
      patterns[1956] = 29'b0_000011110100_100_0_000001111010;
      patterns[1957] = 29'b0_000011110100_101_0_000000111101;
      patterns[1958] = 29'b0_000011110100_110_0_000011110100;
      patterns[1959] = 29'b0_000011110100_111_0_000011110100;
      patterns[1960] = 29'b0_000011110101_000_0_000011110101;
      patterns[1961] = 29'b0_000011110101_001_0_110101000011;
      patterns[1962] = 29'b0_000011110101_010_0_000111101010;
      patterns[1963] = 29'b0_000011110101_011_0_001111010100;
      patterns[1964] = 29'b0_000011110101_100_1_000001111010;
      patterns[1965] = 29'b0_000011110101_101_0_100000111101;
      patterns[1966] = 29'b0_000011110101_110_0_000011110101;
      patterns[1967] = 29'b0_000011110101_111_0_000011110101;
      patterns[1968] = 29'b0_000011110110_000_0_000011110110;
      patterns[1969] = 29'b0_000011110110_001_0_110110000011;
      patterns[1970] = 29'b0_000011110110_010_0_000111101100;
      patterns[1971] = 29'b0_000011110110_011_0_001111011000;
      patterns[1972] = 29'b0_000011110110_100_0_000001111011;
      patterns[1973] = 29'b0_000011110110_101_1_000000111101;
      patterns[1974] = 29'b0_000011110110_110_0_000011110110;
      patterns[1975] = 29'b0_000011110110_111_0_000011110110;
      patterns[1976] = 29'b0_000011110111_000_0_000011110111;
      patterns[1977] = 29'b0_000011110111_001_0_110111000011;
      patterns[1978] = 29'b0_000011110111_010_0_000111101110;
      patterns[1979] = 29'b0_000011110111_011_0_001111011100;
      patterns[1980] = 29'b0_000011110111_100_1_000001111011;
      patterns[1981] = 29'b0_000011110111_101_1_100000111101;
      patterns[1982] = 29'b0_000011110111_110_0_000011110111;
      patterns[1983] = 29'b0_000011110111_111_0_000011110111;
      patterns[1984] = 29'b0_000011111000_000_0_000011111000;
      patterns[1985] = 29'b0_000011111000_001_0_111000000011;
      patterns[1986] = 29'b0_000011111000_010_0_000111110000;
      patterns[1987] = 29'b0_000011111000_011_0_001111100000;
      patterns[1988] = 29'b0_000011111000_100_0_000001111100;
      patterns[1989] = 29'b0_000011111000_101_0_000000111110;
      patterns[1990] = 29'b0_000011111000_110_0_000011111000;
      patterns[1991] = 29'b0_000011111000_111_0_000011111000;
      patterns[1992] = 29'b0_000011111001_000_0_000011111001;
      patterns[1993] = 29'b0_000011111001_001_0_111001000011;
      patterns[1994] = 29'b0_000011111001_010_0_000111110010;
      patterns[1995] = 29'b0_000011111001_011_0_001111100100;
      patterns[1996] = 29'b0_000011111001_100_1_000001111100;
      patterns[1997] = 29'b0_000011111001_101_0_100000111110;
      patterns[1998] = 29'b0_000011111001_110_0_000011111001;
      patterns[1999] = 29'b0_000011111001_111_0_000011111001;
      patterns[2000] = 29'b0_000011111010_000_0_000011111010;
      patterns[2001] = 29'b0_000011111010_001_0_111010000011;
      patterns[2002] = 29'b0_000011111010_010_0_000111110100;
      patterns[2003] = 29'b0_000011111010_011_0_001111101000;
      patterns[2004] = 29'b0_000011111010_100_0_000001111101;
      patterns[2005] = 29'b0_000011111010_101_1_000000111110;
      patterns[2006] = 29'b0_000011111010_110_0_000011111010;
      patterns[2007] = 29'b0_000011111010_111_0_000011111010;
      patterns[2008] = 29'b0_000011111011_000_0_000011111011;
      patterns[2009] = 29'b0_000011111011_001_0_111011000011;
      patterns[2010] = 29'b0_000011111011_010_0_000111110110;
      patterns[2011] = 29'b0_000011111011_011_0_001111101100;
      patterns[2012] = 29'b0_000011111011_100_1_000001111101;
      patterns[2013] = 29'b0_000011111011_101_1_100000111110;
      patterns[2014] = 29'b0_000011111011_110_0_000011111011;
      patterns[2015] = 29'b0_000011111011_111_0_000011111011;
      patterns[2016] = 29'b0_000011111100_000_0_000011111100;
      patterns[2017] = 29'b0_000011111100_001_0_111100000011;
      patterns[2018] = 29'b0_000011111100_010_0_000111111000;
      patterns[2019] = 29'b0_000011111100_011_0_001111110000;
      patterns[2020] = 29'b0_000011111100_100_0_000001111110;
      patterns[2021] = 29'b0_000011111100_101_0_000000111111;
      patterns[2022] = 29'b0_000011111100_110_0_000011111100;
      patterns[2023] = 29'b0_000011111100_111_0_000011111100;
      patterns[2024] = 29'b0_000011111101_000_0_000011111101;
      patterns[2025] = 29'b0_000011111101_001_0_111101000011;
      patterns[2026] = 29'b0_000011111101_010_0_000111111010;
      patterns[2027] = 29'b0_000011111101_011_0_001111110100;
      patterns[2028] = 29'b0_000011111101_100_1_000001111110;
      patterns[2029] = 29'b0_000011111101_101_0_100000111111;
      patterns[2030] = 29'b0_000011111101_110_0_000011111101;
      patterns[2031] = 29'b0_000011111101_111_0_000011111101;
      patterns[2032] = 29'b0_000011111110_000_0_000011111110;
      patterns[2033] = 29'b0_000011111110_001_0_111110000011;
      patterns[2034] = 29'b0_000011111110_010_0_000111111100;
      patterns[2035] = 29'b0_000011111110_011_0_001111111000;
      patterns[2036] = 29'b0_000011111110_100_0_000001111111;
      patterns[2037] = 29'b0_000011111110_101_1_000000111111;
      patterns[2038] = 29'b0_000011111110_110_0_000011111110;
      patterns[2039] = 29'b0_000011111110_111_0_000011111110;
      patterns[2040] = 29'b0_000011111111_000_0_000011111111;
      patterns[2041] = 29'b0_000011111111_001_0_111111000011;
      patterns[2042] = 29'b0_000011111111_010_0_000111111110;
      patterns[2043] = 29'b0_000011111111_011_0_001111111100;
      patterns[2044] = 29'b0_000011111111_100_1_000001111111;
      patterns[2045] = 29'b0_000011111111_101_1_100000111111;
      patterns[2046] = 29'b0_000011111111_110_0_000011111111;
      patterns[2047] = 29'b0_000011111111_111_0_000011111111;
      patterns[2048] = 29'b0_000100000000_000_0_000100000000;
      patterns[2049] = 29'b0_000100000000_001_0_000000000100;
      patterns[2050] = 29'b0_000100000000_010_0_001000000000;
      patterns[2051] = 29'b0_000100000000_011_0_010000000000;
      patterns[2052] = 29'b0_000100000000_100_0_000010000000;
      patterns[2053] = 29'b0_000100000000_101_0_000001000000;
      patterns[2054] = 29'b0_000100000000_110_0_000100000000;
      patterns[2055] = 29'b0_000100000000_111_0_000100000000;
      patterns[2056] = 29'b0_000100000001_000_0_000100000001;
      patterns[2057] = 29'b0_000100000001_001_0_000001000100;
      patterns[2058] = 29'b0_000100000001_010_0_001000000010;
      patterns[2059] = 29'b0_000100000001_011_0_010000000100;
      patterns[2060] = 29'b0_000100000001_100_1_000010000000;
      patterns[2061] = 29'b0_000100000001_101_0_100001000000;
      patterns[2062] = 29'b0_000100000001_110_0_000100000001;
      patterns[2063] = 29'b0_000100000001_111_0_000100000001;
      patterns[2064] = 29'b0_000100000010_000_0_000100000010;
      patterns[2065] = 29'b0_000100000010_001_0_000010000100;
      patterns[2066] = 29'b0_000100000010_010_0_001000000100;
      patterns[2067] = 29'b0_000100000010_011_0_010000001000;
      patterns[2068] = 29'b0_000100000010_100_0_000010000001;
      patterns[2069] = 29'b0_000100000010_101_1_000001000000;
      patterns[2070] = 29'b0_000100000010_110_0_000100000010;
      patterns[2071] = 29'b0_000100000010_111_0_000100000010;
      patterns[2072] = 29'b0_000100000011_000_0_000100000011;
      patterns[2073] = 29'b0_000100000011_001_0_000011000100;
      patterns[2074] = 29'b0_000100000011_010_0_001000000110;
      patterns[2075] = 29'b0_000100000011_011_0_010000001100;
      patterns[2076] = 29'b0_000100000011_100_1_000010000001;
      patterns[2077] = 29'b0_000100000011_101_1_100001000000;
      patterns[2078] = 29'b0_000100000011_110_0_000100000011;
      patterns[2079] = 29'b0_000100000011_111_0_000100000011;
      patterns[2080] = 29'b0_000100000100_000_0_000100000100;
      patterns[2081] = 29'b0_000100000100_001_0_000100000100;
      patterns[2082] = 29'b0_000100000100_010_0_001000001000;
      patterns[2083] = 29'b0_000100000100_011_0_010000010000;
      patterns[2084] = 29'b0_000100000100_100_0_000010000010;
      patterns[2085] = 29'b0_000100000100_101_0_000001000001;
      patterns[2086] = 29'b0_000100000100_110_0_000100000100;
      patterns[2087] = 29'b0_000100000100_111_0_000100000100;
      patterns[2088] = 29'b0_000100000101_000_0_000100000101;
      patterns[2089] = 29'b0_000100000101_001_0_000101000100;
      patterns[2090] = 29'b0_000100000101_010_0_001000001010;
      patterns[2091] = 29'b0_000100000101_011_0_010000010100;
      patterns[2092] = 29'b0_000100000101_100_1_000010000010;
      patterns[2093] = 29'b0_000100000101_101_0_100001000001;
      patterns[2094] = 29'b0_000100000101_110_0_000100000101;
      patterns[2095] = 29'b0_000100000101_111_0_000100000101;
      patterns[2096] = 29'b0_000100000110_000_0_000100000110;
      patterns[2097] = 29'b0_000100000110_001_0_000110000100;
      patterns[2098] = 29'b0_000100000110_010_0_001000001100;
      patterns[2099] = 29'b0_000100000110_011_0_010000011000;
      patterns[2100] = 29'b0_000100000110_100_0_000010000011;
      patterns[2101] = 29'b0_000100000110_101_1_000001000001;
      patterns[2102] = 29'b0_000100000110_110_0_000100000110;
      patterns[2103] = 29'b0_000100000110_111_0_000100000110;
      patterns[2104] = 29'b0_000100000111_000_0_000100000111;
      patterns[2105] = 29'b0_000100000111_001_0_000111000100;
      patterns[2106] = 29'b0_000100000111_010_0_001000001110;
      patterns[2107] = 29'b0_000100000111_011_0_010000011100;
      patterns[2108] = 29'b0_000100000111_100_1_000010000011;
      patterns[2109] = 29'b0_000100000111_101_1_100001000001;
      patterns[2110] = 29'b0_000100000111_110_0_000100000111;
      patterns[2111] = 29'b0_000100000111_111_0_000100000111;
      patterns[2112] = 29'b0_000100001000_000_0_000100001000;
      patterns[2113] = 29'b0_000100001000_001_0_001000000100;
      patterns[2114] = 29'b0_000100001000_010_0_001000010000;
      patterns[2115] = 29'b0_000100001000_011_0_010000100000;
      patterns[2116] = 29'b0_000100001000_100_0_000010000100;
      patterns[2117] = 29'b0_000100001000_101_0_000001000010;
      patterns[2118] = 29'b0_000100001000_110_0_000100001000;
      patterns[2119] = 29'b0_000100001000_111_0_000100001000;
      patterns[2120] = 29'b0_000100001001_000_0_000100001001;
      patterns[2121] = 29'b0_000100001001_001_0_001001000100;
      patterns[2122] = 29'b0_000100001001_010_0_001000010010;
      patterns[2123] = 29'b0_000100001001_011_0_010000100100;
      patterns[2124] = 29'b0_000100001001_100_1_000010000100;
      patterns[2125] = 29'b0_000100001001_101_0_100001000010;
      patterns[2126] = 29'b0_000100001001_110_0_000100001001;
      patterns[2127] = 29'b0_000100001001_111_0_000100001001;
      patterns[2128] = 29'b0_000100001010_000_0_000100001010;
      patterns[2129] = 29'b0_000100001010_001_0_001010000100;
      patterns[2130] = 29'b0_000100001010_010_0_001000010100;
      patterns[2131] = 29'b0_000100001010_011_0_010000101000;
      patterns[2132] = 29'b0_000100001010_100_0_000010000101;
      patterns[2133] = 29'b0_000100001010_101_1_000001000010;
      patterns[2134] = 29'b0_000100001010_110_0_000100001010;
      patterns[2135] = 29'b0_000100001010_111_0_000100001010;
      patterns[2136] = 29'b0_000100001011_000_0_000100001011;
      patterns[2137] = 29'b0_000100001011_001_0_001011000100;
      patterns[2138] = 29'b0_000100001011_010_0_001000010110;
      patterns[2139] = 29'b0_000100001011_011_0_010000101100;
      patterns[2140] = 29'b0_000100001011_100_1_000010000101;
      patterns[2141] = 29'b0_000100001011_101_1_100001000010;
      patterns[2142] = 29'b0_000100001011_110_0_000100001011;
      patterns[2143] = 29'b0_000100001011_111_0_000100001011;
      patterns[2144] = 29'b0_000100001100_000_0_000100001100;
      patterns[2145] = 29'b0_000100001100_001_0_001100000100;
      patterns[2146] = 29'b0_000100001100_010_0_001000011000;
      patterns[2147] = 29'b0_000100001100_011_0_010000110000;
      patterns[2148] = 29'b0_000100001100_100_0_000010000110;
      patterns[2149] = 29'b0_000100001100_101_0_000001000011;
      patterns[2150] = 29'b0_000100001100_110_0_000100001100;
      patterns[2151] = 29'b0_000100001100_111_0_000100001100;
      patterns[2152] = 29'b0_000100001101_000_0_000100001101;
      patterns[2153] = 29'b0_000100001101_001_0_001101000100;
      patterns[2154] = 29'b0_000100001101_010_0_001000011010;
      patterns[2155] = 29'b0_000100001101_011_0_010000110100;
      patterns[2156] = 29'b0_000100001101_100_1_000010000110;
      patterns[2157] = 29'b0_000100001101_101_0_100001000011;
      patterns[2158] = 29'b0_000100001101_110_0_000100001101;
      patterns[2159] = 29'b0_000100001101_111_0_000100001101;
      patterns[2160] = 29'b0_000100001110_000_0_000100001110;
      patterns[2161] = 29'b0_000100001110_001_0_001110000100;
      patterns[2162] = 29'b0_000100001110_010_0_001000011100;
      patterns[2163] = 29'b0_000100001110_011_0_010000111000;
      patterns[2164] = 29'b0_000100001110_100_0_000010000111;
      patterns[2165] = 29'b0_000100001110_101_1_000001000011;
      patterns[2166] = 29'b0_000100001110_110_0_000100001110;
      patterns[2167] = 29'b0_000100001110_111_0_000100001110;
      patterns[2168] = 29'b0_000100001111_000_0_000100001111;
      patterns[2169] = 29'b0_000100001111_001_0_001111000100;
      patterns[2170] = 29'b0_000100001111_010_0_001000011110;
      patterns[2171] = 29'b0_000100001111_011_0_010000111100;
      patterns[2172] = 29'b0_000100001111_100_1_000010000111;
      patterns[2173] = 29'b0_000100001111_101_1_100001000011;
      patterns[2174] = 29'b0_000100001111_110_0_000100001111;
      patterns[2175] = 29'b0_000100001111_111_0_000100001111;
      patterns[2176] = 29'b0_000100010000_000_0_000100010000;
      patterns[2177] = 29'b0_000100010000_001_0_010000000100;
      patterns[2178] = 29'b0_000100010000_010_0_001000100000;
      patterns[2179] = 29'b0_000100010000_011_0_010001000000;
      patterns[2180] = 29'b0_000100010000_100_0_000010001000;
      patterns[2181] = 29'b0_000100010000_101_0_000001000100;
      patterns[2182] = 29'b0_000100010000_110_0_000100010000;
      patterns[2183] = 29'b0_000100010000_111_0_000100010000;
      patterns[2184] = 29'b0_000100010001_000_0_000100010001;
      patterns[2185] = 29'b0_000100010001_001_0_010001000100;
      patterns[2186] = 29'b0_000100010001_010_0_001000100010;
      patterns[2187] = 29'b0_000100010001_011_0_010001000100;
      patterns[2188] = 29'b0_000100010001_100_1_000010001000;
      patterns[2189] = 29'b0_000100010001_101_0_100001000100;
      patterns[2190] = 29'b0_000100010001_110_0_000100010001;
      patterns[2191] = 29'b0_000100010001_111_0_000100010001;
      patterns[2192] = 29'b0_000100010010_000_0_000100010010;
      patterns[2193] = 29'b0_000100010010_001_0_010010000100;
      patterns[2194] = 29'b0_000100010010_010_0_001000100100;
      patterns[2195] = 29'b0_000100010010_011_0_010001001000;
      patterns[2196] = 29'b0_000100010010_100_0_000010001001;
      patterns[2197] = 29'b0_000100010010_101_1_000001000100;
      patterns[2198] = 29'b0_000100010010_110_0_000100010010;
      patterns[2199] = 29'b0_000100010010_111_0_000100010010;
      patterns[2200] = 29'b0_000100010011_000_0_000100010011;
      patterns[2201] = 29'b0_000100010011_001_0_010011000100;
      patterns[2202] = 29'b0_000100010011_010_0_001000100110;
      patterns[2203] = 29'b0_000100010011_011_0_010001001100;
      patterns[2204] = 29'b0_000100010011_100_1_000010001001;
      patterns[2205] = 29'b0_000100010011_101_1_100001000100;
      patterns[2206] = 29'b0_000100010011_110_0_000100010011;
      patterns[2207] = 29'b0_000100010011_111_0_000100010011;
      patterns[2208] = 29'b0_000100010100_000_0_000100010100;
      patterns[2209] = 29'b0_000100010100_001_0_010100000100;
      patterns[2210] = 29'b0_000100010100_010_0_001000101000;
      patterns[2211] = 29'b0_000100010100_011_0_010001010000;
      patterns[2212] = 29'b0_000100010100_100_0_000010001010;
      patterns[2213] = 29'b0_000100010100_101_0_000001000101;
      patterns[2214] = 29'b0_000100010100_110_0_000100010100;
      patterns[2215] = 29'b0_000100010100_111_0_000100010100;
      patterns[2216] = 29'b0_000100010101_000_0_000100010101;
      patterns[2217] = 29'b0_000100010101_001_0_010101000100;
      patterns[2218] = 29'b0_000100010101_010_0_001000101010;
      patterns[2219] = 29'b0_000100010101_011_0_010001010100;
      patterns[2220] = 29'b0_000100010101_100_1_000010001010;
      patterns[2221] = 29'b0_000100010101_101_0_100001000101;
      patterns[2222] = 29'b0_000100010101_110_0_000100010101;
      patterns[2223] = 29'b0_000100010101_111_0_000100010101;
      patterns[2224] = 29'b0_000100010110_000_0_000100010110;
      patterns[2225] = 29'b0_000100010110_001_0_010110000100;
      patterns[2226] = 29'b0_000100010110_010_0_001000101100;
      patterns[2227] = 29'b0_000100010110_011_0_010001011000;
      patterns[2228] = 29'b0_000100010110_100_0_000010001011;
      patterns[2229] = 29'b0_000100010110_101_1_000001000101;
      patterns[2230] = 29'b0_000100010110_110_0_000100010110;
      patterns[2231] = 29'b0_000100010110_111_0_000100010110;
      patterns[2232] = 29'b0_000100010111_000_0_000100010111;
      patterns[2233] = 29'b0_000100010111_001_0_010111000100;
      patterns[2234] = 29'b0_000100010111_010_0_001000101110;
      patterns[2235] = 29'b0_000100010111_011_0_010001011100;
      patterns[2236] = 29'b0_000100010111_100_1_000010001011;
      patterns[2237] = 29'b0_000100010111_101_1_100001000101;
      patterns[2238] = 29'b0_000100010111_110_0_000100010111;
      patterns[2239] = 29'b0_000100010111_111_0_000100010111;
      patterns[2240] = 29'b0_000100011000_000_0_000100011000;
      patterns[2241] = 29'b0_000100011000_001_0_011000000100;
      patterns[2242] = 29'b0_000100011000_010_0_001000110000;
      patterns[2243] = 29'b0_000100011000_011_0_010001100000;
      patterns[2244] = 29'b0_000100011000_100_0_000010001100;
      patterns[2245] = 29'b0_000100011000_101_0_000001000110;
      patterns[2246] = 29'b0_000100011000_110_0_000100011000;
      patterns[2247] = 29'b0_000100011000_111_0_000100011000;
      patterns[2248] = 29'b0_000100011001_000_0_000100011001;
      patterns[2249] = 29'b0_000100011001_001_0_011001000100;
      patterns[2250] = 29'b0_000100011001_010_0_001000110010;
      patterns[2251] = 29'b0_000100011001_011_0_010001100100;
      patterns[2252] = 29'b0_000100011001_100_1_000010001100;
      patterns[2253] = 29'b0_000100011001_101_0_100001000110;
      patterns[2254] = 29'b0_000100011001_110_0_000100011001;
      patterns[2255] = 29'b0_000100011001_111_0_000100011001;
      patterns[2256] = 29'b0_000100011010_000_0_000100011010;
      patterns[2257] = 29'b0_000100011010_001_0_011010000100;
      patterns[2258] = 29'b0_000100011010_010_0_001000110100;
      patterns[2259] = 29'b0_000100011010_011_0_010001101000;
      patterns[2260] = 29'b0_000100011010_100_0_000010001101;
      patterns[2261] = 29'b0_000100011010_101_1_000001000110;
      patterns[2262] = 29'b0_000100011010_110_0_000100011010;
      patterns[2263] = 29'b0_000100011010_111_0_000100011010;
      patterns[2264] = 29'b0_000100011011_000_0_000100011011;
      patterns[2265] = 29'b0_000100011011_001_0_011011000100;
      patterns[2266] = 29'b0_000100011011_010_0_001000110110;
      patterns[2267] = 29'b0_000100011011_011_0_010001101100;
      patterns[2268] = 29'b0_000100011011_100_1_000010001101;
      patterns[2269] = 29'b0_000100011011_101_1_100001000110;
      patterns[2270] = 29'b0_000100011011_110_0_000100011011;
      patterns[2271] = 29'b0_000100011011_111_0_000100011011;
      patterns[2272] = 29'b0_000100011100_000_0_000100011100;
      patterns[2273] = 29'b0_000100011100_001_0_011100000100;
      patterns[2274] = 29'b0_000100011100_010_0_001000111000;
      patterns[2275] = 29'b0_000100011100_011_0_010001110000;
      patterns[2276] = 29'b0_000100011100_100_0_000010001110;
      patterns[2277] = 29'b0_000100011100_101_0_000001000111;
      patterns[2278] = 29'b0_000100011100_110_0_000100011100;
      patterns[2279] = 29'b0_000100011100_111_0_000100011100;
      patterns[2280] = 29'b0_000100011101_000_0_000100011101;
      patterns[2281] = 29'b0_000100011101_001_0_011101000100;
      patterns[2282] = 29'b0_000100011101_010_0_001000111010;
      patterns[2283] = 29'b0_000100011101_011_0_010001110100;
      patterns[2284] = 29'b0_000100011101_100_1_000010001110;
      patterns[2285] = 29'b0_000100011101_101_0_100001000111;
      patterns[2286] = 29'b0_000100011101_110_0_000100011101;
      patterns[2287] = 29'b0_000100011101_111_0_000100011101;
      patterns[2288] = 29'b0_000100011110_000_0_000100011110;
      patterns[2289] = 29'b0_000100011110_001_0_011110000100;
      patterns[2290] = 29'b0_000100011110_010_0_001000111100;
      patterns[2291] = 29'b0_000100011110_011_0_010001111000;
      patterns[2292] = 29'b0_000100011110_100_0_000010001111;
      patterns[2293] = 29'b0_000100011110_101_1_000001000111;
      patterns[2294] = 29'b0_000100011110_110_0_000100011110;
      patterns[2295] = 29'b0_000100011110_111_0_000100011110;
      patterns[2296] = 29'b0_000100011111_000_0_000100011111;
      patterns[2297] = 29'b0_000100011111_001_0_011111000100;
      patterns[2298] = 29'b0_000100011111_010_0_001000111110;
      patterns[2299] = 29'b0_000100011111_011_0_010001111100;
      patterns[2300] = 29'b0_000100011111_100_1_000010001111;
      patterns[2301] = 29'b0_000100011111_101_1_100001000111;
      patterns[2302] = 29'b0_000100011111_110_0_000100011111;
      patterns[2303] = 29'b0_000100011111_111_0_000100011111;
      patterns[2304] = 29'b0_000100100000_000_0_000100100000;
      patterns[2305] = 29'b0_000100100000_001_0_100000000100;
      patterns[2306] = 29'b0_000100100000_010_0_001001000000;
      patterns[2307] = 29'b0_000100100000_011_0_010010000000;
      patterns[2308] = 29'b0_000100100000_100_0_000010010000;
      patterns[2309] = 29'b0_000100100000_101_0_000001001000;
      patterns[2310] = 29'b0_000100100000_110_0_000100100000;
      patterns[2311] = 29'b0_000100100000_111_0_000100100000;
      patterns[2312] = 29'b0_000100100001_000_0_000100100001;
      patterns[2313] = 29'b0_000100100001_001_0_100001000100;
      patterns[2314] = 29'b0_000100100001_010_0_001001000010;
      patterns[2315] = 29'b0_000100100001_011_0_010010000100;
      patterns[2316] = 29'b0_000100100001_100_1_000010010000;
      patterns[2317] = 29'b0_000100100001_101_0_100001001000;
      patterns[2318] = 29'b0_000100100001_110_0_000100100001;
      patterns[2319] = 29'b0_000100100001_111_0_000100100001;
      patterns[2320] = 29'b0_000100100010_000_0_000100100010;
      patterns[2321] = 29'b0_000100100010_001_0_100010000100;
      patterns[2322] = 29'b0_000100100010_010_0_001001000100;
      patterns[2323] = 29'b0_000100100010_011_0_010010001000;
      patterns[2324] = 29'b0_000100100010_100_0_000010010001;
      patterns[2325] = 29'b0_000100100010_101_1_000001001000;
      patterns[2326] = 29'b0_000100100010_110_0_000100100010;
      patterns[2327] = 29'b0_000100100010_111_0_000100100010;
      patterns[2328] = 29'b0_000100100011_000_0_000100100011;
      patterns[2329] = 29'b0_000100100011_001_0_100011000100;
      patterns[2330] = 29'b0_000100100011_010_0_001001000110;
      patterns[2331] = 29'b0_000100100011_011_0_010010001100;
      patterns[2332] = 29'b0_000100100011_100_1_000010010001;
      patterns[2333] = 29'b0_000100100011_101_1_100001001000;
      patterns[2334] = 29'b0_000100100011_110_0_000100100011;
      patterns[2335] = 29'b0_000100100011_111_0_000100100011;
      patterns[2336] = 29'b0_000100100100_000_0_000100100100;
      patterns[2337] = 29'b0_000100100100_001_0_100100000100;
      patterns[2338] = 29'b0_000100100100_010_0_001001001000;
      patterns[2339] = 29'b0_000100100100_011_0_010010010000;
      patterns[2340] = 29'b0_000100100100_100_0_000010010010;
      patterns[2341] = 29'b0_000100100100_101_0_000001001001;
      patterns[2342] = 29'b0_000100100100_110_0_000100100100;
      patterns[2343] = 29'b0_000100100100_111_0_000100100100;
      patterns[2344] = 29'b0_000100100101_000_0_000100100101;
      patterns[2345] = 29'b0_000100100101_001_0_100101000100;
      patterns[2346] = 29'b0_000100100101_010_0_001001001010;
      patterns[2347] = 29'b0_000100100101_011_0_010010010100;
      patterns[2348] = 29'b0_000100100101_100_1_000010010010;
      patterns[2349] = 29'b0_000100100101_101_0_100001001001;
      patterns[2350] = 29'b0_000100100101_110_0_000100100101;
      patterns[2351] = 29'b0_000100100101_111_0_000100100101;
      patterns[2352] = 29'b0_000100100110_000_0_000100100110;
      patterns[2353] = 29'b0_000100100110_001_0_100110000100;
      patterns[2354] = 29'b0_000100100110_010_0_001001001100;
      patterns[2355] = 29'b0_000100100110_011_0_010010011000;
      patterns[2356] = 29'b0_000100100110_100_0_000010010011;
      patterns[2357] = 29'b0_000100100110_101_1_000001001001;
      patterns[2358] = 29'b0_000100100110_110_0_000100100110;
      patterns[2359] = 29'b0_000100100110_111_0_000100100110;
      patterns[2360] = 29'b0_000100100111_000_0_000100100111;
      patterns[2361] = 29'b0_000100100111_001_0_100111000100;
      patterns[2362] = 29'b0_000100100111_010_0_001001001110;
      patterns[2363] = 29'b0_000100100111_011_0_010010011100;
      patterns[2364] = 29'b0_000100100111_100_1_000010010011;
      patterns[2365] = 29'b0_000100100111_101_1_100001001001;
      patterns[2366] = 29'b0_000100100111_110_0_000100100111;
      patterns[2367] = 29'b0_000100100111_111_0_000100100111;
      patterns[2368] = 29'b0_000100101000_000_0_000100101000;
      patterns[2369] = 29'b0_000100101000_001_0_101000000100;
      patterns[2370] = 29'b0_000100101000_010_0_001001010000;
      patterns[2371] = 29'b0_000100101000_011_0_010010100000;
      patterns[2372] = 29'b0_000100101000_100_0_000010010100;
      patterns[2373] = 29'b0_000100101000_101_0_000001001010;
      patterns[2374] = 29'b0_000100101000_110_0_000100101000;
      patterns[2375] = 29'b0_000100101000_111_0_000100101000;
      patterns[2376] = 29'b0_000100101001_000_0_000100101001;
      patterns[2377] = 29'b0_000100101001_001_0_101001000100;
      patterns[2378] = 29'b0_000100101001_010_0_001001010010;
      patterns[2379] = 29'b0_000100101001_011_0_010010100100;
      patterns[2380] = 29'b0_000100101001_100_1_000010010100;
      patterns[2381] = 29'b0_000100101001_101_0_100001001010;
      patterns[2382] = 29'b0_000100101001_110_0_000100101001;
      patterns[2383] = 29'b0_000100101001_111_0_000100101001;
      patterns[2384] = 29'b0_000100101010_000_0_000100101010;
      patterns[2385] = 29'b0_000100101010_001_0_101010000100;
      patterns[2386] = 29'b0_000100101010_010_0_001001010100;
      patterns[2387] = 29'b0_000100101010_011_0_010010101000;
      patterns[2388] = 29'b0_000100101010_100_0_000010010101;
      patterns[2389] = 29'b0_000100101010_101_1_000001001010;
      patterns[2390] = 29'b0_000100101010_110_0_000100101010;
      patterns[2391] = 29'b0_000100101010_111_0_000100101010;
      patterns[2392] = 29'b0_000100101011_000_0_000100101011;
      patterns[2393] = 29'b0_000100101011_001_0_101011000100;
      patterns[2394] = 29'b0_000100101011_010_0_001001010110;
      patterns[2395] = 29'b0_000100101011_011_0_010010101100;
      patterns[2396] = 29'b0_000100101011_100_1_000010010101;
      patterns[2397] = 29'b0_000100101011_101_1_100001001010;
      patterns[2398] = 29'b0_000100101011_110_0_000100101011;
      patterns[2399] = 29'b0_000100101011_111_0_000100101011;
      patterns[2400] = 29'b0_000100101100_000_0_000100101100;
      patterns[2401] = 29'b0_000100101100_001_0_101100000100;
      patterns[2402] = 29'b0_000100101100_010_0_001001011000;
      patterns[2403] = 29'b0_000100101100_011_0_010010110000;
      patterns[2404] = 29'b0_000100101100_100_0_000010010110;
      patterns[2405] = 29'b0_000100101100_101_0_000001001011;
      patterns[2406] = 29'b0_000100101100_110_0_000100101100;
      patterns[2407] = 29'b0_000100101100_111_0_000100101100;
      patterns[2408] = 29'b0_000100101101_000_0_000100101101;
      patterns[2409] = 29'b0_000100101101_001_0_101101000100;
      patterns[2410] = 29'b0_000100101101_010_0_001001011010;
      patterns[2411] = 29'b0_000100101101_011_0_010010110100;
      patterns[2412] = 29'b0_000100101101_100_1_000010010110;
      patterns[2413] = 29'b0_000100101101_101_0_100001001011;
      patterns[2414] = 29'b0_000100101101_110_0_000100101101;
      patterns[2415] = 29'b0_000100101101_111_0_000100101101;
      patterns[2416] = 29'b0_000100101110_000_0_000100101110;
      patterns[2417] = 29'b0_000100101110_001_0_101110000100;
      patterns[2418] = 29'b0_000100101110_010_0_001001011100;
      patterns[2419] = 29'b0_000100101110_011_0_010010111000;
      patterns[2420] = 29'b0_000100101110_100_0_000010010111;
      patterns[2421] = 29'b0_000100101110_101_1_000001001011;
      patterns[2422] = 29'b0_000100101110_110_0_000100101110;
      patterns[2423] = 29'b0_000100101110_111_0_000100101110;
      patterns[2424] = 29'b0_000100101111_000_0_000100101111;
      patterns[2425] = 29'b0_000100101111_001_0_101111000100;
      patterns[2426] = 29'b0_000100101111_010_0_001001011110;
      patterns[2427] = 29'b0_000100101111_011_0_010010111100;
      patterns[2428] = 29'b0_000100101111_100_1_000010010111;
      patterns[2429] = 29'b0_000100101111_101_1_100001001011;
      patterns[2430] = 29'b0_000100101111_110_0_000100101111;
      patterns[2431] = 29'b0_000100101111_111_0_000100101111;
      patterns[2432] = 29'b0_000100110000_000_0_000100110000;
      patterns[2433] = 29'b0_000100110000_001_0_110000000100;
      patterns[2434] = 29'b0_000100110000_010_0_001001100000;
      patterns[2435] = 29'b0_000100110000_011_0_010011000000;
      patterns[2436] = 29'b0_000100110000_100_0_000010011000;
      patterns[2437] = 29'b0_000100110000_101_0_000001001100;
      patterns[2438] = 29'b0_000100110000_110_0_000100110000;
      patterns[2439] = 29'b0_000100110000_111_0_000100110000;
      patterns[2440] = 29'b0_000100110001_000_0_000100110001;
      patterns[2441] = 29'b0_000100110001_001_0_110001000100;
      patterns[2442] = 29'b0_000100110001_010_0_001001100010;
      patterns[2443] = 29'b0_000100110001_011_0_010011000100;
      patterns[2444] = 29'b0_000100110001_100_1_000010011000;
      patterns[2445] = 29'b0_000100110001_101_0_100001001100;
      patterns[2446] = 29'b0_000100110001_110_0_000100110001;
      patterns[2447] = 29'b0_000100110001_111_0_000100110001;
      patterns[2448] = 29'b0_000100110010_000_0_000100110010;
      patterns[2449] = 29'b0_000100110010_001_0_110010000100;
      patterns[2450] = 29'b0_000100110010_010_0_001001100100;
      patterns[2451] = 29'b0_000100110010_011_0_010011001000;
      patterns[2452] = 29'b0_000100110010_100_0_000010011001;
      patterns[2453] = 29'b0_000100110010_101_1_000001001100;
      patterns[2454] = 29'b0_000100110010_110_0_000100110010;
      patterns[2455] = 29'b0_000100110010_111_0_000100110010;
      patterns[2456] = 29'b0_000100110011_000_0_000100110011;
      patterns[2457] = 29'b0_000100110011_001_0_110011000100;
      patterns[2458] = 29'b0_000100110011_010_0_001001100110;
      patterns[2459] = 29'b0_000100110011_011_0_010011001100;
      patterns[2460] = 29'b0_000100110011_100_1_000010011001;
      patterns[2461] = 29'b0_000100110011_101_1_100001001100;
      patterns[2462] = 29'b0_000100110011_110_0_000100110011;
      patterns[2463] = 29'b0_000100110011_111_0_000100110011;
      patterns[2464] = 29'b0_000100110100_000_0_000100110100;
      patterns[2465] = 29'b0_000100110100_001_0_110100000100;
      patterns[2466] = 29'b0_000100110100_010_0_001001101000;
      patterns[2467] = 29'b0_000100110100_011_0_010011010000;
      patterns[2468] = 29'b0_000100110100_100_0_000010011010;
      patterns[2469] = 29'b0_000100110100_101_0_000001001101;
      patterns[2470] = 29'b0_000100110100_110_0_000100110100;
      patterns[2471] = 29'b0_000100110100_111_0_000100110100;
      patterns[2472] = 29'b0_000100110101_000_0_000100110101;
      patterns[2473] = 29'b0_000100110101_001_0_110101000100;
      patterns[2474] = 29'b0_000100110101_010_0_001001101010;
      patterns[2475] = 29'b0_000100110101_011_0_010011010100;
      patterns[2476] = 29'b0_000100110101_100_1_000010011010;
      patterns[2477] = 29'b0_000100110101_101_0_100001001101;
      patterns[2478] = 29'b0_000100110101_110_0_000100110101;
      patterns[2479] = 29'b0_000100110101_111_0_000100110101;
      patterns[2480] = 29'b0_000100110110_000_0_000100110110;
      patterns[2481] = 29'b0_000100110110_001_0_110110000100;
      patterns[2482] = 29'b0_000100110110_010_0_001001101100;
      patterns[2483] = 29'b0_000100110110_011_0_010011011000;
      patterns[2484] = 29'b0_000100110110_100_0_000010011011;
      patterns[2485] = 29'b0_000100110110_101_1_000001001101;
      patterns[2486] = 29'b0_000100110110_110_0_000100110110;
      patterns[2487] = 29'b0_000100110110_111_0_000100110110;
      patterns[2488] = 29'b0_000100110111_000_0_000100110111;
      patterns[2489] = 29'b0_000100110111_001_0_110111000100;
      patterns[2490] = 29'b0_000100110111_010_0_001001101110;
      patterns[2491] = 29'b0_000100110111_011_0_010011011100;
      patterns[2492] = 29'b0_000100110111_100_1_000010011011;
      patterns[2493] = 29'b0_000100110111_101_1_100001001101;
      patterns[2494] = 29'b0_000100110111_110_0_000100110111;
      patterns[2495] = 29'b0_000100110111_111_0_000100110111;
      patterns[2496] = 29'b0_000100111000_000_0_000100111000;
      patterns[2497] = 29'b0_000100111000_001_0_111000000100;
      patterns[2498] = 29'b0_000100111000_010_0_001001110000;
      patterns[2499] = 29'b0_000100111000_011_0_010011100000;
      patterns[2500] = 29'b0_000100111000_100_0_000010011100;
      patterns[2501] = 29'b0_000100111000_101_0_000001001110;
      patterns[2502] = 29'b0_000100111000_110_0_000100111000;
      patterns[2503] = 29'b0_000100111000_111_0_000100111000;
      patterns[2504] = 29'b0_000100111001_000_0_000100111001;
      patterns[2505] = 29'b0_000100111001_001_0_111001000100;
      patterns[2506] = 29'b0_000100111001_010_0_001001110010;
      patterns[2507] = 29'b0_000100111001_011_0_010011100100;
      patterns[2508] = 29'b0_000100111001_100_1_000010011100;
      patterns[2509] = 29'b0_000100111001_101_0_100001001110;
      patterns[2510] = 29'b0_000100111001_110_0_000100111001;
      patterns[2511] = 29'b0_000100111001_111_0_000100111001;
      patterns[2512] = 29'b0_000100111010_000_0_000100111010;
      patterns[2513] = 29'b0_000100111010_001_0_111010000100;
      patterns[2514] = 29'b0_000100111010_010_0_001001110100;
      patterns[2515] = 29'b0_000100111010_011_0_010011101000;
      patterns[2516] = 29'b0_000100111010_100_0_000010011101;
      patterns[2517] = 29'b0_000100111010_101_1_000001001110;
      patterns[2518] = 29'b0_000100111010_110_0_000100111010;
      patterns[2519] = 29'b0_000100111010_111_0_000100111010;
      patterns[2520] = 29'b0_000100111011_000_0_000100111011;
      patterns[2521] = 29'b0_000100111011_001_0_111011000100;
      patterns[2522] = 29'b0_000100111011_010_0_001001110110;
      patterns[2523] = 29'b0_000100111011_011_0_010011101100;
      patterns[2524] = 29'b0_000100111011_100_1_000010011101;
      patterns[2525] = 29'b0_000100111011_101_1_100001001110;
      patterns[2526] = 29'b0_000100111011_110_0_000100111011;
      patterns[2527] = 29'b0_000100111011_111_0_000100111011;
      patterns[2528] = 29'b0_000100111100_000_0_000100111100;
      patterns[2529] = 29'b0_000100111100_001_0_111100000100;
      patterns[2530] = 29'b0_000100111100_010_0_001001111000;
      patterns[2531] = 29'b0_000100111100_011_0_010011110000;
      patterns[2532] = 29'b0_000100111100_100_0_000010011110;
      patterns[2533] = 29'b0_000100111100_101_0_000001001111;
      patterns[2534] = 29'b0_000100111100_110_0_000100111100;
      patterns[2535] = 29'b0_000100111100_111_0_000100111100;
      patterns[2536] = 29'b0_000100111101_000_0_000100111101;
      patterns[2537] = 29'b0_000100111101_001_0_111101000100;
      patterns[2538] = 29'b0_000100111101_010_0_001001111010;
      patterns[2539] = 29'b0_000100111101_011_0_010011110100;
      patterns[2540] = 29'b0_000100111101_100_1_000010011110;
      patterns[2541] = 29'b0_000100111101_101_0_100001001111;
      patterns[2542] = 29'b0_000100111101_110_0_000100111101;
      patterns[2543] = 29'b0_000100111101_111_0_000100111101;
      patterns[2544] = 29'b0_000100111110_000_0_000100111110;
      patterns[2545] = 29'b0_000100111110_001_0_111110000100;
      patterns[2546] = 29'b0_000100111110_010_0_001001111100;
      patterns[2547] = 29'b0_000100111110_011_0_010011111000;
      patterns[2548] = 29'b0_000100111110_100_0_000010011111;
      patterns[2549] = 29'b0_000100111110_101_1_000001001111;
      patterns[2550] = 29'b0_000100111110_110_0_000100111110;
      patterns[2551] = 29'b0_000100111110_111_0_000100111110;
      patterns[2552] = 29'b0_000100111111_000_0_000100111111;
      patterns[2553] = 29'b0_000100111111_001_0_111111000100;
      patterns[2554] = 29'b0_000100111111_010_0_001001111110;
      patterns[2555] = 29'b0_000100111111_011_0_010011111100;
      patterns[2556] = 29'b0_000100111111_100_1_000010011111;
      patterns[2557] = 29'b0_000100111111_101_1_100001001111;
      patterns[2558] = 29'b0_000100111111_110_0_000100111111;
      patterns[2559] = 29'b0_000100111111_111_0_000100111111;
      patterns[2560] = 29'b0_000101000000_000_0_000101000000;
      patterns[2561] = 29'b0_000101000000_001_0_000000000101;
      patterns[2562] = 29'b0_000101000000_010_0_001010000000;
      patterns[2563] = 29'b0_000101000000_011_0_010100000000;
      patterns[2564] = 29'b0_000101000000_100_0_000010100000;
      patterns[2565] = 29'b0_000101000000_101_0_000001010000;
      patterns[2566] = 29'b0_000101000000_110_0_000101000000;
      patterns[2567] = 29'b0_000101000000_111_0_000101000000;
      patterns[2568] = 29'b0_000101000001_000_0_000101000001;
      patterns[2569] = 29'b0_000101000001_001_0_000001000101;
      patterns[2570] = 29'b0_000101000001_010_0_001010000010;
      patterns[2571] = 29'b0_000101000001_011_0_010100000100;
      patterns[2572] = 29'b0_000101000001_100_1_000010100000;
      patterns[2573] = 29'b0_000101000001_101_0_100001010000;
      patterns[2574] = 29'b0_000101000001_110_0_000101000001;
      patterns[2575] = 29'b0_000101000001_111_0_000101000001;
      patterns[2576] = 29'b0_000101000010_000_0_000101000010;
      patterns[2577] = 29'b0_000101000010_001_0_000010000101;
      patterns[2578] = 29'b0_000101000010_010_0_001010000100;
      patterns[2579] = 29'b0_000101000010_011_0_010100001000;
      patterns[2580] = 29'b0_000101000010_100_0_000010100001;
      patterns[2581] = 29'b0_000101000010_101_1_000001010000;
      patterns[2582] = 29'b0_000101000010_110_0_000101000010;
      patterns[2583] = 29'b0_000101000010_111_0_000101000010;
      patterns[2584] = 29'b0_000101000011_000_0_000101000011;
      patterns[2585] = 29'b0_000101000011_001_0_000011000101;
      patterns[2586] = 29'b0_000101000011_010_0_001010000110;
      patterns[2587] = 29'b0_000101000011_011_0_010100001100;
      patterns[2588] = 29'b0_000101000011_100_1_000010100001;
      patterns[2589] = 29'b0_000101000011_101_1_100001010000;
      patterns[2590] = 29'b0_000101000011_110_0_000101000011;
      patterns[2591] = 29'b0_000101000011_111_0_000101000011;
      patterns[2592] = 29'b0_000101000100_000_0_000101000100;
      patterns[2593] = 29'b0_000101000100_001_0_000100000101;
      patterns[2594] = 29'b0_000101000100_010_0_001010001000;
      patterns[2595] = 29'b0_000101000100_011_0_010100010000;
      patterns[2596] = 29'b0_000101000100_100_0_000010100010;
      patterns[2597] = 29'b0_000101000100_101_0_000001010001;
      patterns[2598] = 29'b0_000101000100_110_0_000101000100;
      patterns[2599] = 29'b0_000101000100_111_0_000101000100;
      patterns[2600] = 29'b0_000101000101_000_0_000101000101;
      patterns[2601] = 29'b0_000101000101_001_0_000101000101;
      patterns[2602] = 29'b0_000101000101_010_0_001010001010;
      patterns[2603] = 29'b0_000101000101_011_0_010100010100;
      patterns[2604] = 29'b0_000101000101_100_1_000010100010;
      patterns[2605] = 29'b0_000101000101_101_0_100001010001;
      patterns[2606] = 29'b0_000101000101_110_0_000101000101;
      patterns[2607] = 29'b0_000101000101_111_0_000101000101;
      patterns[2608] = 29'b0_000101000110_000_0_000101000110;
      patterns[2609] = 29'b0_000101000110_001_0_000110000101;
      patterns[2610] = 29'b0_000101000110_010_0_001010001100;
      patterns[2611] = 29'b0_000101000110_011_0_010100011000;
      patterns[2612] = 29'b0_000101000110_100_0_000010100011;
      patterns[2613] = 29'b0_000101000110_101_1_000001010001;
      patterns[2614] = 29'b0_000101000110_110_0_000101000110;
      patterns[2615] = 29'b0_000101000110_111_0_000101000110;
      patterns[2616] = 29'b0_000101000111_000_0_000101000111;
      patterns[2617] = 29'b0_000101000111_001_0_000111000101;
      patterns[2618] = 29'b0_000101000111_010_0_001010001110;
      patterns[2619] = 29'b0_000101000111_011_0_010100011100;
      patterns[2620] = 29'b0_000101000111_100_1_000010100011;
      patterns[2621] = 29'b0_000101000111_101_1_100001010001;
      patterns[2622] = 29'b0_000101000111_110_0_000101000111;
      patterns[2623] = 29'b0_000101000111_111_0_000101000111;
      patterns[2624] = 29'b0_000101001000_000_0_000101001000;
      patterns[2625] = 29'b0_000101001000_001_0_001000000101;
      patterns[2626] = 29'b0_000101001000_010_0_001010010000;
      patterns[2627] = 29'b0_000101001000_011_0_010100100000;
      patterns[2628] = 29'b0_000101001000_100_0_000010100100;
      patterns[2629] = 29'b0_000101001000_101_0_000001010010;
      patterns[2630] = 29'b0_000101001000_110_0_000101001000;
      patterns[2631] = 29'b0_000101001000_111_0_000101001000;
      patterns[2632] = 29'b0_000101001001_000_0_000101001001;
      patterns[2633] = 29'b0_000101001001_001_0_001001000101;
      patterns[2634] = 29'b0_000101001001_010_0_001010010010;
      patterns[2635] = 29'b0_000101001001_011_0_010100100100;
      patterns[2636] = 29'b0_000101001001_100_1_000010100100;
      patterns[2637] = 29'b0_000101001001_101_0_100001010010;
      patterns[2638] = 29'b0_000101001001_110_0_000101001001;
      patterns[2639] = 29'b0_000101001001_111_0_000101001001;
      patterns[2640] = 29'b0_000101001010_000_0_000101001010;
      patterns[2641] = 29'b0_000101001010_001_0_001010000101;
      patterns[2642] = 29'b0_000101001010_010_0_001010010100;
      patterns[2643] = 29'b0_000101001010_011_0_010100101000;
      patterns[2644] = 29'b0_000101001010_100_0_000010100101;
      patterns[2645] = 29'b0_000101001010_101_1_000001010010;
      patterns[2646] = 29'b0_000101001010_110_0_000101001010;
      patterns[2647] = 29'b0_000101001010_111_0_000101001010;
      patterns[2648] = 29'b0_000101001011_000_0_000101001011;
      patterns[2649] = 29'b0_000101001011_001_0_001011000101;
      patterns[2650] = 29'b0_000101001011_010_0_001010010110;
      patterns[2651] = 29'b0_000101001011_011_0_010100101100;
      patterns[2652] = 29'b0_000101001011_100_1_000010100101;
      patterns[2653] = 29'b0_000101001011_101_1_100001010010;
      patterns[2654] = 29'b0_000101001011_110_0_000101001011;
      patterns[2655] = 29'b0_000101001011_111_0_000101001011;
      patterns[2656] = 29'b0_000101001100_000_0_000101001100;
      patterns[2657] = 29'b0_000101001100_001_0_001100000101;
      patterns[2658] = 29'b0_000101001100_010_0_001010011000;
      patterns[2659] = 29'b0_000101001100_011_0_010100110000;
      patterns[2660] = 29'b0_000101001100_100_0_000010100110;
      patterns[2661] = 29'b0_000101001100_101_0_000001010011;
      patterns[2662] = 29'b0_000101001100_110_0_000101001100;
      patterns[2663] = 29'b0_000101001100_111_0_000101001100;
      patterns[2664] = 29'b0_000101001101_000_0_000101001101;
      patterns[2665] = 29'b0_000101001101_001_0_001101000101;
      patterns[2666] = 29'b0_000101001101_010_0_001010011010;
      patterns[2667] = 29'b0_000101001101_011_0_010100110100;
      patterns[2668] = 29'b0_000101001101_100_1_000010100110;
      patterns[2669] = 29'b0_000101001101_101_0_100001010011;
      patterns[2670] = 29'b0_000101001101_110_0_000101001101;
      patterns[2671] = 29'b0_000101001101_111_0_000101001101;
      patterns[2672] = 29'b0_000101001110_000_0_000101001110;
      patterns[2673] = 29'b0_000101001110_001_0_001110000101;
      patterns[2674] = 29'b0_000101001110_010_0_001010011100;
      patterns[2675] = 29'b0_000101001110_011_0_010100111000;
      patterns[2676] = 29'b0_000101001110_100_0_000010100111;
      patterns[2677] = 29'b0_000101001110_101_1_000001010011;
      patterns[2678] = 29'b0_000101001110_110_0_000101001110;
      patterns[2679] = 29'b0_000101001110_111_0_000101001110;
      patterns[2680] = 29'b0_000101001111_000_0_000101001111;
      patterns[2681] = 29'b0_000101001111_001_0_001111000101;
      patterns[2682] = 29'b0_000101001111_010_0_001010011110;
      patterns[2683] = 29'b0_000101001111_011_0_010100111100;
      patterns[2684] = 29'b0_000101001111_100_1_000010100111;
      patterns[2685] = 29'b0_000101001111_101_1_100001010011;
      patterns[2686] = 29'b0_000101001111_110_0_000101001111;
      patterns[2687] = 29'b0_000101001111_111_0_000101001111;
      patterns[2688] = 29'b0_000101010000_000_0_000101010000;
      patterns[2689] = 29'b0_000101010000_001_0_010000000101;
      patterns[2690] = 29'b0_000101010000_010_0_001010100000;
      patterns[2691] = 29'b0_000101010000_011_0_010101000000;
      patterns[2692] = 29'b0_000101010000_100_0_000010101000;
      patterns[2693] = 29'b0_000101010000_101_0_000001010100;
      patterns[2694] = 29'b0_000101010000_110_0_000101010000;
      patterns[2695] = 29'b0_000101010000_111_0_000101010000;
      patterns[2696] = 29'b0_000101010001_000_0_000101010001;
      patterns[2697] = 29'b0_000101010001_001_0_010001000101;
      patterns[2698] = 29'b0_000101010001_010_0_001010100010;
      patterns[2699] = 29'b0_000101010001_011_0_010101000100;
      patterns[2700] = 29'b0_000101010001_100_1_000010101000;
      patterns[2701] = 29'b0_000101010001_101_0_100001010100;
      patterns[2702] = 29'b0_000101010001_110_0_000101010001;
      patterns[2703] = 29'b0_000101010001_111_0_000101010001;
      patterns[2704] = 29'b0_000101010010_000_0_000101010010;
      patterns[2705] = 29'b0_000101010010_001_0_010010000101;
      patterns[2706] = 29'b0_000101010010_010_0_001010100100;
      patterns[2707] = 29'b0_000101010010_011_0_010101001000;
      patterns[2708] = 29'b0_000101010010_100_0_000010101001;
      patterns[2709] = 29'b0_000101010010_101_1_000001010100;
      patterns[2710] = 29'b0_000101010010_110_0_000101010010;
      patterns[2711] = 29'b0_000101010010_111_0_000101010010;
      patterns[2712] = 29'b0_000101010011_000_0_000101010011;
      patterns[2713] = 29'b0_000101010011_001_0_010011000101;
      patterns[2714] = 29'b0_000101010011_010_0_001010100110;
      patterns[2715] = 29'b0_000101010011_011_0_010101001100;
      patterns[2716] = 29'b0_000101010011_100_1_000010101001;
      patterns[2717] = 29'b0_000101010011_101_1_100001010100;
      patterns[2718] = 29'b0_000101010011_110_0_000101010011;
      patterns[2719] = 29'b0_000101010011_111_0_000101010011;
      patterns[2720] = 29'b0_000101010100_000_0_000101010100;
      patterns[2721] = 29'b0_000101010100_001_0_010100000101;
      patterns[2722] = 29'b0_000101010100_010_0_001010101000;
      patterns[2723] = 29'b0_000101010100_011_0_010101010000;
      patterns[2724] = 29'b0_000101010100_100_0_000010101010;
      patterns[2725] = 29'b0_000101010100_101_0_000001010101;
      patterns[2726] = 29'b0_000101010100_110_0_000101010100;
      patterns[2727] = 29'b0_000101010100_111_0_000101010100;
      patterns[2728] = 29'b0_000101010101_000_0_000101010101;
      patterns[2729] = 29'b0_000101010101_001_0_010101000101;
      patterns[2730] = 29'b0_000101010101_010_0_001010101010;
      patterns[2731] = 29'b0_000101010101_011_0_010101010100;
      patterns[2732] = 29'b0_000101010101_100_1_000010101010;
      patterns[2733] = 29'b0_000101010101_101_0_100001010101;
      patterns[2734] = 29'b0_000101010101_110_0_000101010101;
      patterns[2735] = 29'b0_000101010101_111_0_000101010101;
      patterns[2736] = 29'b0_000101010110_000_0_000101010110;
      patterns[2737] = 29'b0_000101010110_001_0_010110000101;
      patterns[2738] = 29'b0_000101010110_010_0_001010101100;
      patterns[2739] = 29'b0_000101010110_011_0_010101011000;
      patterns[2740] = 29'b0_000101010110_100_0_000010101011;
      patterns[2741] = 29'b0_000101010110_101_1_000001010101;
      patterns[2742] = 29'b0_000101010110_110_0_000101010110;
      patterns[2743] = 29'b0_000101010110_111_0_000101010110;
      patterns[2744] = 29'b0_000101010111_000_0_000101010111;
      patterns[2745] = 29'b0_000101010111_001_0_010111000101;
      patterns[2746] = 29'b0_000101010111_010_0_001010101110;
      patterns[2747] = 29'b0_000101010111_011_0_010101011100;
      patterns[2748] = 29'b0_000101010111_100_1_000010101011;
      patterns[2749] = 29'b0_000101010111_101_1_100001010101;
      patterns[2750] = 29'b0_000101010111_110_0_000101010111;
      patterns[2751] = 29'b0_000101010111_111_0_000101010111;
      patterns[2752] = 29'b0_000101011000_000_0_000101011000;
      patterns[2753] = 29'b0_000101011000_001_0_011000000101;
      patterns[2754] = 29'b0_000101011000_010_0_001010110000;
      patterns[2755] = 29'b0_000101011000_011_0_010101100000;
      patterns[2756] = 29'b0_000101011000_100_0_000010101100;
      patterns[2757] = 29'b0_000101011000_101_0_000001010110;
      patterns[2758] = 29'b0_000101011000_110_0_000101011000;
      patterns[2759] = 29'b0_000101011000_111_0_000101011000;
      patterns[2760] = 29'b0_000101011001_000_0_000101011001;
      patterns[2761] = 29'b0_000101011001_001_0_011001000101;
      patterns[2762] = 29'b0_000101011001_010_0_001010110010;
      patterns[2763] = 29'b0_000101011001_011_0_010101100100;
      patterns[2764] = 29'b0_000101011001_100_1_000010101100;
      patterns[2765] = 29'b0_000101011001_101_0_100001010110;
      patterns[2766] = 29'b0_000101011001_110_0_000101011001;
      patterns[2767] = 29'b0_000101011001_111_0_000101011001;
      patterns[2768] = 29'b0_000101011010_000_0_000101011010;
      patterns[2769] = 29'b0_000101011010_001_0_011010000101;
      patterns[2770] = 29'b0_000101011010_010_0_001010110100;
      patterns[2771] = 29'b0_000101011010_011_0_010101101000;
      patterns[2772] = 29'b0_000101011010_100_0_000010101101;
      patterns[2773] = 29'b0_000101011010_101_1_000001010110;
      patterns[2774] = 29'b0_000101011010_110_0_000101011010;
      patterns[2775] = 29'b0_000101011010_111_0_000101011010;
      patterns[2776] = 29'b0_000101011011_000_0_000101011011;
      patterns[2777] = 29'b0_000101011011_001_0_011011000101;
      patterns[2778] = 29'b0_000101011011_010_0_001010110110;
      patterns[2779] = 29'b0_000101011011_011_0_010101101100;
      patterns[2780] = 29'b0_000101011011_100_1_000010101101;
      patterns[2781] = 29'b0_000101011011_101_1_100001010110;
      patterns[2782] = 29'b0_000101011011_110_0_000101011011;
      patterns[2783] = 29'b0_000101011011_111_0_000101011011;
      patterns[2784] = 29'b0_000101011100_000_0_000101011100;
      patterns[2785] = 29'b0_000101011100_001_0_011100000101;
      patterns[2786] = 29'b0_000101011100_010_0_001010111000;
      patterns[2787] = 29'b0_000101011100_011_0_010101110000;
      patterns[2788] = 29'b0_000101011100_100_0_000010101110;
      patterns[2789] = 29'b0_000101011100_101_0_000001010111;
      patterns[2790] = 29'b0_000101011100_110_0_000101011100;
      patterns[2791] = 29'b0_000101011100_111_0_000101011100;
      patterns[2792] = 29'b0_000101011101_000_0_000101011101;
      patterns[2793] = 29'b0_000101011101_001_0_011101000101;
      patterns[2794] = 29'b0_000101011101_010_0_001010111010;
      patterns[2795] = 29'b0_000101011101_011_0_010101110100;
      patterns[2796] = 29'b0_000101011101_100_1_000010101110;
      patterns[2797] = 29'b0_000101011101_101_0_100001010111;
      patterns[2798] = 29'b0_000101011101_110_0_000101011101;
      patterns[2799] = 29'b0_000101011101_111_0_000101011101;
      patterns[2800] = 29'b0_000101011110_000_0_000101011110;
      patterns[2801] = 29'b0_000101011110_001_0_011110000101;
      patterns[2802] = 29'b0_000101011110_010_0_001010111100;
      patterns[2803] = 29'b0_000101011110_011_0_010101111000;
      patterns[2804] = 29'b0_000101011110_100_0_000010101111;
      patterns[2805] = 29'b0_000101011110_101_1_000001010111;
      patterns[2806] = 29'b0_000101011110_110_0_000101011110;
      patterns[2807] = 29'b0_000101011110_111_0_000101011110;
      patterns[2808] = 29'b0_000101011111_000_0_000101011111;
      patterns[2809] = 29'b0_000101011111_001_0_011111000101;
      patterns[2810] = 29'b0_000101011111_010_0_001010111110;
      patterns[2811] = 29'b0_000101011111_011_0_010101111100;
      patterns[2812] = 29'b0_000101011111_100_1_000010101111;
      patterns[2813] = 29'b0_000101011111_101_1_100001010111;
      patterns[2814] = 29'b0_000101011111_110_0_000101011111;
      patterns[2815] = 29'b0_000101011111_111_0_000101011111;
      patterns[2816] = 29'b0_000101100000_000_0_000101100000;
      patterns[2817] = 29'b0_000101100000_001_0_100000000101;
      patterns[2818] = 29'b0_000101100000_010_0_001011000000;
      patterns[2819] = 29'b0_000101100000_011_0_010110000000;
      patterns[2820] = 29'b0_000101100000_100_0_000010110000;
      patterns[2821] = 29'b0_000101100000_101_0_000001011000;
      patterns[2822] = 29'b0_000101100000_110_0_000101100000;
      patterns[2823] = 29'b0_000101100000_111_0_000101100000;
      patterns[2824] = 29'b0_000101100001_000_0_000101100001;
      patterns[2825] = 29'b0_000101100001_001_0_100001000101;
      patterns[2826] = 29'b0_000101100001_010_0_001011000010;
      patterns[2827] = 29'b0_000101100001_011_0_010110000100;
      patterns[2828] = 29'b0_000101100001_100_1_000010110000;
      patterns[2829] = 29'b0_000101100001_101_0_100001011000;
      patterns[2830] = 29'b0_000101100001_110_0_000101100001;
      patterns[2831] = 29'b0_000101100001_111_0_000101100001;
      patterns[2832] = 29'b0_000101100010_000_0_000101100010;
      patterns[2833] = 29'b0_000101100010_001_0_100010000101;
      patterns[2834] = 29'b0_000101100010_010_0_001011000100;
      patterns[2835] = 29'b0_000101100010_011_0_010110001000;
      patterns[2836] = 29'b0_000101100010_100_0_000010110001;
      patterns[2837] = 29'b0_000101100010_101_1_000001011000;
      patterns[2838] = 29'b0_000101100010_110_0_000101100010;
      patterns[2839] = 29'b0_000101100010_111_0_000101100010;
      patterns[2840] = 29'b0_000101100011_000_0_000101100011;
      patterns[2841] = 29'b0_000101100011_001_0_100011000101;
      patterns[2842] = 29'b0_000101100011_010_0_001011000110;
      patterns[2843] = 29'b0_000101100011_011_0_010110001100;
      patterns[2844] = 29'b0_000101100011_100_1_000010110001;
      patterns[2845] = 29'b0_000101100011_101_1_100001011000;
      patterns[2846] = 29'b0_000101100011_110_0_000101100011;
      patterns[2847] = 29'b0_000101100011_111_0_000101100011;
      patterns[2848] = 29'b0_000101100100_000_0_000101100100;
      patterns[2849] = 29'b0_000101100100_001_0_100100000101;
      patterns[2850] = 29'b0_000101100100_010_0_001011001000;
      patterns[2851] = 29'b0_000101100100_011_0_010110010000;
      patterns[2852] = 29'b0_000101100100_100_0_000010110010;
      patterns[2853] = 29'b0_000101100100_101_0_000001011001;
      patterns[2854] = 29'b0_000101100100_110_0_000101100100;
      patterns[2855] = 29'b0_000101100100_111_0_000101100100;
      patterns[2856] = 29'b0_000101100101_000_0_000101100101;
      patterns[2857] = 29'b0_000101100101_001_0_100101000101;
      patterns[2858] = 29'b0_000101100101_010_0_001011001010;
      patterns[2859] = 29'b0_000101100101_011_0_010110010100;
      patterns[2860] = 29'b0_000101100101_100_1_000010110010;
      patterns[2861] = 29'b0_000101100101_101_0_100001011001;
      patterns[2862] = 29'b0_000101100101_110_0_000101100101;
      patterns[2863] = 29'b0_000101100101_111_0_000101100101;
      patterns[2864] = 29'b0_000101100110_000_0_000101100110;
      patterns[2865] = 29'b0_000101100110_001_0_100110000101;
      patterns[2866] = 29'b0_000101100110_010_0_001011001100;
      patterns[2867] = 29'b0_000101100110_011_0_010110011000;
      patterns[2868] = 29'b0_000101100110_100_0_000010110011;
      patterns[2869] = 29'b0_000101100110_101_1_000001011001;
      patterns[2870] = 29'b0_000101100110_110_0_000101100110;
      patterns[2871] = 29'b0_000101100110_111_0_000101100110;
      patterns[2872] = 29'b0_000101100111_000_0_000101100111;
      patterns[2873] = 29'b0_000101100111_001_0_100111000101;
      patterns[2874] = 29'b0_000101100111_010_0_001011001110;
      patterns[2875] = 29'b0_000101100111_011_0_010110011100;
      patterns[2876] = 29'b0_000101100111_100_1_000010110011;
      patterns[2877] = 29'b0_000101100111_101_1_100001011001;
      patterns[2878] = 29'b0_000101100111_110_0_000101100111;
      patterns[2879] = 29'b0_000101100111_111_0_000101100111;
      patterns[2880] = 29'b0_000101101000_000_0_000101101000;
      patterns[2881] = 29'b0_000101101000_001_0_101000000101;
      patterns[2882] = 29'b0_000101101000_010_0_001011010000;
      patterns[2883] = 29'b0_000101101000_011_0_010110100000;
      patterns[2884] = 29'b0_000101101000_100_0_000010110100;
      patterns[2885] = 29'b0_000101101000_101_0_000001011010;
      patterns[2886] = 29'b0_000101101000_110_0_000101101000;
      patterns[2887] = 29'b0_000101101000_111_0_000101101000;
      patterns[2888] = 29'b0_000101101001_000_0_000101101001;
      patterns[2889] = 29'b0_000101101001_001_0_101001000101;
      patterns[2890] = 29'b0_000101101001_010_0_001011010010;
      patterns[2891] = 29'b0_000101101001_011_0_010110100100;
      patterns[2892] = 29'b0_000101101001_100_1_000010110100;
      patterns[2893] = 29'b0_000101101001_101_0_100001011010;
      patterns[2894] = 29'b0_000101101001_110_0_000101101001;
      patterns[2895] = 29'b0_000101101001_111_0_000101101001;
      patterns[2896] = 29'b0_000101101010_000_0_000101101010;
      patterns[2897] = 29'b0_000101101010_001_0_101010000101;
      patterns[2898] = 29'b0_000101101010_010_0_001011010100;
      patterns[2899] = 29'b0_000101101010_011_0_010110101000;
      patterns[2900] = 29'b0_000101101010_100_0_000010110101;
      patterns[2901] = 29'b0_000101101010_101_1_000001011010;
      patterns[2902] = 29'b0_000101101010_110_0_000101101010;
      patterns[2903] = 29'b0_000101101010_111_0_000101101010;
      patterns[2904] = 29'b0_000101101011_000_0_000101101011;
      patterns[2905] = 29'b0_000101101011_001_0_101011000101;
      patterns[2906] = 29'b0_000101101011_010_0_001011010110;
      patterns[2907] = 29'b0_000101101011_011_0_010110101100;
      patterns[2908] = 29'b0_000101101011_100_1_000010110101;
      patterns[2909] = 29'b0_000101101011_101_1_100001011010;
      patterns[2910] = 29'b0_000101101011_110_0_000101101011;
      patterns[2911] = 29'b0_000101101011_111_0_000101101011;
      patterns[2912] = 29'b0_000101101100_000_0_000101101100;
      patterns[2913] = 29'b0_000101101100_001_0_101100000101;
      patterns[2914] = 29'b0_000101101100_010_0_001011011000;
      patterns[2915] = 29'b0_000101101100_011_0_010110110000;
      patterns[2916] = 29'b0_000101101100_100_0_000010110110;
      patterns[2917] = 29'b0_000101101100_101_0_000001011011;
      patterns[2918] = 29'b0_000101101100_110_0_000101101100;
      patterns[2919] = 29'b0_000101101100_111_0_000101101100;
      patterns[2920] = 29'b0_000101101101_000_0_000101101101;
      patterns[2921] = 29'b0_000101101101_001_0_101101000101;
      patterns[2922] = 29'b0_000101101101_010_0_001011011010;
      patterns[2923] = 29'b0_000101101101_011_0_010110110100;
      patterns[2924] = 29'b0_000101101101_100_1_000010110110;
      patterns[2925] = 29'b0_000101101101_101_0_100001011011;
      patterns[2926] = 29'b0_000101101101_110_0_000101101101;
      patterns[2927] = 29'b0_000101101101_111_0_000101101101;
      patterns[2928] = 29'b0_000101101110_000_0_000101101110;
      patterns[2929] = 29'b0_000101101110_001_0_101110000101;
      patterns[2930] = 29'b0_000101101110_010_0_001011011100;
      patterns[2931] = 29'b0_000101101110_011_0_010110111000;
      patterns[2932] = 29'b0_000101101110_100_0_000010110111;
      patterns[2933] = 29'b0_000101101110_101_1_000001011011;
      patterns[2934] = 29'b0_000101101110_110_0_000101101110;
      patterns[2935] = 29'b0_000101101110_111_0_000101101110;
      patterns[2936] = 29'b0_000101101111_000_0_000101101111;
      patterns[2937] = 29'b0_000101101111_001_0_101111000101;
      patterns[2938] = 29'b0_000101101111_010_0_001011011110;
      patterns[2939] = 29'b0_000101101111_011_0_010110111100;
      patterns[2940] = 29'b0_000101101111_100_1_000010110111;
      patterns[2941] = 29'b0_000101101111_101_1_100001011011;
      patterns[2942] = 29'b0_000101101111_110_0_000101101111;
      patterns[2943] = 29'b0_000101101111_111_0_000101101111;
      patterns[2944] = 29'b0_000101110000_000_0_000101110000;
      patterns[2945] = 29'b0_000101110000_001_0_110000000101;
      patterns[2946] = 29'b0_000101110000_010_0_001011100000;
      patterns[2947] = 29'b0_000101110000_011_0_010111000000;
      patterns[2948] = 29'b0_000101110000_100_0_000010111000;
      patterns[2949] = 29'b0_000101110000_101_0_000001011100;
      patterns[2950] = 29'b0_000101110000_110_0_000101110000;
      patterns[2951] = 29'b0_000101110000_111_0_000101110000;
      patterns[2952] = 29'b0_000101110001_000_0_000101110001;
      patterns[2953] = 29'b0_000101110001_001_0_110001000101;
      patterns[2954] = 29'b0_000101110001_010_0_001011100010;
      patterns[2955] = 29'b0_000101110001_011_0_010111000100;
      patterns[2956] = 29'b0_000101110001_100_1_000010111000;
      patterns[2957] = 29'b0_000101110001_101_0_100001011100;
      patterns[2958] = 29'b0_000101110001_110_0_000101110001;
      patterns[2959] = 29'b0_000101110001_111_0_000101110001;
      patterns[2960] = 29'b0_000101110010_000_0_000101110010;
      patterns[2961] = 29'b0_000101110010_001_0_110010000101;
      patterns[2962] = 29'b0_000101110010_010_0_001011100100;
      patterns[2963] = 29'b0_000101110010_011_0_010111001000;
      patterns[2964] = 29'b0_000101110010_100_0_000010111001;
      patterns[2965] = 29'b0_000101110010_101_1_000001011100;
      patterns[2966] = 29'b0_000101110010_110_0_000101110010;
      patterns[2967] = 29'b0_000101110010_111_0_000101110010;
      patterns[2968] = 29'b0_000101110011_000_0_000101110011;
      patterns[2969] = 29'b0_000101110011_001_0_110011000101;
      patterns[2970] = 29'b0_000101110011_010_0_001011100110;
      patterns[2971] = 29'b0_000101110011_011_0_010111001100;
      patterns[2972] = 29'b0_000101110011_100_1_000010111001;
      patterns[2973] = 29'b0_000101110011_101_1_100001011100;
      patterns[2974] = 29'b0_000101110011_110_0_000101110011;
      patterns[2975] = 29'b0_000101110011_111_0_000101110011;
      patterns[2976] = 29'b0_000101110100_000_0_000101110100;
      patterns[2977] = 29'b0_000101110100_001_0_110100000101;
      patterns[2978] = 29'b0_000101110100_010_0_001011101000;
      patterns[2979] = 29'b0_000101110100_011_0_010111010000;
      patterns[2980] = 29'b0_000101110100_100_0_000010111010;
      patterns[2981] = 29'b0_000101110100_101_0_000001011101;
      patterns[2982] = 29'b0_000101110100_110_0_000101110100;
      patterns[2983] = 29'b0_000101110100_111_0_000101110100;
      patterns[2984] = 29'b0_000101110101_000_0_000101110101;
      patterns[2985] = 29'b0_000101110101_001_0_110101000101;
      patterns[2986] = 29'b0_000101110101_010_0_001011101010;
      patterns[2987] = 29'b0_000101110101_011_0_010111010100;
      patterns[2988] = 29'b0_000101110101_100_1_000010111010;
      patterns[2989] = 29'b0_000101110101_101_0_100001011101;
      patterns[2990] = 29'b0_000101110101_110_0_000101110101;
      patterns[2991] = 29'b0_000101110101_111_0_000101110101;
      patterns[2992] = 29'b0_000101110110_000_0_000101110110;
      patterns[2993] = 29'b0_000101110110_001_0_110110000101;
      patterns[2994] = 29'b0_000101110110_010_0_001011101100;
      patterns[2995] = 29'b0_000101110110_011_0_010111011000;
      patterns[2996] = 29'b0_000101110110_100_0_000010111011;
      patterns[2997] = 29'b0_000101110110_101_1_000001011101;
      patterns[2998] = 29'b0_000101110110_110_0_000101110110;
      patterns[2999] = 29'b0_000101110110_111_0_000101110110;
      patterns[3000] = 29'b0_000101110111_000_0_000101110111;
      patterns[3001] = 29'b0_000101110111_001_0_110111000101;
      patterns[3002] = 29'b0_000101110111_010_0_001011101110;
      patterns[3003] = 29'b0_000101110111_011_0_010111011100;
      patterns[3004] = 29'b0_000101110111_100_1_000010111011;
      patterns[3005] = 29'b0_000101110111_101_1_100001011101;
      patterns[3006] = 29'b0_000101110111_110_0_000101110111;
      patterns[3007] = 29'b0_000101110111_111_0_000101110111;
      patterns[3008] = 29'b0_000101111000_000_0_000101111000;
      patterns[3009] = 29'b0_000101111000_001_0_111000000101;
      patterns[3010] = 29'b0_000101111000_010_0_001011110000;
      patterns[3011] = 29'b0_000101111000_011_0_010111100000;
      patterns[3012] = 29'b0_000101111000_100_0_000010111100;
      patterns[3013] = 29'b0_000101111000_101_0_000001011110;
      patterns[3014] = 29'b0_000101111000_110_0_000101111000;
      patterns[3015] = 29'b0_000101111000_111_0_000101111000;
      patterns[3016] = 29'b0_000101111001_000_0_000101111001;
      patterns[3017] = 29'b0_000101111001_001_0_111001000101;
      patterns[3018] = 29'b0_000101111001_010_0_001011110010;
      patterns[3019] = 29'b0_000101111001_011_0_010111100100;
      patterns[3020] = 29'b0_000101111001_100_1_000010111100;
      patterns[3021] = 29'b0_000101111001_101_0_100001011110;
      patterns[3022] = 29'b0_000101111001_110_0_000101111001;
      patterns[3023] = 29'b0_000101111001_111_0_000101111001;
      patterns[3024] = 29'b0_000101111010_000_0_000101111010;
      patterns[3025] = 29'b0_000101111010_001_0_111010000101;
      patterns[3026] = 29'b0_000101111010_010_0_001011110100;
      patterns[3027] = 29'b0_000101111010_011_0_010111101000;
      patterns[3028] = 29'b0_000101111010_100_0_000010111101;
      patterns[3029] = 29'b0_000101111010_101_1_000001011110;
      patterns[3030] = 29'b0_000101111010_110_0_000101111010;
      patterns[3031] = 29'b0_000101111010_111_0_000101111010;
      patterns[3032] = 29'b0_000101111011_000_0_000101111011;
      patterns[3033] = 29'b0_000101111011_001_0_111011000101;
      patterns[3034] = 29'b0_000101111011_010_0_001011110110;
      patterns[3035] = 29'b0_000101111011_011_0_010111101100;
      patterns[3036] = 29'b0_000101111011_100_1_000010111101;
      patterns[3037] = 29'b0_000101111011_101_1_100001011110;
      patterns[3038] = 29'b0_000101111011_110_0_000101111011;
      patterns[3039] = 29'b0_000101111011_111_0_000101111011;
      patterns[3040] = 29'b0_000101111100_000_0_000101111100;
      patterns[3041] = 29'b0_000101111100_001_0_111100000101;
      patterns[3042] = 29'b0_000101111100_010_0_001011111000;
      patterns[3043] = 29'b0_000101111100_011_0_010111110000;
      patterns[3044] = 29'b0_000101111100_100_0_000010111110;
      patterns[3045] = 29'b0_000101111100_101_0_000001011111;
      patterns[3046] = 29'b0_000101111100_110_0_000101111100;
      patterns[3047] = 29'b0_000101111100_111_0_000101111100;
      patterns[3048] = 29'b0_000101111101_000_0_000101111101;
      patterns[3049] = 29'b0_000101111101_001_0_111101000101;
      patterns[3050] = 29'b0_000101111101_010_0_001011111010;
      patterns[3051] = 29'b0_000101111101_011_0_010111110100;
      patterns[3052] = 29'b0_000101111101_100_1_000010111110;
      patterns[3053] = 29'b0_000101111101_101_0_100001011111;
      patterns[3054] = 29'b0_000101111101_110_0_000101111101;
      patterns[3055] = 29'b0_000101111101_111_0_000101111101;
      patterns[3056] = 29'b0_000101111110_000_0_000101111110;
      patterns[3057] = 29'b0_000101111110_001_0_111110000101;
      patterns[3058] = 29'b0_000101111110_010_0_001011111100;
      patterns[3059] = 29'b0_000101111110_011_0_010111111000;
      patterns[3060] = 29'b0_000101111110_100_0_000010111111;
      patterns[3061] = 29'b0_000101111110_101_1_000001011111;
      patterns[3062] = 29'b0_000101111110_110_0_000101111110;
      patterns[3063] = 29'b0_000101111110_111_0_000101111110;
      patterns[3064] = 29'b0_000101111111_000_0_000101111111;
      patterns[3065] = 29'b0_000101111111_001_0_111111000101;
      patterns[3066] = 29'b0_000101111111_010_0_001011111110;
      patterns[3067] = 29'b0_000101111111_011_0_010111111100;
      patterns[3068] = 29'b0_000101111111_100_1_000010111111;
      patterns[3069] = 29'b0_000101111111_101_1_100001011111;
      patterns[3070] = 29'b0_000101111111_110_0_000101111111;
      patterns[3071] = 29'b0_000101111111_111_0_000101111111;
      patterns[3072] = 29'b0_000110000000_000_0_000110000000;
      patterns[3073] = 29'b0_000110000000_001_0_000000000110;
      patterns[3074] = 29'b0_000110000000_010_0_001100000000;
      patterns[3075] = 29'b0_000110000000_011_0_011000000000;
      patterns[3076] = 29'b0_000110000000_100_0_000011000000;
      patterns[3077] = 29'b0_000110000000_101_0_000001100000;
      patterns[3078] = 29'b0_000110000000_110_0_000110000000;
      patterns[3079] = 29'b0_000110000000_111_0_000110000000;
      patterns[3080] = 29'b0_000110000001_000_0_000110000001;
      patterns[3081] = 29'b0_000110000001_001_0_000001000110;
      patterns[3082] = 29'b0_000110000001_010_0_001100000010;
      patterns[3083] = 29'b0_000110000001_011_0_011000000100;
      patterns[3084] = 29'b0_000110000001_100_1_000011000000;
      patterns[3085] = 29'b0_000110000001_101_0_100001100000;
      patterns[3086] = 29'b0_000110000001_110_0_000110000001;
      patterns[3087] = 29'b0_000110000001_111_0_000110000001;
      patterns[3088] = 29'b0_000110000010_000_0_000110000010;
      patterns[3089] = 29'b0_000110000010_001_0_000010000110;
      patterns[3090] = 29'b0_000110000010_010_0_001100000100;
      patterns[3091] = 29'b0_000110000010_011_0_011000001000;
      patterns[3092] = 29'b0_000110000010_100_0_000011000001;
      patterns[3093] = 29'b0_000110000010_101_1_000001100000;
      patterns[3094] = 29'b0_000110000010_110_0_000110000010;
      patterns[3095] = 29'b0_000110000010_111_0_000110000010;
      patterns[3096] = 29'b0_000110000011_000_0_000110000011;
      patterns[3097] = 29'b0_000110000011_001_0_000011000110;
      patterns[3098] = 29'b0_000110000011_010_0_001100000110;
      patterns[3099] = 29'b0_000110000011_011_0_011000001100;
      patterns[3100] = 29'b0_000110000011_100_1_000011000001;
      patterns[3101] = 29'b0_000110000011_101_1_100001100000;
      patterns[3102] = 29'b0_000110000011_110_0_000110000011;
      patterns[3103] = 29'b0_000110000011_111_0_000110000011;
      patterns[3104] = 29'b0_000110000100_000_0_000110000100;
      patterns[3105] = 29'b0_000110000100_001_0_000100000110;
      patterns[3106] = 29'b0_000110000100_010_0_001100001000;
      patterns[3107] = 29'b0_000110000100_011_0_011000010000;
      patterns[3108] = 29'b0_000110000100_100_0_000011000010;
      patterns[3109] = 29'b0_000110000100_101_0_000001100001;
      patterns[3110] = 29'b0_000110000100_110_0_000110000100;
      patterns[3111] = 29'b0_000110000100_111_0_000110000100;
      patterns[3112] = 29'b0_000110000101_000_0_000110000101;
      patterns[3113] = 29'b0_000110000101_001_0_000101000110;
      patterns[3114] = 29'b0_000110000101_010_0_001100001010;
      patterns[3115] = 29'b0_000110000101_011_0_011000010100;
      patterns[3116] = 29'b0_000110000101_100_1_000011000010;
      patterns[3117] = 29'b0_000110000101_101_0_100001100001;
      patterns[3118] = 29'b0_000110000101_110_0_000110000101;
      patterns[3119] = 29'b0_000110000101_111_0_000110000101;
      patterns[3120] = 29'b0_000110000110_000_0_000110000110;
      patterns[3121] = 29'b0_000110000110_001_0_000110000110;
      patterns[3122] = 29'b0_000110000110_010_0_001100001100;
      patterns[3123] = 29'b0_000110000110_011_0_011000011000;
      patterns[3124] = 29'b0_000110000110_100_0_000011000011;
      patterns[3125] = 29'b0_000110000110_101_1_000001100001;
      patterns[3126] = 29'b0_000110000110_110_0_000110000110;
      patterns[3127] = 29'b0_000110000110_111_0_000110000110;
      patterns[3128] = 29'b0_000110000111_000_0_000110000111;
      patterns[3129] = 29'b0_000110000111_001_0_000111000110;
      patterns[3130] = 29'b0_000110000111_010_0_001100001110;
      patterns[3131] = 29'b0_000110000111_011_0_011000011100;
      patterns[3132] = 29'b0_000110000111_100_1_000011000011;
      patterns[3133] = 29'b0_000110000111_101_1_100001100001;
      patterns[3134] = 29'b0_000110000111_110_0_000110000111;
      patterns[3135] = 29'b0_000110000111_111_0_000110000111;
      patterns[3136] = 29'b0_000110001000_000_0_000110001000;
      patterns[3137] = 29'b0_000110001000_001_0_001000000110;
      patterns[3138] = 29'b0_000110001000_010_0_001100010000;
      patterns[3139] = 29'b0_000110001000_011_0_011000100000;
      patterns[3140] = 29'b0_000110001000_100_0_000011000100;
      patterns[3141] = 29'b0_000110001000_101_0_000001100010;
      patterns[3142] = 29'b0_000110001000_110_0_000110001000;
      patterns[3143] = 29'b0_000110001000_111_0_000110001000;
      patterns[3144] = 29'b0_000110001001_000_0_000110001001;
      patterns[3145] = 29'b0_000110001001_001_0_001001000110;
      patterns[3146] = 29'b0_000110001001_010_0_001100010010;
      patterns[3147] = 29'b0_000110001001_011_0_011000100100;
      patterns[3148] = 29'b0_000110001001_100_1_000011000100;
      patterns[3149] = 29'b0_000110001001_101_0_100001100010;
      patterns[3150] = 29'b0_000110001001_110_0_000110001001;
      patterns[3151] = 29'b0_000110001001_111_0_000110001001;
      patterns[3152] = 29'b0_000110001010_000_0_000110001010;
      patterns[3153] = 29'b0_000110001010_001_0_001010000110;
      patterns[3154] = 29'b0_000110001010_010_0_001100010100;
      patterns[3155] = 29'b0_000110001010_011_0_011000101000;
      patterns[3156] = 29'b0_000110001010_100_0_000011000101;
      patterns[3157] = 29'b0_000110001010_101_1_000001100010;
      patterns[3158] = 29'b0_000110001010_110_0_000110001010;
      patterns[3159] = 29'b0_000110001010_111_0_000110001010;
      patterns[3160] = 29'b0_000110001011_000_0_000110001011;
      patterns[3161] = 29'b0_000110001011_001_0_001011000110;
      patterns[3162] = 29'b0_000110001011_010_0_001100010110;
      patterns[3163] = 29'b0_000110001011_011_0_011000101100;
      patterns[3164] = 29'b0_000110001011_100_1_000011000101;
      patterns[3165] = 29'b0_000110001011_101_1_100001100010;
      patterns[3166] = 29'b0_000110001011_110_0_000110001011;
      patterns[3167] = 29'b0_000110001011_111_0_000110001011;
      patterns[3168] = 29'b0_000110001100_000_0_000110001100;
      patterns[3169] = 29'b0_000110001100_001_0_001100000110;
      patterns[3170] = 29'b0_000110001100_010_0_001100011000;
      patterns[3171] = 29'b0_000110001100_011_0_011000110000;
      patterns[3172] = 29'b0_000110001100_100_0_000011000110;
      patterns[3173] = 29'b0_000110001100_101_0_000001100011;
      patterns[3174] = 29'b0_000110001100_110_0_000110001100;
      patterns[3175] = 29'b0_000110001100_111_0_000110001100;
      patterns[3176] = 29'b0_000110001101_000_0_000110001101;
      patterns[3177] = 29'b0_000110001101_001_0_001101000110;
      patterns[3178] = 29'b0_000110001101_010_0_001100011010;
      patterns[3179] = 29'b0_000110001101_011_0_011000110100;
      patterns[3180] = 29'b0_000110001101_100_1_000011000110;
      patterns[3181] = 29'b0_000110001101_101_0_100001100011;
      patterns[3182] = 29'b0_000110001101_110_0_000110001101;
      patterns[3183] = 29'b0_000110001101_111_0_000110001101;
      patterns[3184] = 29'b0_000110001110_000_0_000110001110;
      patterns[3185] = 29'b0_000110001110_001_0_001110000110;
      patterns[3186] = 29'b0_000110001110_010_0_001100011100;
      patterns[3187] = 29'b0_000110001110_011_0_011000111000;
      patterns[3188] = 29'b0_000110001110_100_0_000011000111;
      patterns[3189] = 29'b0_000110001110_101_1_000001100011;
      patterns[3190] = 29'b0_000110001110_110_0_000110001110;
      patterns[3191] = 29'b0_000110001110_111_0_000110001110;
      patterns[3192] = 29'b0_000110001111_000_0_000110001111;
      patterns[3193] = 29'b0_000110001111_001_0_001111000110;
      patterns[3194] = 29'b0_000110001111_010_0_001100011110;
      patterns[3195] = 29'b0_000110001111_011_0_011000111100;
      patterns[3196] = 29'b0_000110001111_100_1_000011000111;
      patterns[3197] = 29'b0_000110001111_101_1_100001100011;
      patterns[3198] = 29'b0_000110001111_110_0_000110001111;
      patterns[3199] = 29'b0_000110001111_111_0_000110001111;
      patterns[3200] = 29'b0_000110010000_000_0_000110010000;
      patterns[3201] = 29'b0_000110010000_001_0_010000000110;
      patterns[3202] = 29'b0_000110010000_010_0_001100100000;
      patterns[3203] = 29'b0_000110010000_011_0_011001000000;
      patterns[3204] = 29'b0_000110010000_100_0_000011001000;
      patterns[3205] = 29'b0_000110010000_101_0_000001100100;
      patterns[3206] = 29'b0_000110010000_110_0_000110010000;
      patterns[3207] = 29'b0_000110010000_111_0_000110010000;
      patterns[3208] = 29'b0_000110010001_000_0_000110010001;
      patterns[3209] = 29'b0_000110010001_001_0_010001000110;
      patterns[3210] = 29'b0_000110010001_010_0_001100100010;
      patterns[3211] = 29'b0_000110010001_011_0_011001000100;
      patterns[3212] = 29'b0_000110010001_100_1_000011001000;
      patterns[3213] = 29'b0_000110010001_101_0_100001100100;
      patterns[3214] = 29'b0_000110010001_110_0_000110010001;
      patterns[3215] = 29'b0_000110010001_111_0_000110010001;
      patterns[3216] = 29'b0_000110010010_000_0_000110010010;
      patterns[3217] = 29'b0_000110010010_001_0_010010000110;
      patterns[3218] = 29'b0_000110010010_010_0_001100100100;
      patterns[3219] = 29'b0_000110010010_011_0_011001001000;
      patterns[3220] = 29'b0_000110010010_100_0_000011001001;
      patterns[3221] = 29'b0_000110010010_101_1_000001100100;
      patterns[3222] = 29'b0_000110010010_110_0_000110010010;
      patterns[3223] = 29'b0_000110010010_111_0_000110010010;
      patterns[3224] = 29'b0_000110010011_000_0_000110010011;
      patterns[3225] = 29'b0_000110010011_001_0_010011000110;
      patterns[3226] = 29'b0_000110010011_010_0_001100100110;
      patterns[3227] = 29'b0_000110010011_011_0_011001001100;
      patterns[3228] = 29'b0_000110010011_100_1_000011001001;
      patterns[3229] = 29'b0_000110010011_101_1_100001100100;
      patterns[3230] = 29'b0_000110010011_110_0_000110010011;
      patterns[3231] = 29'b0_000110010011_111_0_000110010011;
      patterns[3232] = 29'b0_000110010100_000_0_000110010100;
      patterns[3233] = 29'b0_000110010100_001_0_010100000110;
      patterns[3234] = 29'b0_000110010100_010_0_001100101000;
      patterns[3235] = 29'b0_000110010100_011_0_011001010000;
      patterns[3236] = 29'b0_000110010100_100_0_000011001010;
      patterns[3237] = 29'b0_000110010100_101_0_000001100101;
      patterns[3238] = 29'b0_000110010100_110_0_000110010100;
      patterns[3239] = 29'b0_000110010100_111_0_000110010100;
      patterns[3240] = 29'b0_000110010101_000_0_000110010101;
      patterns[3241] = 29'b0_000110010101_001_0_010101000110;
      patterns[3242] = 29'b0_000110010101_010_0_001100101010;
      patterns[3243] = 29'b0_000110010101_011_0_011001010100;
      patterns[3244] = 29'b0_000110010101_100_1_000011001010;
      patterns[3245] = 29'b0_000110010101_101_0_100001100101;
      patterns[3246] = 29'b0_000110010101_110_0_000110010101;
      patterns[3247] = 29'b0_000110010101_111_0_000110010101;
      patterns[3248] = 29'b0_000110010110_000_0_000110010110;
      patterns[3249] = 29'b0_000110010110_001_0_010110000110;
      patterns[3250] = 29'b0_000110010110_010_0_001100101100;
      patterns[3251] = 29'b0_000110010110_011_0_011001011000;
      patterns[3252] = 29'b0_000110010110_100_0_000011001011;
      patterns[3253] = 29'b0_000110010110_101_1_000001100101;
      patterns[3254] = 29'b0_000110010110_110_0_000110010110;
      patterns[3255] = 29'b0_000110010110_111_0_000110010110;
      patterns[3256] = 29'b0_000110010111_000_0_000110010111;
      patterns[3257] = 29'b0_000110010111_001_0_010111000110;
      patterns[3258] = 29'b0_000110010111_010_0_001100101110;
      patterns[3259] = 29'b0_000110010111_011_0_011001011100;
      patterns[3260] = 29'b0_000110010111_100_1_000011001011;
      patterns[3261] = 29'b0_000110010111_101_1_100001100101;
      patterns[3262] = 29'b0_000110010111_110_0_000110010111;
      patterns[3263] = 29'b0_000110010111_111_0_000110010111;
      patterns[3264] = 29'b0_000110011000_000_0_000110011000;
      patterns[3265] = 29'b0_000110011000_001_0_011000000110;
      patterns[3266] = 29'b0_000110011000_010_0_001100110000;
      patterns[3267] = 29'b0_000110011000_011_0_011001100000;
      patterns[3268] = 29'b0_000110011000_100_0_000011001100;
      patterns[3269] = 29'b0_000110011000_101_0_000001100110;
      patterns[3270] = 29'b0_000110011000_110_0_000110011000;
      patterns[3271] = 29'b0_000110011000_111_0_000110011000;
      patterns[3272] = 29'b0_000110011001_000_0_000110011001;
      patterns[3273] = 29'b0_000110011001_001_0_011001000110;
      patterns[3274] = 29'b0_000110011001_010_0_001100110010;
      patterns[3275] = 29'b0_000110011001_011_0_011001100100;
      patterns[3276] = 29'b0_000110011001_100_1_000011001100;
      patterns[3277] = 29'b0_000110011001_101_0_100001100110;
      patterns[3278] = 29'b0_000110011001_110_0_000110011001;
      patterns[3279] = 29'b0_000110011001_111_0_000110011001;
      patterns[3280] = 29'b0_000110011010_000_0_000110011010;
      patterns[3281] = 29'b0_000110011010_001_0_011010000110;
      patterns[3282] = 29'b0_000110011010_010_0_001100110100;
      patterns[3283] = 29'b0_000110011010_011_0_011001101000;
      patterns[3284] = 29'b0_000110011010_100_0_000011001101;
      patterns[3285] = 29'b0_000110011010_101_1_000001100110;
      patterns[3286] = 29'b0_000110011010_110_0_000110011010;
      patterns[3287] = 29'b0_000110011010_111_0_000110011010;
      patterns[3288] = 29'b0_000110011011_000_0_000110011011;
      patterns[3289] = 29'b0_000110011011_001_0_011011000110;
      patterns[3290] = 29'b0_000110011011_010_0_001100110110;
      patterns[3291] = 29'b0_000110011011_011_0_011001101100;
      patterns[3292] = 29'b0_000110011011_100_1_000011001101;
      patterns[3293] = 29'b0_000110011011_101_1_100001100110;
      patterns[3294] = 29'b0_000110011011_110_0_000110011011;
      patterns[3295] = 29'b0_000110011011_111_0_000110011011;
      patterns[3296] = 29'b0_000110011100_000_0_000110011100;
      patterns[3297] = 29'b0_000110011100_001_0_011100000110;
      patterns[3298] = 29'b0_000110011100_010_0_001100111000;
      patterns[3299] = 29'b0_000110011100_011_0_011001110000;
      patterns[3300] = 29'b0_000110011100_100_0_000011001110;
      patterns[3301] = 29'b0_000110011100_101_0_000001100111;
      patterns[3302] = 29'b0_000110011100_110_0_000110011100;
      patterns[3303] = 29'b0_000110011100_111_0_000110011100;
      patterns[3304] = 29'b0_000110011101_000_0_000110011101;
      patterns[3305] = 29'b0_000110011101_001_0_011101000110;
      patterns[3306] = 29'b0_000110011101_010_0_001100111010;
      patterns[3307] = 29'b0_000110011101_011_0_011001110100;
      patterns[3308] = 29'b0_000110011101_100_1_000011001110;
      patterns[3309] = 29'b0_000110011101_101_0_100001100111;
      patterns[3310] = 29'b0_000110011101_110_0_000110011101;
      patterns[3311] = 29'b0_000110011101_111_0_000110011101;
      patterns[3312] = 29'b0_000110011110_000_0_000110011110;
      patterns[3313] = 29'b0_000110011110_001_0_011110000110;
      patterns[3314] = 29'b0_000110011110_010_0_001100111100;
      patterns[3315] = 29'b0_000110011110_011_0_011001111000;
      patterns[3316] = 29'b0_000110011110_100_0_000011001111;
      patterns[3317] = 29'b0_000110011110_101_1_000001100111;
      patterns[3318] = 29'b0_000110011110_110_0_000110011110;
      patterns[3319] = 29'b0_000110011110_111_0_000110011110;
      patterns[3320] = 29'b0_000110011111_000_0_000110011111;
      patterns[3321] = 29'b0_000110011111_001_0_011111000110;
      patterns[3322] = 29'b0_000110011111_010_0_001100111110;
      patterns[3323] = 29'b0_000110011111_011_0_011001111100;
      patterns[3324] = 29'b0_000110011111_100_1_000011001111;
      patterns[3325] = 29'b0_000110011111_101_1_100001100111;
      patterns[3326] = 29'b0_000110011111_110_0_000110011111;
      patterns[3327] = 29'b0_000110011111_111_0_000110011111;
      patterns[3328] = 29'b0_000110100000_000_0_000110100000;
      patterns[3329] = 29'b0_000110100000_001_0_100000000110;
      patterns[3330] = 29'b0_000110100000_010_0_001101000000;
      patterns[3331] = 29'b0_000110100000_011_0_011010000000;
      patterns[3332] = 29'b0_000110100000_100_0_000011010000;
      patterns[3333] = 29'b0_000110100000_101_0_000001101000;
      patterns[3334] = 29'b0_000110100000_110_0_000110100000;
      patterns[3335] = 29'b0_000110100000_111_0_000110100000;
      patterns[3336] = 29'b0_000110100001_000_0_000110100001;
      patterns[3337] = 29'b0_000110100001_001_0_100001000110;
      patterns[3338] = 29'b0_000110100001_010_0_001101000010;
      patterns[3339] = 29'b0_000110100001_011_0_011010000100;
      patterns[3340] = 29'b0_000110100001_100_1_000011010000;
      patterns[3341] = 29'b0_000110100001_101_0_100001101000;
      patterns[3342] = 29'b0_000110100001_110_0_000110100001;
      patterns[3343] = 29'b0_000110100001_111_0_000110100001;
      patterns[3344] = 29'b0_000110100010_000_0_000110100010;
      patterns[3345] = 29'b0_000110100010_001_0_100010000110;
      patterns[3346] = 29'b0_000110100010_010_0_001101000100;
      patterns[3347] = 29'b0_000110100010_011_0_011010001000;
      patterns[3348] = 29'b0_000110100010_100_0_000011010001;
      patterns[3349] = 29'b0_000110100010_101_1_000001101000;
      patterns[3350] = 29'b0_000110100010_110_0_000110100010;
      patterns[3351] = 29'b0_000110100010_111_0_000110100010;
      patterns[3352] = 29'b0_000110100011_000_0_000110100011;
      patterns[3353] = 29'b0_000110100011_001_0_100011000110;
      patterns[3354] = 29'b0_000110100011_010_0_001101000110;
      patterns[3355] = 29'b0_000110100011_011_0_011010001100;
      patterns[3356] = 29'b0_000110100011_100_1_000011010001;
      patterns[3357] = 29'b0_000110100011_101_1_100001101000;
      patterns[3358] = 29'b0_000110100011_110_0_000110100011;
      patterns[3359] = 29'b0_000110100011_111_0_000110100011;
      patterns[3360] = 29'b0_000110100100_000_0_000110100100;
      patterns[3361] = 29'b0_000110100100_001_0_100100000110;
      patterns[3362] = 29'b0_000110100100_010_0_001101001000;
      patterns[3363] = 29'b0_000110100100_011_0_011010010000;
      patterns[3364] = 29'b0_000110100100_100_0_000011010010;
      patterns[3365] = 29'b0_000110100100_101_0_000001101001;
      patterns[3366] = 29'b0_000110100100_110_0_000110100100;
      patterns[3367] = 29'b0_000110100100_111_0_000110100100;
      patterns[3368] = 29'b0_000110100101_000_0_000110100101;
      patterns[3369] = 29'b0_000110100101_001_0_100101000110;
      patterns[3370] = 29'b0_000110100101_010_0_001101001010;
      patterns[3371] = 29'b0_000110100101_011_0_011010010100;
      patterns[3372] = 29'b0_000110100101_100_1_000011010010;
      patterns[3373] = 29'b0_000110100101_101_0_100001101001;
      patterns[3374] = 29'b0_000110100101_110_0_000110100101;
      patterns[3375] = 29'b0_000110100101_111_0_000110100101;
      patterns[3376] = 29'b0_000110100110_000_0_000110100110;
      patterns[3377] = 29'b0_000110100110_001_0_100110000110;
      patterns[3378] = 29'b0_000110100110_010_0_001101001100;
      patterns[3379] = 29'b0_000110100110_011_0_011010011000;
      patterns[3380] = 29'b0_000110100110_100_0_000011010011;
      patterns[3381] = 29'b0_000110100110_101_1_000001101001;
      patterns[3382] = 29'b0_000110100110_110_0_000110100110;
      patterns[3383] = 29'b0_000110100110_111_0_000110100110;
      patterns[3384] = 29'b0_000110100111_000_0_000110100111;
      patterns[3385] = 29'b0_000110100111_001_0_100111000110;
      patterns[3386] = 29'b0_000110100111_010_0_001101001110;
      patterns[3387] = 29'b0_000110100111_011_0_011010011100;
      patterns[3388] = 29'b0_000110100111_100_1_000011010011;
      patterns[3389] = 29'b0_000110100111_101_1_100001101001;
      patterns[3390] = 29'b0_000110100111_110_0_000110100111;
      patterns[3391] = 29'b0_000110100111_111_0_000110100111;
      patterns[3392] = 29'b0_000110101000_000_0_000110101000;
      patterns[3393] = 29'b0_000110101000_001_0_101000000110;
      patterns[3394] = 29'b0_000110101000_010_0_001101010000;
      patterns[3395] = 29'b0_000110101000_011_0_011010100000;
      patterns[3396] = 29'b0_000110101000_100_0_000011010100;
      patterns[3397] = 29'b0_000110101000_101_0_000001101010;
      patterns[3398] = 29'b0_000110101000_110_0_000110101000;
      patterns[3399] = 29'b0_000110101000_111_0_000110101000;
      patterns[3400] = 29'b0_000110101001_000_0_000110101001;
      patterns[3401] = 29'b0_000110101001_001_0_101001000110;
      patterns[3402] = 29'b0_000110101001_010_0_001101010010;
      patterns[3403] = 29'b0_000110101001_011_0_011010100100;
      patterns[3404] = 29'b0_000110101001_100_1_000011010100;
      patterns[3405] = 29'b0_000110101001_101_0_100001101010;
      patterns[3406] = 29'b0_000110101001_110_0_000110101001;
      patterns[3407] = 29'b0_000110101001_111_0_000110101001;
      patterns[3408] = 29'b0_000110101010_000_0_000110101010;
      patterns[3409] = 29'b0_000110101010_001_0_101010000110;
      patterns[3410] = 29'b0_000110101010_010_0_001101010100;
      patterns[3411] = 29'b0_000110101010_011_0_011010101000;
      patterns[3412] = 29'b0_000110101010_100_0_000011010101;
      patterns[3413] = 29'b0_000110101010_101_1_000001101010;
      patterns[3414] = 29'b0_000110101010_110_0_000110101010;
      patterns[3415] = 29'b0_000110101010_111_0_000110101010;
      patterns[3416] = 29'b0_000110101011_000_0_000110101011;
      patterns[3417] = 29'b0_000110101011_001_0_101011000110;
      patterns[3418] = 29'b0_000110101011_010_0_001101010110;
      patterns[3419] = 29'b0_000110101011_011_0_011010101100;
      patterns[3420] = 29'b0_000110101011_100_1_000011010101;
      patterns[3421] = 29'b0_000110101011_101_1_100001101010;
      patterns[3422] = 29'b0_000110101011_110_0_000110101011;
      patterns[3423] = 29'b0_000110101011_111_0_000110101011;
      patterns[3424] = 29'b0_000110101100_000_0_000110101100;
      patterns[3425] = 29'b0_000110101100_001_0_101100000110;
      patterns[3426] = 29'b0_000110101100_010_0_001101011000;
      patterns[3427] = 29'b0_000110101100_011_0_011010110000;
      patterns[3428] = 29'b0_000110101100_100_0_000011010110;
      patterns[3429] = 29'b0_000110101100_101_0_000001101011;
      patterns[3430] = 29'b0_000110101100_110_0_000110101100;
      patterns[3431] = 29'b0_000110101100_111_0_000110101100;
      patterns[3432] = 29'b0_000110101101_000_0_000110101101;
      patterns[3433] = 29'b0_000110101101_001_0_101101000110;
      patterns[3434] = 29'b0_000110101101_010_0_001101011010;
      patterns[3435] = 29'b0_000110101101_011_0_011010110100;
      patterns[3436] = 29'b0_000110101101_100_1_000011010110;
      patterns[3437] = 29'b0_000110101101_101_0_100001101011;
      patterns[3438] = 29'b0_000110101101_110_0_000110101101;
      patterns[3439] = 29'b0_000110101101_111_0_000110101101;
      patterns[3440] = 29'b0_000110101110_000_0_000110101110;
      patterns[3441] = 29'b0_000110101110_001_0_101110000110;
      patterns[3442] = 29'b0_000110101110_010_0_001101011100;
      patterns[3443] = 29'b0_000110101110_011_0_011010111000;
      patterns[3444] = 29'b0_000110101110_100_0_000011010111;
      patterns[3445] = 29'b0_000110101110_101_1_000001101011;
      patterns[3446] = 29'b0_000110101110_110_0_000110101110;
      patterns[3447] = 29'b0_000110101110_111_0_000110101110;
      patterns[3448] = 29'b0_000110101111_000_0_000110101111;
      patterns[3449] = 29'b0_000110101111_001_0_101111000110;
      patterns[3450] = 29'b0_000110101111_010_0_001101011110;
      patterns[3451] = 29'b0_000110101111_011_0_011010111100;
      patterns[3452] = 29'b0_000110101111_100_1_000011010111;
      patterns[3453] = 29'b0_000110101111_101_1_100001101011;
      patterns[3454] = 29'b0_000110101111_110_0_000110101111;
      patterns[3455] = 29'b0_000110101111_111_0_000110101111;
      patterns[3456] = 29'b0_000110110000_000_0_000110110000;
      patterns[3457] = 29'b0_000110110000_001_0_110000000110;
      patterns[3458] = 29'b0_000110110000_010_0_001101100000;
      patterns[3459] = 29'b0_000110110000_011_0_011011000000;
      patterns[3460] = 29'b0_000110110000_100_0_000011011000;
      patterns[3461] = 29'b0_000110110000_101_0_000001101100;
      patterns[3462] = 29'b0_000110110000_110_0_000110110000;
      patterns[3463] = 29'b0_000110110000_111_0_000110110000;
      patterns[3464] = 29'b0_000110110001_000_0_000110110001;
      patterns[3465] = 29'b0_000110110001_001_0_110001000110;
      patterns[3466] = 29'b0_000110110001_010_0_001101100010;
      patterns[3467] = 29'b0_000110110001_011_0_011011000100;
      patterns[3468] = 29'b0_000110110001_100_1_000011011000;
      patterns[3469] = 29'b0_000110110001_101_0_100001101100;
      patterns[3470] = 29'b0_000110110001_110_0_000110110001;
      patterns[3471] = 29'b0_000110110001_111_0_000110110001;
      patterns[3472] = 29'b0_000110110010_000_0_000110110010;
      patterns[3473] = 29'b0_000110110010_001_0_110010000110;
      patterns[3474] = 29'b0_000110110010_010_0_001101100100;
      patterns[3475] = 29'b0_000110110010_011_0_011011001000;
      patterns[3476] = 29'b0_000110110010_100_0_000011011001;
      patterns[3477] = 29'b0_000110110010_101_1_000001101100;
      patterns[3478] = 29'b0_000110110010_110_0_000110110010;
      patterns[3479] = 29'b0_000110110010_111_0_000110110010;
      patterns[3480] = 29'b0_000110110011_000_0_000110110011;
      patterns[3481] = 29'b0_000110110011_001_0_110011000110;
      patterns[3482] = 29'b0_000110110011_010_0_001101100110;
      patterns[3483] = 29'b0_000110110011_011_0_011011001100;
      patterns[3484] = 29'b0_000110110011_100_1_000011011001;
      patterns[3485] = 29'b0_000110110011_101_1_100001101100;
      patterns[3486] = 29'b0_000110110011_110_0_000110110011;
      patterns[3487] = 29'b0_000110110011_111_0_000110110011;
      patterns[3488] = 29'b0_000110110100_000_0_000110110100;
      patterns[3489] = 29'b0_000110110100_001_0_110100000110;
      patterns[3490] = 29'b0_000110110100_010_0_001101101000;
      patterns[3491] = 29'b0_000110110100_011_0_011011010000;
      patterns[3492] = 29'b0_000110110100_100_0_000011011010;
      patterns[3493] = 29'b0_000110110100_101_0_000001101101;
      patterns[3494] = 29'b0_000110110100_110_0_000110110100;
      patterns[3495] = 29'b0_000110110100_111_0_000110110100;
      patterns[3496] = 29'b0_000110110101_000_0_000110110101;
      patterns[3497] = 29'b0_000110110101_001_0_110101000110;
      patterns[3498] = 29'b0_000110110101_010_0_001101101010;
      patterns[3499] = 29'b0_000110110101_011_0_011011010100;
      patterns[3500] = 29'b0_000110110101_100_1_000011011010;
      patterns[3501] = 29'b0_000110110101_101_0_100001101101;
      patterns[3502] = 29'b0_000110110101_110_0_000110110101;
      patterns[3503] = 29'b0_000110110101_111_0_000110110101;
      patterns[3504] = 29'b0_000110110110_000_0_000110110110;
      patterns[3505] = 29'b0_000110110110_001_0_110110000110;
      patterns[3506] = 29'b0_000110110110_010_0_001101101100;
      patterns[3507] = 29'b0_000110110110_011_0_011011011000;
      patterns[3508] = 29'b0_000110110110_100_0_000011011011;
      patterns[3509] = 29'b0_000110110110_101_1_000001101101;
      patterns[3510] = 29'b0_000110110110_110_0_000110110110;
      patterns[3511] = 29'b0_000110110110_111_0_000110110110;
      patterns[3512] = 29'b0_000110110111_000_0_000110110111;
      patterns[3513] = 29'b0_000110110111_001_0_110111000110;
      patterns[3514] = 29'b0_000110110111_010_0_001101101110;
      patterns[3515] = 29'b0_000110110111_011_0_011011011100;
      patterns[3516] = 29'b0_000110110111_100_1_000011011011;
      patterns[3517] = 29'b0_000110110111_101_1_100001101101;
      patterns[3518] = 29'b0_000110110111_110_0_000110110111;
      patterns[3519] = 29'b0_000110110111_111_0_000110110111;
      patterns[3520] = 29'b0_000110111000_000_0_000110111000;
      patterns[3521] = 29'b0_000110111000_001_0_111000000110;
      patterns[3522] = 29'b0_000110111000_010_0_001101110000;
      patterns[3523] = 29'b0_000110111000_011_0_011011100000;
      patterns[3524] = 29'b0_000110111000_100_0_000011011100;
      patterns[3525] = 29'b0_000110111000_101_0_000001101110;
      patterns[3526] = 29'b0_000110111000_110_0_000110111000;
      patterns[3527] = 29'b0_000110111000_111_0_000110111000;
      patterns[3528] = 29'b0_000110111001_000_0_000110111001;
      patterns[3529] = 29'b0_000110111001_001_0_111001000110;
      patterns[3530] = 29'b0_000110111001_010_0_001101110010;
      patterns[3531] = 29'b0_000110111001_011_0_011011100100;
      patterns[3532] = 29'b0_000110111001_100_1_000011011100;
      patterns[3533] = 29'b0_000110111001_101_0_100001101110;
      patterns[3534] = 29'b0_000110111001_110_0_000110111001;
      patterns[3535] = 29'b0_000110111001_111_0_000110111001;
      patterns[3536] = 29'b0_000110111010_000_0_000110111010;
      patterns[3537] = 29'b0_000110111010_001_0_111010000110;
      patterns[3538] = 29'b0_000110111010_010_0_001101110100;
      patterns[3539] = 29'b0_000110111010_011_0_011011101000;
      patterns[3540] = 29'b0_000110111010_100_0_000011011101;
      patterns[3541] = 29'b0_000110111010_101_1_000001101110;
      patterns[3542] = 29'b0_000110111010_110_0_000110111010;
      patterns[3543] = 29'b0_000110111010_111_0_000110111010;
      patterns[3544] = 29'b0_000110111011_000_0_000110111011;
      patterns[3545] = 29'b0_000110111011_001_0_111011000110;
      patterns[3546] = 29'b0_000110111011_010_0_001101110110;
      patterns[3547] = 29'b0_000110111011_011_0_011011101100;
      patterns[3548] = 29'b0_000110111011_100_1_000011011101;
      patterns[3549] = 29'b0_000110111011_101_1_100001101110;
      patterns[3550] = 29'b0_000110111011_110_0_000110111011;
      patterns[3551] = 29'b0_000110111011_111_0_000110111011;
      patterns[3552] = 29'b0_000110111100_000_0_000110111100;
      patterns[3553] = 29'b0_000110111100_001_0_111100000110;
      patterns[3554] = 29'b0_000110111100_010_0_001101111000;
      patterns[3555] = 29'b0_000110111100_011_0_011011110000;
      patterns[3556] = 29'b0_000110111100_100_0_000011011110;
      patterns[3557] = 29'b0_000110111100_101_0_000001101111;
      patterns[3558] = 29'b0_000110111100_110_0_000110111100;
      patterns[3559] = 29'b0_000110111100_111_0_000110111100;
      patterns[3560] = 29'b0_000110111101_000_0_000110111101;
      patterns[3561] = 29'b0_000110111101_001_0_111101000110;
      patterns[3562] = 29'b0_000110111101_010_0_001101111010;
      patterns[3563] = 29'b0_000110111101_011_0_011011110100;
      patterns[3564] = 29'b0_000110111101_100_1_000011011110;
      patterns[3565] = 29'b0_000110111101_101_0_100001101111;
      patterns[3566] = 29'b0_000110111101_110_0_000110111101;
      patterns[3567] = 29'b0_000110111101_111_0_000110111101;
      patterns[3568] = 29'b0_000110111110_000_0_000110111110;
      patterns[3569] = 29'b0_000110111110_001_0_111110000110;
      patterns[3570] = 29'b0_000110111110_010_0_001101111100;
      patterns[3571] = 29'b0_000110111110_011_0_011011111000;
      patterns[3572] = 29'b0_000110111110_100_0_000011011111;
      patterns[3573] = 29'b0_000110111110_101_1_000001101111;
      patterns[3574] = 29'b0_000110111110_110_0_000110111110;
      patterns[3575] = 29'b0_000110111110_111_0_000110111110;
      patterns[3576] = 29'b0_000110111111_000_0_000110111111;
      patterns[3577] = 29'b0_000110111111_001_0_111111000110;
      patterns[3578] = 29'b0_000110111111_010_0_001101111110;
      patterns[3579] = 29'b0_000110111111_011_0_011011111100;
      patterns[3580] = 29'b0_000110111111_100_1_000011011111;
      patterns[3581] = 29'b0_000110111111_101_1_100001101111;
      patterns[3582] = 29'b0_000110111111_110_0_000110111111;
      patterns[3583] = 29'b0_000110111111_111_0_000110111111;
      patterns[3584] = 29'b0_000111000000_000_0_000111000000;
      patterns[3585] = 29'b0_000111000000_001_0_000000000111;
      patterns[3586] = 29'b0_000111000000_010_0_001110000000;
      patterns[3587] = 29'b0_000111000000_011_0_011100000000;
      patterns[3588] = 29'b0_000111000000_100_0_000011100000;
      patterns[3589] = 29'b0_000111000000_101_0_000001110000;
      patterns[3590] = 29'b0_000111000000_110_0_000111000000;
      patterns[3591] = 29'b0_000111000000_111_0_000111000000;
      patterns[3592] = 29'b0_000111000001_000_0_000111000001;
      patterns[3593] = 29'b0_000111000001_001_0_000001000111;
      patterns[3594] = 29'b0_000111000001_010_0_001110000010;
      patterns[3595] = 29'b0_000111000001_011_0_011100000100;
      patterns[3596] = 29'b0_000111000001_100_1_000011100000;
      patterns[3597] = 29'b0_000111000001_101_0_100001110000;
      patterns[3598] = 29'b0_000111000001_110_0_000111000001;
      patterns[3599] = 29'b0_000111000001_111_0_000111000001;
      patterns[3600] = 29'b0_000111000010_000_0_000111000010;
      patterns[3601] = 29'b0_000111000010_001_0_000010000111;
      patterns[3602] = 29'b0_000111000010_010_0_001110000100;
      patterns[3603] = 29'b0_000111000010_011_0_011100001000;
      patterns[3604] = 29'b0_000111000010_100_0_000011100001;
      patterns[3605] = 29'b0_000111000010_101_1_000001110000;
      patterns[3606] = 29'b0_000111000010_110_0_000111000010;
      patterns[3607] = 29'b0_000111000010_111_0_000111000010;
      patterns[3608] = 29'b0_000111000011_000_0_000111000011;
      patterns[3609] = 29'b0_000111000011_001_0_000011000111;
      patterns[3610] = 29'b0_000111000011_010_0_001110000110;
      patterns[3611] = 29'b0_000111000011_011_0_011100001100;
      patterns[3612] = 29'b0_000111000011_100_1_000011100001;
      patterns[3613] = 29'b0_000111000011_101_1_100001110000;
      patterns[3614] = 29'b0_000111000011_110_0_000111000011;
      patterns[3615] = 29'b0_000111000011_111_0_000111000011;
      patterns[3616] = 29'b0_000111000100_000_0_000111000100;
      patterns[3617] = 29'b0_000111000100_001_0_000100000111;
      patterns[3618] = 29'b0_000111000100_010_0_001110001000;
      patterns[3619] = 29'b0_000111000100_011_0_011100010000;
      patterns[3620] = 29'b0_000111000100_100_0_000011100010;
      patterns[3621] = 29'b0_000111000100_101_0_000001110001;
      patterns[3622] = 29'b0_000111000100_110_0_000111000100;
      patterns[3623] = 29'b0_000111000100_111_0_000111000100;
      patterns[3624] = 29'b0_000111000101_000_0_000111000101;
      patterns[3625] = 29'b0_000111000101_001_0_000101000111;
      patterns[3626] = 29'b0_000111000101_010_0_001110001010;
      patterns[3627] = 29'b0_000111000101_011_0_011100010100;
      patterns[3628] = 29'b0_000111000101_100_1_000011100010;
      patterns[3629] = 29'b0_000111000101_101_0_100001110001;
      patterns[3630] = 29'b0_000111000101_110_0_000111000101;
      patterns[3631] = 29'b0_000111000101_111_0_000111000101;
      patterns[3632] = 29'b0_000111000110_000_0_000111000110;
      patterns[3633] = 29'b0_000111000110_001_0_000110000111;
      patterns[3634] = 29'b0_000111000110_010_0_001110001100;
      patterns[3635] = 29'b0_000111000110_011_0_011100011000;
      patterns[3636] = 29'b0_000111000110_100_0_000011100011;
      patterns[3637] = 29'b0_000111000110_101_1_000001110001;
      patterns[3638] = 29'b0_000111000110_110_0_000111000110;
      patterns[3639] = 29'b0_000111000110_111_0_000111000110;
      patterns[3640] = 29'b0_000111000111_000_0_000111000111;
      patterns[3641] = 29'b0_000111000111_001_0_000111000111;
      patterns[3642] = 29'b0_000111000111_010_0_001110001110;
      patterns[3643] = 29'b0_000111000111_011_0_011100011100;
      patterns[3644] = 29'b0_000111000111_100_1_000011100011;
      patterns[3645] = 29'b0_000111000111_101_1_100001110001;
      patterns[3646] = 29'b0_000111000111_110_0_000111000111;
      patterns[3647] = 29'b0_000111000111_111_0_000111000111;
      patterns[3648] = 29'b0_000111001000_000_0_000111001000;
      patterns[3649] = 29'b0_000111001000_001_0_001000000111;
      patterns[3650] = 29'b0_000111001000_010_0_001110010000;
      patterns[3651] = 29'b0_000111001000_011_0_011100100000;
      patterns[3652] = 29'b0_000111001000_100_0_000011100100;
      patterns[3653] = 29'b0_000111001000_101_0_000001110010;
      patterns[3654] = 29'b0_000111001000_110_0_000111001000;
      patterns[3655] = 29'b0_000111001000_111_0_000111001000;
      patterns[3656] = 29'b0_000111001001_000_0_000111001001;
      patterns[3657] = 29'b0_000111001001_001_0_001001000111;
      patterns[3658] = 29'b0_000111001001_010_0_001110010010;
      patterns[3659] = 29'b0_000111001001_011_0_011100100100;
      patterns[3660] = 29'b0_000111001001_100_1_000011100100;
      patterns[3661] = 29'b0_000111001001_101_0_100001110010;
      patterns[3662] = 29'b0_000111001001_110_0_000111001001;
      patterns[3663] = 29'b0_000111001001_111_0_000111001001;
      patterns[3664] = 29'b0_000111001010_000_0_000111001010;
      patterns[3665] = 29'b0_000111001010_001_0_001010000111;
      patterns[3666] = 29'b0_000111001010_010_0_001110010100;
      patterns[3667] = 29'b0_000111001010_011_0_011100101000;
      patterns[3668] = 29'b0_000111001010_100_0_000011100101;
      patterns[3669] = 29'b0_000111001010_101_1_000001110010;
      patterns[3670] = 29'b0_000111001010_110_0_000111001010;
      patterns[3671] = 29'b0_000111001010_111_0_000111001010;
      patterns[3672] = 29'b0_000111001011_000_0_000111001011;
      patterns[3673] = 29'b0_000111001011_001_0_001011000111;
      patterns[3674] = 29'b0_000111001011_010_0_001110010110;
      patterns[3675] = 29'b0_000111001011_011_0_011100101100;
      patterns[3676] = 29'b0_000111001011_100_1_000011100101;
      patterns[3677] = 29'b0_000111001011_101_1_100001110010;
      patterns[3678] = 29'b0_000111001011_110_0_000111001011;
      patterns[3679] = 29'b0_000111001011_111_0_000111001011;
      patterns[3680] = 29'b0_000111001100_000_0_000111001100;
      patterns[3681] = 29'b0_000111001100_001_0_001100000111;
      patterns[3682] = 29'b0_000111001100_010_0_001110011000;
      patterns[3683] = 29'b0_000111001100_011_0_011100110000;
      patterns[3684] = 29'b0_000111001100_100_0_000011100110;
      patterns[3685] = 29'b0_000111001100_101_0_000001110011;
      patterns[3686] = 29'b0_000111001100_110_0_000111001100;
      patterns[3687] = 29'b0_000111001100_111_0_000111001100;
      patterns[3688] = 29'b0_000111001101_000_0_000111001101;
      patterns[3689] = 29'b0_000111001101_001_0_001101000111;
      patterns[3690] = 29'b0_000111001101_010_0_001110011010;
      patterns[3691] = 29'b0_000111001101_011_0_011100110100;
      patterns[3692] = 29'b0_000111001101_100_1_000011100110;
      patterns[3693] = 29'b0_000111001101_101_0_100001110011;
      patterns[3694] = 29'b0_000111001101_110_0_000111001101;
      patterns[3695] = 29'b0_000111001101_111_0_000111001101;
      patterns[3696] = 29'b0_000111001110_000_0_000111001110;
      patterns[3697] = 29'b0_000111001110_001_0_001110000111;
      patterns[3698] = 29'b0_000111001110_010_0_001110011100;
      patterns[3699] = 29'b0_000111001110_011_0_011100111000;
      patterns[3700] = 29'b0_000111001110_100_0_000011100111;
      patterns[3701] = 29'b0_000111001110_101_1_000001110011;
      patterns[3702] = 29'b0_000111001110_110_0_000111001110;
      patterns[3703] = 29'b0_000111001110_111_0_000111001110;
      patterns[3704] = 29'b0_000111001111_000_0_000111001111;
      patterns[3705] = 29'b0_000111001111_001_0_001111000111;
      patterns[3706] = 29'b0_000111001111_010_0_001110011110;
      patterns[3707] = 29'b0_000111001111_011_0_011100111100;
      patterns[3708] = 29'b0_000111001111_100_1_000011100111;
      patterns[3709] = 29'b0_000111001111_101_1_100001110011;
      patterns[3710] = 29'b0_000111001111_110_0_000111001111;
      patterns[3711] = 29'b0_000111001111_111_0_000111001111;
      patterns[3712] = 29'b0_000111010000_000_0_000111010000;
      patterns[3713] = 29'b0_000111010000_001_0_010000000111;
      patterns[3714] = 29'b0_000111010000_010_0_001110100000;
      patterns[3715] = 29'b0_000111010000_011_0_011101000000;
      patterns[3716] = 29'b0_000111010000_100_0_000011101000;
      patterns[3717] = 29'b0_000111010000_101_0_000001110100;
      patterns[3718] = 29'b0_000111010000_110_0_000111010000;
      patterns[3719] = 29'b0_000111010000_111_0_000111010000;
      patterns[3720] = 29'b0_000111010001_000_0_000111010001;
      patterns[3721] = 29'b0_000111010001_001_0_010001000111;
      patterns[3722] = 29'b0_000111010001_010_0_001110100010;
      patterns[3723] = 29'b0_000111010001_011_0_011101000100;
      patterns[3724] = 29'b0_000111010001_100_1_000011101000;
      patterns[3725] = 29'b0_000111010001_101_0_100001110100;
      patterns[3726] = 29'b0_000111010001_110_0_000111010001;
      patterns[3727] = 29'b0_000111010001_111_0_000111010001;
      patterns[3728] = 29'b0_000111010010_000_0_000111010010;
      patterns[3729] = 29'b0_000111010010_001_0_010010000111;
      patterns[3730] = 29'b0_000111010010_010_0_001110100100;
      patterns[3731] = 29'b0_000111010010_011_0_011101001000;
      patterns[3732] = 29'b0_000111010010_100_0_000011101001;
      patterns[3733] = 29'b0_000111010010_101_1_000001110100;
      patterns[3734] = 29'b0_000111010010_110_0_000111010010;
      patterns[3735] = 29'b0_000111010010_111_0_000111010010;
      patterns[3736] = 29'b0_000111010011_000_0_000111010011;
      patterns[3737] = 29'b0_000111010011_001_0_010011000111;
      patterns[3738] = 29'b0_000111010011_010_0_001110100110;
      patterns[3739] = 29'b0_000111010011_011_0_011101001100;
      patterns[3740] = 29'b0_000111010011_100_1_000011101001;
      patterns[3741] = 29'b0_000111010011_101_1_100001110100;
      patterns[3742] = 29'b0_000111010011_110_0_000111010011;
      patterns[3743] = 29'b0_000111010011_111_0_000111010011;
      patterns[3744] = 29'b0_000111010100_000_0_000111010100;
      patterns[3745] = 29'b0_000111010100_001_0_010100000111;
      patterns[3746] = 29'b0_000111010100_010_0_001110101000;
      patterns[3747] = 29'b0_000111010100_011_0_011101010000;
      patterns[3748] = 29'b0_000111010100_100_0_000011101010;
      patterns[3749] = 29'b0_000111010100_101_0_000001110101;
      patterns[3750] = 29'b0_000111010100_110_0_000111010100;
      patterns[3751] = 29'b0_000111010100_111_0_000111010100;
      patterns[3752] = 29'b0_000111010101_000_0_000111010101;
      patterns[3753] = 29'b0_000111010101_001_0_010101000111;
      patterns[3754] = 29'b0_000111010101_010_0_001110101010;
      patterns[3755] = 29'b0_000111010101_011_0_011101010100;
      patterns[3756] = 29'b0_000111010101_100_1_000011101010;
      patterns[3757] = 29'b0_000111010101_101_0_100001110101;
      patterns[3758] = 29'b0_000111010101_110_0_000111010101;
      patterns[3759] = 29'b0_000111010101_111_0_000111010101;
      patterns[3760] = 29'b0_000111010110_000_0_000111010110;
      patterns[3761] = 29'b0_000111010110_001_0_010110000111;
      patterns[3762] = 29'b0_000111010110_010_0_001110101100;
      patterns[3763] = 29'b0_000111010110_011_0_011101011000;
      patterns[3764] = 29'b0_000111010110_100_0_000011101011;
      patterns[3765] = 29'b0_000111010110_101_1_000001110101;
      patterns[3766] = 29'b0_000111010110_110_0_000111010110;
      patterns[3767] = 29'b0_000111010110_111_0_000111010110;
      patterns[3768] = 29'b0_000111010111_000_0_000111010111;
      patterns[3769] = 29'b0_000111010111_001_0_010111000111;
      patterns[3770] = 29'b0_000111010111_010_0_001110101110;
      patterns[3771] = 29'b0_000111010111_011_0_011101011100;
      patterns[3772] = 29'b0_000111010111_100_1_000011101011;
      patterns[3773] = 29'b0_000111010111_101_1_100001110101;
      patterns[3774] = 29'b0_000111010111_110_0_000111010111;
      patterns[3775] = 29'b0_000111010111_111_0_000111010111;
      patterns[3776] = 29'b0_000111011000_000_0_000111011000;
      patterns[3777] = 29'b0_000111011000_001_0_011000000111;
      patterns[3778] = 29'b0_000111011000_010_0_001110110000;
      patterns[3779] = 29'b0_000111011000_011_0_011101100000;
      patterns[3780] = 29'b0_000111011000_100_0_000011101100;
      patterns[3781] = 29'b0_000111011000_101_0_000001110110;
      patterns[3782] = 29'b0_000111011000_110_0_000111011000;
      patterns[3783] = 29'b0_000111011000_111_0_000111011000;
      patterns[3784] = 29'b0_000111011001_000_0_000111011001;
      patterns[3785] = 29'b0_000111011001_001_0_011001000111;
      patterns[3786] = 29'b0_000111011001_010_0_001110110010;
      patterns[3787] = 29'b0_000111011001_011_0_011101100100;
      patterns[3788] = 29'b0_000111011001_100_1_000011101100;
      patterns[3789] = 29'b0_000111011001_101_0_100001110110;
      patterns[3790] = 29'b0_000111011001_110_0_000111011001;
      patterns[3791] = 29'b0_000111011001_111_0_000111011001;
      patterns[3792] = 29'b0_000111011010_000_0_000111011010;
      patterns[3793] = 29'b0_000111011010_001_0_011010000111;
      patterns[3794] = 29'b0_000111011010_010_0_001110110100;
      patterns[3795] = 29'b0_000111011010_011_0_011101101000;
      patterns[3796] = 29'b0_000111011010_100_0_000011101101;
      patterns[3797] = 29'b0_000111011010_101_1_000001110110;
      patterns[3798] = 29'b0_000111011010_110_0_000111011010;
      patterns[3799] = 29'b0_000111011010_111_0_000111011010;
      patterns[3800] = 29'b0_000111011011_000_0_000111011011;
      patterns[3801] = 29'b0_000111011011_001_0_011011000111;
      patterns[3802] = 29'b0_000111011011_010_0_001110110110;
      patterns[3803] = 29'b0_000111011011_011_0_011101101100;
      patterns[3804] = 29'b0_000111011011_100_1_000011101101;
      patterns[3805] = 29'b0_000111011011_101_1_100001110110;
      patterns[3806] = 29'b0_000111011011_110_0_000111011011;
      patterns[3807] = 29'b0_000111011011_111_0_000111011011;
      patterns[3808] = 29'b0_000111011100_000_0_000111011100;
      patterns[3809] = 29'b0_000111011100_001_0_011100000111;
      patterns[3810] = 29'b0_000111011100_010_0_001110111000;
      patterns[3811] = 29'b0_000111011100_011_0_011101110000;
      patterns[3812] = 29'b0_000111011100_100_0_000011101110;
      patterns[3813] = 29'b0_000111011100_101_0_000001110111;
      patterns[3814] = 29'b0_000111011100_110_0_000111011100;
      patterns[3815] = 29'b0_000111011100_111_0_000111011100;
      patterns[3816] = 29'b0_000111011101_000_0_000111011101;
      patterns[3817] = 29'b0_000111011101_001_0_011101000111;
      patterns[3818] = 29'b0_000111011101_010_0_001110111010;
      patterns[3819] = 29'b0_000111011101_011_0_011101110100;
      patterns[3820] = 29'b0_000111011101_100_1_000011101110;
      patterns[3821] = 29'b0_000111011101_101_0_100001110111;
      patterns[3822] = 29'b0_000111011101_110_0_000111011101;
      patterns[3823] = 29'b0_000111011101_111_0_000111011101;
      patterns[3824] = 29'b0_000111011110_000_0_000111011110;
      patterns[3825] = 29'b0_000111011110_001_0_011110000111;
      patterns[3826] = 29'b0_000111011110_010_0_001110111100;
      patterns[3827] = 29'b0_000111011110_011_0_011101111000;
      patterns[3828] = 29'b0_000111011110_100_0_000011101111;
      patterns[3829] = 29'b0_000111011110_101_1_000001110111;
      patterns[3830] = 29'b0_000111011110_110_0_000111011110;
      patterns[3831] = 29'b0_000111011110_111_0_000111011110;
      patterns[3832] = 29'b0_000111011111_000_0_000111011111;
      patterns[3833] = 29'b0_000111011111_001_0_011111000111;
      patterns[3834] = 29'b0_000111011111_010_0_001110111110;
      patterns[3835] = 29'b0_000111011111_011_0_011101111100;
      patterns[3836] = 29'b0_000111011111_100_1_000011101111;
      patterns[3837] = 29'b0_000111011111_101_1_100001110111;
      patterns[3838] = 29'b0_000111011111_110_0_000111011111;
      patterns[3839] = 29'b0_000111011111_111_0_000111011111;
      patterns[3840] = 29'b0_000111100000_000_0_000111100000;
      patterns[3841] = 29'b0_000111100000_001_0_100000000111;
      patterns[3842] = 29'b0_000111100000_010_0_001111000000;
      patterns[3843] = 29'b0_000111100000_011_0_011110000000;
      patterns[3844] = 29'b0_000111100000_100_0_000011110000;
      patterns[3845] = 29'b0_000111100000_101_0_000001111000;
      patterns[3846] = 29'b0_000111100000_110_0_000111100000;
      patterns[3847] = 29'b0_000111100000_111_0_000111100000;
      patterns[3848] = 29'b0_000111100001_000_0_000111100001;
      patterns[3849] = 29'b0_000111100001_001_0_100001000111;
      patterns[3850] = 29'b0_000111100001_010_0_001111000010;
      patterns[3851] = 29'b0_000111100001_011_0_011110000100;
      patterns[3852] = 29'b0_000111100001_100_1_000011110000;
      patterns[3853] = 29'b0_000111100001_101_0_100001111000;
      patterns[3854] = 29'b0_000111100001_110_0_000111100001;
      patterns[3855] = 29'b0_000111100001_111_0_000111100001;
      patterns[3856] = 29'b0_000111100010_000_0_000111100010;
      patterns[3857] = 29'b0_000111100010_001_0_100010000111;
      patterns[3858] = 29'b0_000111100010_010_0_001111000100;
      patterns[3859] = 29'b0_000111100010_011_0_011110001000;
      patterns[3860] = 29'b0_000111100010_100_0_000011110001;
      patterns[3861] = 29'b0_000111100010_101_1_000001111000;
      patterns[3862] = 29'b0_000111100010_110_0_000111100010;
      patterns[3863] = 29'b0_000111100010_111_0_000111100010;
      patterns[3864] = 29'b0_000111100011_000_0_000111100011;
      patterns[3865] = 29'b0_000111100011_001_0_100011000111;
      patterns[3866] = 29'b0_000111100011_010_0_001111000110;
      patterns[3867] = 29'b0_000111100011_011_0_011110001100;
      patterns[3868] = 29'b0_000111100011_100_1_000011110001;
      patterns[3869] = 29'b0_000111100011_101_1_100001111000;
      patterns[3870] = 29'b0_000111100011_110_0_000111100011;
      patterns[3871] = 29'b0_000111100011_111_0_000111100011;
      patterns[3872] = 29'b0_000111100100_000_0_000111100100;
      patterns[3873] = 29'b0_000111100100_001_0_100100000111;
      patterns[3874] = 29'b0_000111100100_010_0_001111001000;
      patterns[3875] = 29'b0_000111100100_011_0_011110010000;
      patterns[3876] = 29'b0_000111100100_100_0_000011110010;
      patterns[3877] = 29'b0_000111100100_101_0_000001111001;
      patterns[3878] = 29'b0_000111100100_110_0_000111100100;
      patterns[3879] = 29'b0_000111100100_111_0_000111100100;
      patterns[3880] = 29'b0_000111100101_000_0_000111100101;
      patterns[3881] = 29'b0_000111100101_001_0_100101000111;
      patterns[3882] = 29'b0_000111100101_010_0_001111001010;
      patterns[3883] = 29'b0_000111100101_011_0_011110010100;
      patterns[3884] = 29'b0_000111100101_100_1_000011110010;
      patterns[3885] = 29'b0_000111100101_101_0_100001111001;
      patterns[3886] = 29'b0_000111100101_110_0_000111100101;
      patterns[3887] = 29'b0_000111100101_111_0_000111100101;
      patterns[3888] = 29'b0_000111100110_000_0_000111100110;
      patterns[3889] = 29'b0_000111100110_001_0_100110000111;
      patterns[3890] = 29'b0_000111100110_010_0_001111001100;
      patterns[3891] = 29'b0_000111100110_011_0_011110011000;
      patterns[3892] = 29'b0_000111100110_100_0_000011110011;
      patterns[3893] = 29'b0_000111100110_101_1_000001111001;
      patterns[3894] = 29'b0_000111100110_110_0_000111100110;
      patterns[3895] = 29'b0_000111100110_111_0_000111100110;
      patterns[3896] = 29'b0_000111100111_000_0_000111100111;
      patterns[3897] = 29'b0_000111100111_001_0_100111000111;
      patterns[3898] = 29'b0_000111100111_010_0_001111001110;
      patterns[3899] = 29'b0_000111100111_011_0_011110011100;
      patterns[3900] = 29'b0_000111100111_100_1_000011110011;
      patterns[3901] = 29'b0_000111100111_101_1_100001111001;
      patterns[3902] = 29'b0_000111100111_110_0_000111100111;
      patterns[3903] = 29'b0_000111100111_111_0_000111100111;
      patterns[3904] = 29'b0_000111101000_000_0_000111101000;
      patterns[3905] = 29'b0_000111101000_001_0_101000000111;
      patterns[3906] = 29'b0_000111101000_010_0_001111010000;
      patterns[3907] = 29'b0_000111101000_011_0_011110100000;
      patterns[3908] = 29'b0_000111101000_100_0_000011110100;
      patterns[3909] = 29'b0_000111101000_101_0_000001111010;
      patterns[3910] = 29'b0_000111101000_110_0_000111101000;
      patterns[3911] = 29'b0_000111101000_111_0_000111101000;
      patterns[3912] = 29'b0_000111101001_000_0_000111101001;
      patterns[3913] = 29'b0_000111101001_001_0_101001000111;
      patterns[3914] = 29'b0_000111101001_010_0_001111010010;
      patterns[3915] = 29'b0_000111101001_011_0_011110100100;
      patterns[3916] = 29'b0_000111101001_100_1_000011110100;
      patterns[3917] = 29'b0_000111101001_101_0_100001111010;
      patterns[3918] = 29'b0_000111101001_110_0_000111101001;
      patterns[3919] = 29'b0_000111101001_111_0_000111101001;
      patterns[3920] = 29'b0_000111101010_000_0_000111101010;
      patterns[3921] = 29'b0_000111101010_001_0_101010000111;
      patterns[3922] = 29'b0_000111101010_010_0_001111010100;
      patterns[3923] = 29'b0_000111101010_011_0_011110101000;
      patterns[3924] = 29'b0_000111101010_100_0_000011110101;
      patterns[3925] = 29'b0_000111101010_101_1_000001111010;
      patterns[3926] = 29'b0_000111101010_110_0_000111101010;
      patterns[3927] = 29'b0_000111101010_111_0_000111101010;
      patterns[3928] = 29'b0_000111101011_000_0_000111101011;
      patterns[3929] = 29'b0_000111101011_001_0_101011000111;
      patterns[3930] = 29'b0_000111101011_010_0_001111010110;
      patterns[3931] = 29'b0_000111101011_011_0_011110101100;
      patterns[3932] = 29'b0_000111101011_100_1_000011110101;
      patterns[3933] = 29'b0_000111101011_101_1_100001111010;
      patterns[3934] = 29'b0_000111101011_110_0_000111101011;
      patterns[3935] = 29'b0_000111101011_111_0_000111101011;
      patterns[3936] = 29'b0_000111101100_000_0_000111101100;
      patterns[3937] = 29'b0_000111101100_001_0_101100000111;
      patterns[3938] = 29'b0_000111101100_010_0_001111011000;
      patterns[3939] = 29'b0_000111101100_011_0_011110110000;
      patterns[3940] = 29'b0_000111101100_100_0_000011110110;
      patterns[3941] = 29'b0_000111101100_101_0_000001111011;
      patterns[3942] = 29'b0_000111101100_110_0_000111101100;
      patterns[3943] = 29'b0_000111101100_111_0_000111101100;
      patterns[3944] = 29'b0_000111101101_000_0_000111101101;
      patterns[3945] = 29'b0_000111101101_001_0_101101000111;
      patterns[3946] = 29'b0_000111101101_010_0_001111011010;
      patterns[3947] = 29'b0_000111101101_011_0_011110110100;
      patterns[3948] = 29'b0_000111101101_100_1_000011110110;
      patterns[3949] = 29'b0_000111101101_101_0_100001111011;
      patterns[3950] = 29'b0_000111101101_110_0_000111101101;
      patterns[3951] = 29'b0_000111101101_111_0_000111101101;
      patterns[3952] = 29'b0_000111101110_000_0_000111101110;
      patterns[3953] = 29'b0_000111101110_001_0_101110000111;
      patterns[3954] = 29'b0_000111101110_010_0_001111011100;
      patterns[3955] = 29'b0_000111101110_011_0_011110111000;
      patterns[3956] = 29'b0_000111101110_100_0_000011110111;
      patterns[3957] = 29'b0_000111101110_101_1_000001111011;
      patterns[3958] = 29'b0_000111101110_110_0_000111101110;
      patterns[3959] = 29'b0_000111101110_111_0_000111101110;
      patterns[3960] = 29'b0_000111101111_000_0_000111101111;
      patterns[3961] = 29'b0_000111101111_001_0_101111000111;
      patterns[3962] = 29'b0_000111101111_010_0_001111011110;
      patterns[3963] = 29'b0_000111101111_011_0_011110111100;
      patterns[3964] = 29'b0_000111101111_100_1_000011110111;
      patterns[3965] = 29'b0_000111101111_101_1_100001111011;
      patterns[3966] = 29'b0_000111101111_110_0_000111101111;
      patterns[3967] = 29'b0_000111101111_111_0_000111101111;
      patterns[3968] = 29'b0_000111110000_000_0_000111110000;
      patterns[3969] = 29'b0_000111110000_001_0_110000000111;
      patterns[3970] = 29'b0_000111110000_010_0_001111100000;
      patterns[3971] = 29'b0_000111110000_011_0_011111000000;
      patterns[3972] = 29'b0_000111110000_100_0_000011111000;
      patterns[3973] = 29'b0_000111110000_101_0_000001111100;
      patterns[3974] = 29'b0_000111110000_110_0_000111110000;
      patterns[3975] = 29'b0_000111110000_111_0_000111110000;
      patterns[3976] = 29'b0_000111110001_000_0_000111110001;
      patterns[3977] = 29'b0_000111110001_001_0_110001000111;
      patterns[3978] = 29'b0_000111110001_010_0_001111100010;
      patterns[3979] = 29'b0_000111110001_011_0_011111000100;
      patterns[3980] = 29'b0_000111110001_100_1_000011111000;
      patterns[3981] = 29'b0_000111110001_101_0_100001111100;
      patterns[3982] = 29'b0_000111110001_110_0_000111110001;
      patterns[3983] = 29'b0_000111110001_111_0_000111110001;
      patterns[3984] = 29'b0_000111110010_000_0_000111110010;
      patterns[3985] = 29'b0_000111110010_001_0_110010000111;
      patterns[3986] = 29'b0_000111110010_010_0_001111100100;
      patterns[3987] = 29'b0_000111110010_011_0_011111001000;
      patterns[3988] = 29'b0_000111110010_100_0_000011111001;
      patterns[3989] = 29'b0_000111110010_101_1_000001111100;
      patterns[3990] = 29'b0_000111110010_110_0_000111110010;
      patterns[3991] = 29'b0_000111110010_111_0_000111110010;
      patterns[3992] = 29'b0_000111110011_000_0_000111110011;
      patterns[3993] = 29'b0_000111110011_001_0_110011000111;
      patterns[3994] = 29'b0_000111110011_010_0_001111100110;
      patterns[3995] = 29'b0_000111110011_011_0_011111001100;
      patterns[3996] = 29'b0_000111110011_100_1_000011111001;
      patterns[3997] = 29'b0_000111110011_101_1_100001111100;
      patterns[3998] = 29'b0_000111110011_110_0_000111110011;
      patterns[3999] = 29'b0_000111110011_111_0_000111110011;
      patterns[4000] = 29'b0_000111110100_000_0_000111110100;
      patterns[4001] = 29'b0_000111110100_001_0_110100000111;
      patterns[4002] = 29'b0_000111110100_010_0_001111101000;
      patterns[4003] = 29'b0_000111110100_011_0_011111010000;
      patterns[4004] = 29'b0_000111110100_100_0_000011111010;
      patterns[4005] = 29'b0_000111110100_101_0_000001111101;
      patterns[4006] = 29'b0_000111110100_110_0_000111110100;
      patterns[4007] = 29'b0_000111110100_111_0_000111110100;
      patterns[4008] = 29'b0_000111110101_000_0_000111110101;
      patterns[4009] = 29'b0_000111110101_001_0_110101000111;
      patterns[4010] = 29'b0_000111110101_010_0_001111101010;
      patterns[4011] = 29'b0_000111110101_011_0_011111010100;
      patterns[4012] = 29'b0_000111110101_100_1_000011111010;
      patterns[4013] = 29'b0_000111110101_101_0_100001111101;
      patterns[4014] = 29'b0_000111110101_110_0_000111110101;
      patterns[4015] = 29'b0_000111110101_111_0_000111110101;
      patterns[4016] = 29'b0_000111110110_000_0_000111110110;
      patterns[4017] = 29'b0_000111110110_001_0_110110000111;
      patterns[4018] = 29'b0_000111110110_010_0_001111101100;
      patterns[4019] = 29'b0_000111110110_011_0_011111011000;
      patterns[4020] = 29'b0_000111110110_100_0_000011111011;
      patterns[4021] = 29'b0_000111110110_101_1_000001111101;
      patterns[4022] = 29'b0_000111110110_110_0_000111110110;
      patterns[4023] = 29'b0_000111110110_111_0_000111110110;
      patterns[4024] = 29'b0_000111110111_000_0_000111110111;
      patterns[4025] = 29'b0_000111110111_001_0_110111000111;
      patterns[4026] = 29'b0_000111110111_010_0_001111101110;
      patterns[4027] = 29'b0_000111110111_011_0_011111011100;
      patterns[4028] = 29'b0_000111110111_100_1_000011111011;
      patterns[4029] = 29'b0_000111110111_101_1_100001111101;
      patterns[4030] = 29'b0_000111110111_110_0_000111110111;
      patterns[4031] = 29'b0_000111110111_111_0_000111110111;
      patterns[4032] = 29'b0_000111111000_000_0_000111111000;
      patterns[4033] = 29'b0_000111111000_001_0_111000000111;
      patterns[4034] = 29'b0_000111111000_010_0_001111110000;
      patterns[4035] = 29'b0_000111111000_011_0_011111100000;
      patterns[4036] = 29'b0_000111111000_100_0_000011111100;
      patterns[4037] = 29'b0_000111111000_101_0_000001111110;
      patterns[4038] = 29'b0_000111111000_110_0_000111111000;
      patterns[4039] = 29'b0_000111111000_111_0_000111111000;
      patterns[4040] = 29'b0_000111111001_000_0_000111111001;
      patterns[4041] = 29'b0_000111111001_001_0_111001000111;
      patterns[4042] = 29'b0_000111111001_010_0_001111110010;
      patterns[4043] = 29'b0_000111111001_011_0_011111100100;
      patterns[4044] = 29'b0_000111111001_100_1_000011111100;
      patterns[4045] = 29'b0_000111111001_101_0_100001111110;
      patterns[4046] = 29'b0_000111111001_110_0_000111111001;
      patterns[4047] = 29'b0_000111111001_111_0_000111111001;
      patterns[4048] = 29'b0_000111111010_000_0_000111111010;
      patterns[4049] = 29'b0_000111111010_001_0_111010000111;
      patterns[4050] = 29'b0_000111111010_010_0_001111110100;
      patterns[4051] = 29'b0_000111111010_011_0_011111101000;
      patterns[4052] = 29'b0_000111111010_100_0_000011111101;
      patterns[4053] = 29'b0_000111111010_101_1_000001111110;
      patterns[4054] = 29'b0_000111111010_110_0_000111111010;
      patterns[4055] = 29'b0_000111111010_111_0_000111111010;
      patterns[4056] = 29'b0_000111111011_000_0_000111111011;
      patterns[4057] = 29'b0_000111111011_001_0_111011000111;
      patterns[4058] = 29'b0_000111111011_010_0_001111110110;
      patterns[4059] = 29'b0_000111111011_011_0_011111101100;
      patterns[4060] = 29'b0_000111111011_100_1_000011111101;
      patterns[4061] = 29'b0_000111111011_101_1_100001111110;
      patterns[4062] = 29'b0_000111111011_110_0_000111111011;
      patterns[4063] = 29'b0_000111111011_111_0_000111111011;
      patterns[4064] = 29'b0_000111111100_000_0_000111111100;
      patterns[4065] = 29'b0_000111111100_001_0_111100000111;
      patterns[4066] = 29'b0_000111111100_010_0_001111111000;
      patterns[4067] = 29'b0_000111111100_011_0_011111110000;
      patterns[4068] = 29'b0_000111111100_100_0_000011111110;
      patterns[4069] = 29'b0_000111111100_101_0_000001111111;
      patterns[4070] = 29'b0_000111111100_110_0_000111111100;
      patterns[4071] = 29'b0_000111111100_111_0_000111111100;
      patterns[4072] = 29'b0_000111111101_000_0_000111111101;
      patterns[4073] = 29'b0_000111111101_001_0_111101000111;
      patterns[4074] = 29'b0_000111111101_010_0_001111111010;
      patterns[4075] = 29'b0_000111111101_011_0_011111110100;
      patterns[4076] = 29'b0_000111111101_100_1_000011111110;
      patterns[4077] = 29'b0_000111111101_101_0_100001111111;
      patterns[4078] = 29'b0_000111111101_110_0_000111111101;
      patterns[4079] = 29'b0_000111111101_111_0_000111111101;
      patterns[4080] = 29'b0_000111111110_000_0_000111111110;
      patterns[4081] = 29'b0_000111111110_001_0_111110000111;
      patterns[4082] = 29'b0_000111111110_010_0_001111111100;
      patterns[4083] = 29'b0_000111111110_011_0_011111111000;
      patterns[4084] = 29'b0_000111111110_100_0_000011111111;
      patterns[4085] = 29'b0_000111111110_101_1_000001111111;
      patterns[4086] = 29'b0_000111111110_110_0_000111111110;
      patterns[4087] = 29'b0_000111111110_111_0_000111111110;
      patterns[4088] = 29'b0_000111111111_000_0_000111111111;
      patterns[4089] = 29'b0_000111111111_001_0_111111000111;
      patterns[4090] = 29'b0_000111111111_010_0_001111111110;
      patterns[4091] = 29'b0_000111111111_011_0_011111111100;
      patterns[4092] = 29'b0_000111111111_100_1_000011111111;
      patterns[4093] = 29'b0_000111111111_101_1_100001111111;
      patterns[4094] = 29'b0_000111111111_110_0_000111111111;
      patterns[4095] = 29'b0_000111111111_111_0_000111111111;
      patterns[4096] = 29'b0_001000000000_000_0_001000000000;
      patterns[4097] = 29'b0_001000000000_001_0_000000001000;
      patterns[4098] = 29'b0_001000000000_010_0_010000000000;
      patterns[4099] = 29'b0_001000000000_011_0_100000000000;
      patterns[4100] = 29'b0_001000000000_100_0_000100000000;
      patterns[4101] = 29'b0_001000000000_101_0_000010000000;
      patterns[4102] = 29'b0_001000000000_110_0_001000000000;
      patterns[4103] = 29'b0_001000000000_111_0_001000000000;
      patterns[4104] = 29'b0_001000000001_000_0_001000000001;
      patterns[4105] = 29'b0_001000000001_001_0_000001001000;
      patterns[4106] = 29'b0_001000000001_010_0_010000000010;
      patterns[4107] = 29'b0_001000000001_011_0_100000000100;
      patterns[4108] = 29'b0_001000000001_100_1_000100000000;
      patterns[4109] = 29'b0_001000000001_101_0_100010000000;
      patterns[4110] = 29'b0_001000000001_110_0_001000000001;
      patterns[4111] = 29'b0_001000000001_111_0_001000000001;
      patterns[4112] = 29'b0_001000000010_000_0_001000000010;
      patterns[4113] = 29'b0_001000000010_001_0_000010001000;
      patterns[4114] = 29'b0_001000000010_010_0_010000000100;
      patterns[4115] = 29'b0_001000000010_011_0_100000001000;
      patterns[4116] = 29'b0_001000000010_100_0_000100000001;
      patterns[4117] = 29'b0_001000000010_101_1_000010000000;
      patterns[4118] = 29'b0_001000000010_110_0_001000000010;
      patterns[4119] = 29'b0_001000000010_111_0_001000000010;
      patterns[4120] = 29'b0_001000000011_000_0_001000000011;
      patterns[4121] = 29'b0_001000000011_001_0_000011001000;
      patterns[4122] = 29'b0_001000000011_010_0_010000000110;
      patterns[4123] = 29'b0_001000000011_011_0_100000001100;
      patterns[4124] = 29'b0_001000000011_100_1_000100000001;
      patterns[4125] = 29'b0_001000000011_101_1_100010000000;
      patterns[4126] = 29'b0_001000000011_110_0_001000000011;
      patterns[4127] = 29'b0_001000000011_111_0_001000000011;
      patterns[4128] = 29'b0_001000000100_000_0_001000000100;
      patterns[4129] = 29'b0_001000000100_001_0_000100001000;
      patterns[4130] = 29'b0_001000000100_010_0_010000001000;
      patterns[4131] = 29'b0_001000000100_011_0_100000010000;
      patterns[4132] = 29'b0_001000000100_100_0_000100000010;
      patterns[4133] = 29'b0_001000000100_101_0_000010000001;
      patterns[4134] = 29'b0_001000000100_110_0_001000000100;
      patterns[4135] = 29'b0_001000000100_111_0_001000000100;
      patterns[4136] = 29'b0_001000000101_000_0_001000000101;
      patterns[4137] = 29'b0_001000000101_001_0_000101001000;
      patterns[4138] = 29'b0_001000000101_010_0_010000001010;
      patterns[4139] = 29'b0_001000000101_011_0_100000010100;
      patterns[4140] = 29'b0_001000000101_100_1_000100000010;
      patterns[4141] = 29'b0_001000000101_101_0_100010000001;
      patterns[4142] = 29'b0_001000000101_110_0_001000000101;
      patterns[4143] = 29'b0_001000000101_111_0_001000000101;
      patterns[4144] = 29'b0_001000000110_000_0_001000000110;
      patterns[4145] = 29'b0_001000000110_001_0_000110001000;
      patterns[4146] = 29'b0_001000000110_010_0_010000001100;
      patterns[4147] = 29'b0_001000000110_011_0_100000011000;
      patterns[4148] = 29'b0_001000000110_100_0_000100000011;
      patterns[4149] = 29'b0_001000000110_101_1_000010000001;
      patterns[4150] = 29'b0_001000000110_110_0_001000000110;
      patterns[4151] = 29'b0_001000000110_111_0_001000000110;
      patterns[4152] = 29'b0_001000000111_000_0_001000000111;
      patterns[4153] = 29'b0_001000000111_001_0_000111001000;
      patterns[4154] = 29'b0_001000000111_010_0_010000001110;
      patterns[4155] = 29'b0_001000000111_011_0_100000011100;
      patterns[4156] = 29'b0_001000000111_100_1_000100000011;
      patterns[4157] = 29'b0_001000000111_101_1_100010000001;
      patterns[4158] = 29'b0_001000000111_110_0_001000000111;
      patterns[4159] = 29'b0_001000000111_111_0_001000000111;
      patterns[4160] = 29'b0_001000001000_000_0_001000001000;
      patterns[4161] = 29'b0_001000001000_001_0_001000001000;
      patterns[4162] = 29'b0_001000001000_010_0_010000010000;
      patterns[4163] = 29'b0_001000001000_011_0_100000100000;
      patterns[4164] = 29'b0_001000001000_100_0_000100000100;
      patterns[4165] = 29'b0_001000001000_101_0_000010000010;
      patterns[4166] = 29'b0_001000001000_110_0_001000001000;
      patterns[4167] = 29'b0_001000001000_111_0_001000001000;
      patterns[4168] = 29'b0_001000001001_000_0_001000001001;
      patterns[4169] = 29'b0_001000001001_001_0_001001001000;
      patterns[4170] = 29'b0_001000001001_010_0_010000010010;
      patterns[4171] = 29'b0_001000001001_011_0_100000100100;
      patterns[4172] = 29'b0_001000001001_100_1_000100000100;
      patterns[4173] = 29'b0_001000001001_101_0_100010000010;
      patterns[4174] = 29'b0_001000001001_110_0_001000001001;
      patterns[4175] = 29'b0_001000001001_111_0_001000001001;
      patterns[4176] = 29'b0_001000001010_000_0_001000001010;
      patterns[4177] = 29'b0_001000001010_001_0_001010001000;
      patterns[4178] = 29'b0_001000001010_010_0_010000010100;
      patterns[4179] = 29'b0_001000001010_011_0_100000101000;
      patterns[4180] = 29'b0_001000001010_100_0_000100000101;
      patterns[4181] = 29'b0_001000001010_101_1_000010000010;
      patterns[4182] = 29'b0_001000001010_110_0_001000001010;
      patterns[4183] = 29'b0_001000001010_111_0_001000001010;
      patterns[4184] = 29'b0_001000001011_000_0_001000001011;
      patterns[4185] = 29'b0_001000001011_001_0_001011001000;
      patterns[4186] = 29'b0_001000001011_010_0_010000010110;
      patterns[4187] = 29'b0_001000001011_011_0_100000101100;
      patterns[4188] = 29'b0_001000001011_100_1_000100000101;
      patterns[4189] = 29'b0_001000001011_101_1_100010000010;
      patterns[4190] = 29'b0_001000001011_110_0_001000001011;
      patterns[4191] = 29'b0_001000001011_111_0_001000001011;
      patterns[4192] = 29'b0_001000001100_000_0_001000001100;
      patterns[4193] = 29'b0_001000001100_001_0_001100001000;
      patterns[4194] = 29'b0_001000001100_010_0_010000011000;
      patterns[4195] = 29'b0_001000001100_011_0_100000110000;
      patterns[4196] = 29'b0_001000001100_100_0_000100000110;
      patterns[4197] = 29'b0_001000001100_101_0_000010000011;
      patterns[4198] = 29'b0_001000001100_110_0_001000001100;
      patterns[4199] = 29'b0_001000001100_111_0_001000001100;
      patterns[4200] = 29'b0_001000001101_000_0_001000001101;
      patterns[4201] = 29'b0_001000001101_001_0_001101001000;
      patterns[4202] = 29'b0_001000001101_010_0_010000011010;
      patterns[4203] = 29'b0_001000001101_011_0_100000110100;
      patterns[4204] = 29'b0_001000001101_100_1_000100000110;
      patterns[4205] = 29'b0_001000001101_101_0_100010000011;
      patterns[4206] = 29'b0_001000001101_110_0_001000001101;
      patterns[4207] = 29'b0_001000001101_111_0_001000001101;
      patterns[4208] = 29'b0_001000001110_000_0_001000001110;
      patterns[4209] = 29'b0_001000001110_001_0_001110001000;
      patterns[4210] = 29'b0_001000001110_010_0_010000011100;
      patterns[4211] = 29'b0_001000001110_011_0_100000111000;
      patterns[4212] = 29'b0_001000001110_100_0_000100000111;
      patterns[4213] = 29'b0_001000001110_101_1_000010000011;
      patterns[4214] = 29'b0_001000001110_110_0_001000001110;
      patterns[4215] = 29'b0_001000001110_111_0_001000001110;
      patterns[4216] = 29'b0_001000001111_000_0_001000001111;
      patterns[4217] = 29'b0_001000001111_001_0_001111001000;
      patterns[4218] = 29'b0_001000001111_010_0_010000011110;
      patterns[4219] = 29'b0_001000001111_011_0_100000111100;
      patterns[4220] = 29'b0_001000001111_100_1_000100000111;
      patterns[4221] = 29'b0_001000001111_101_1_100010000011;
      patterns[4222] = 29'b0_001000001111_110_0_001000001111;
      patterns[4223] = 29'b0_001000001111_111_0_001000001111;
      patterns[4224] = 29'b0_001000010000_000_0_001000010000;
      patterns[4225] = 29'b0_001000010000_001_0_010000001000;
      patterns[4226] = 29'b0_001000010000_010_0_010000100000;
      patterns[4227] = 29'b0_001000010000_011_0_100001000000;
      patterns[4228] = 29'b0_001000010000_100_0_000100001000;
      patterns[4229] = 29'b0_001000010000_101_0_000010000100;
      patterns[4230] = 29'b0_001000010000_110_0_001000010000;
      patterns[4231] = 29'b0_001000010000_111_0_001000010000;
      patterns[4232] = 29'b0_001000010001_000_0_001000010001;
      patterns[4233] = 29'b0_001000010001_001_0_010001001000;
      patterns[4234] = 29'b0_001000010001_010_0_010000100010;
      patterns[4235] = 29'b0_001000010001_011_0_100001000100;
      patterns[4236] = 29'b0_001000010001_100_1_000100001000;
      patterns[4237] = 29'b0_001000010001_101_0_100010000100;
      patterns[4238] = 29'b0_001000010001_110_0_001000010001;
      patterns[4239] = 29'b0_001000010001_111_0_001000010001;
      patterns[4240] = 29'b0_001000010010_000_0_001000010010;
      patterns[4241] = 29'b0_001000010010_001_0_010010001000;
      patterns[4242] = 29'b0_001000010010_010_0_010000100100;
      patterns[4243] = 29'b0_001000010010_011_0_100001001000;
      patterns[4244] = 29'b0_001000010010_100_0_000100001001;
      patterns[4245] = 29'b0_001000010010_101_1_000010000100;
      patterns[4246] = 29'b0_001000010010_110_0_001000010010;
      patterns[4247] = 29'b0_001000010010_111_0_001000010010;
      patterns[4248] = 29'b0_001000010011_000_0_001000010011;
      patterns[4249] = 29'b0_001000010011_001_0_010011001000;
      patterns[4250] = 29'b0_001000010011_010_0_010000100110;
      patterns[4251] = 29'b0_001000010011_011_0_100001001100;
      patterns[4252] = 29'b0_001000010011_100_1_000100001001;
      patterns[4253] = 29'b0_001000010011_101_1_100010000100;
      patterns[4254] = 29'b0_001000010011_110_0_001000010011;
      patterns[4255] = 29'b0_001000010011_111_0_001000010011;
      patterns[4256] = 29'b0_001000010100_000_0_001000010100;
      patterns[4257] = 29'b0_001000010100_001_0_010100001000;
      patterns[4258] = 29'b0_001000010100_010_0_010000101000;
      patterns[4259] = 29'b0_001000010100_011_0_100001010000;
      patterns[4260] = 29'b0_001000010100_100_0_000100001010;
      patterns[4261] = 29'b0_001000010100_101_0_000010000101;
      patterns[4262] = 29'b0_001000010100_110_0_001000010100;
      patterns[4263] = 29'b0_001000010100_111_0_001000010100;
      patterns[4264] = 29'b0_001000010101_000_0_001000010101;
      patterns[4265] = 29'b0_001000010101_001_0_010101001000;
      patterns[4266] = 29'b0_001000010101_010_0_010000101010;
      patterns[4267] = 29'b0_001000010101_011_0_100001010100;
      patterns[4268] = 29'b0_001000010101_100_1_000100001010;
      patterns[4269] = 29'b0_001000010101_101_0_100010000101;
      patterns[4270] = 29'b0_001000010101_110_0_001000010101;
      patterns[4271] = 29'b0_001000010101_111_0_001000010101;
      patterns[4272] = 29'b0_001000010110_000_0_001000010110;
      patterns[4273] = 29'b0_001000010110_001_0_010110001000;
      patterns[4274] = 29'b0_001000010110_010_0_010000101100;
      patterns[4275] = 29'b0_001000010110_011_0_100001011000;
      patterns[4276] = 29'b0_001000010110_100_0_000100001011;
      patterns[4277] = 29'b0_001000010110_101_1_000010000101;
      patterns[4278] = 29'b0_001000010110_110_0_001000010110;
      patterns[4279] = 29'b0_001000010110_111_0_001000010110;
      patterns[4280] = 29'b0_001000010111_000_0_001000010111;
      patterns[4281] = 29'b0_001000010111_001_0_010111001000;
      patterns[4282] = 29'b0_001000010111_010_0_010000101110;
      patterns[4283] = 29'b0_001000010111_011_0_100001011100;
      patterns[4284] = 29'b0_001000010111_100_1_000100001011;
      patterns[4285] = 29'b0_001000010111_101_1_100010000101;
      patterns[4286] = 29'b0_001000010111_110_0_001000010111;
      patterns[4287] = 29'b0_001000010111_111_0_001000010111;
      patterns[4288] = 29'b0_001000011000_000_0_001000011000;
      patterns[4289] = 29'b0_001000011000_001_0_011000001000;
      patterns[4290] = 29'b0_001000011000_010_0_010000110000;
      patterns[4291] = 29'b0_001000011000_011_0_100001100000;
      patterns[4292] = 29'b0_001000011000_100_0_000100001100;
      patterns[4293] = 29'b0_001000011000_101_0_000010000110;
      patterns[4294] = 29'b0_001000011000_110_0_001000011000;
      patterns[4295] = 29'b0_001000011000_111_0_001000011000;
      patterns[4296] = 29'b0_001000011001_000_0_001000011001;
      patterns[4297] = 29'b0_001000011001_001_0_011001001000;
      patterns[4298] = 29'b0_001000011001_010_0_010000110010;
      patterns[4299] = 29'b0_001000011001_011_0_100001100100;
      patterns[4300] = 29'b0_001000011001_100_1_000100001100;
      patterns[4301] = 29'b0_001000011001_101_0_100010000110;
      patterns[4302] = 29'b0_001000011001_110_0_001000011001;
      patterns[4303] = 29'b0_001000011001_111_0_001000011001;
      patterns[4304] = 29'b0_001000011010_000_0_001000011010;
      patterns[4305] = 29'b0_001000011010_001_0_011010001000;
      patterns[4306] = 29'b0_001000011010_010_0_010000110100;
      patterns[4307] = 29'b0_001000011010_011_0_100001101000;
      patterns[4308] = 29'b0_001000011010_100_0_000100001101;
      patterns[4309] = 29'b0_001000011010_101_1_000010000110;
      patterns[4310] = 29'b0_001000011010_110_0_001000011010;
      patterns[4311] = 29'b0_001000011010_111_0_001000011010;
      patterns[4312] = 29'b0_001000011011_000_0_001000011011;
      patterns[4313] = 29'b0_001000011011_001_0_011011001000;
      patterns[4314] = 29'b0_001000011011_010_0_010000110110;
      patterns[4315] = 29'b0_001000011011_011_0_100001101100;
      patterns[4316] = 29'b0_001000011011_100_1_000100001101;
      patterns[4317] = 29'b0_001000011011_101_1_100010000110;
      patterns[4318] = 29'b0_001000011011_110_0_001000011011;
      patterns[4319] = 29'b0_001000011011_111_0_001000011011;
      patterns[4320] = 29'b0_001000011100_000_0_001000011100;
      patterns[4321] = 29'b0_001000011100_001_0_011100001000;
      patterns[4322] = 29'b0_001000011100_010_0_010000111000;
      patterns[4323] = 29'b0_001000011100_011_0_100001110000;
      patterns[4324] = 29'b0_001000011100_100_0_000100001110;
      patterns[4325] = 29'b0_001000011100_101_0_000010000111;
      patterns[4326] = 29'b0_001000011100_110_0_001000011100;
      patterns[4327] = 29'b0_001000011100_111_0_001000011100;
      patterns[4328] = 29'b0_001000011101_000_0_001000011101;
      patterns[4329] = 29'b0_001000011101_001_0_011101001000;
      patterns[4330] = 29'b0_001000011101_010_0_010000111010;
      patterns[4331] = 29'b0_001000011101_011_0_100001110100;
      patterns[4332] = 29'b0_001000011101_100_1_000100001110;
      patterns[4333] = 29'b0_001000011101_101_0_100010000111;
      patterns[4334] = 29'b0_001000011101_110_0_001000011101;
      patterns[4335] = 29'b0_001000011101_111_0_001000011101;
      patterns[4336] = 29'b0_001000011110_000_0_001000011110;
      patterns[4337] = 29'b0_001000011110_001_0_011110001000;
      patterns[4338] = 29'b0_001000011110_010_0_010000111100;
      patterns[4339] = 29'b0_001000011110_011_0_100001111000;
      patterns[4340] = 29'b0_001000011110_100_0_000100001111;
      patterns[4341] = 29'b0_001000011110_101_1_000010000111;
      patterns[4342] = 29'b0_001000011110_110_0_001000011110;
      patterns[4343] = 29'b0_001000011110_111_0_001000011110;
      patterns[4344] = 29'b0_001000011111_000_0_001000011111;
      patterns[4345] = 29'b0_001000011111_001_0_011111001000;
      patterns[4346] = 29'b0_001000011111_010_0_010000111110;
      patterns[4347] = 29'b0_001000011111_011_0_100001111100;
      patterns[4348] = 29'b0_001000011111_100_1_000100001111;
      patterns[4349] = 29'b0_001000011111_101_1_100010000111;
      patterns[4350] = 29'b0_001000011111_110_0_001000011111;
      patterns[4351] = 29'b0_001000011111_111_0_001000011111;
      patterns[4352] = 29'b0_001000100000_000_0_001000100000;
      patterns[4353] = 29'b0_001000100000_001_0_100000001000;
      patterns[4354] = 29'b0_001000100000_010_0_010001000000;
      patterns[4355] = 29'b0_001000100000_011_0_100010000000;
      patterns[4356] = 29'b0_001000100000_100_0_000100010000;
      patterns[4357] = 29'b0_001000100000_101_0_000010001000;
      patterns[4358] = 29'b0_001000100000_110_0_001000100000;
      patterns[4359] = 29'b0_001000100000_111_0_001000100000;
      patterns[4360] = 29'b0_001000100001_000_0_001000100001;
      patterns[4361] = 29'b0_001000100001_001_0_100001001000;
      patterns[4362] = 29'b0_001000100001_010_0_010001000010;
      patterns[4363] = 29'b0_001000100001_011_0_100010000100;
      patterns[4364] = 29'b0_001000100001_100_1_000100010000;
      patterns[4365] = 29'b0_001000100001_101_0_100010001000;
      patterns[4366] = 29'b0_001000100001_110_0_001000100001;
      patterns[4367] = 29'b0_001000100001_111_0_001000100001;
      patterns[4368] = 29'b0_001000100010_000_0_001000100010;
      patterns[4369] = 29'b0_001000100010_001_0_100010001000;
      patterns[4370] = 29'b0_001000100010_010_0_010001000100;
      patterns[4371] = 29'b0_001000100010_011_0_100010001000;
      patterns[4372] = 29'b0_001000100010_100_0_000100010001;
      patterns[4373] = 29'b0_001000100010_101_1_000010001000;
      patterns[4374] = 29'b0_001000100010_110_0_001000100010;
      patterns[4375] = 29'b0_001000100010_111_0_001000100010;
      patterns[4376] = 29'b0_001000100011_000_0_001000100011;
      patterns[4377] = 29'b0_001000100011_001_0_100011001000;
      patterns[4378] = 29'b0_001000100011_010_0_010001000110;
      patterns[4379] = 29'b0_001000100011_011_0_100010001100;
      patterns[4380] = 29'b0_001000100011_100_1_000100010001;
      patterns[4381] = 29'b0_001000100011_101_1_100010001000;
      patterns[4382] = 29'b0_001000100011_110_0_001000100011;
      patterns[4383] = 29'b0_001000100011_111_0_001000100011;
      patterns[4384] = 29'b0_001000100100_000_0_001000100100;
      patterns[4385] = 29'b0_001000100100_001_0_100100001000;
      patterns[4386] = 29'b0_001000100100_010_0_010001001000;
      patterns[4387] = 29'b0_001000100100_011_0_100010010000;
      patterns[4388] = 29'b0_001000100100_100_0_000100010010;
      patterns[4389] = 29'b0_001000100100_101_0_000010001001;
      patterns[4390] = 29'b0_001000100100_110_0_001000100100;
      patterns[4391] = 29'b0_001000100100_111_0_001000100100;
      patterns[4392] = 29'b0_001000100101_000_0_001000100101;
      patterns[4393] = 29'b0_001000100101_001_0_100101001000;
      patterns[4394] = 29'b0_001000100101_010_0_010001001010;
      patterns[4395] = 29'b0_001000100101_011_0_100010010100;
      patterns[4396] = 29'b0_001000100101_100_1_000100010010;
      patterns[4397] = 29'b0_001000100101_101_0_100010001001;
      patterns[4398] = 29'b0_001000100101_110_0_001000100101;
      patterns[4399] = 29'b0_001000100101_111_0_001000100101;
      patterns[4400] = 29'b0_001000100110_000_0_001000100110;
      patterns[4401] = 29'b0_001000100110_001_0_100110001000;
      patterns[4402] = 29'b0_001000100110_010_0_010001001100;
      patterns[4403] = 29'b0_001000100110_011_0_100010011000;
      patterns[4404] = 29'b0_001000100110_100_0_000100010011;
      patterns[4405] = 29'b0_001000100110_101_1_000010001001;
      patterns[4406] = 29'b0_001000100110_110_0_001000100110;
      patterns[4407] = 29'b0_001000100110_111_0_001000100110;
      patterns[4408] = 29'b0_001000100111_000_0_001000100111;
      patterns[4409] = 29'b0_001000100111_001_0_100111001000;
      patterns[4410] = 29'b0_001000100111_010_0_010001001110;
      patterns[4411] = 29'b0_001000100111_011_0_100010011100;
      patterns[4412] = 29'b0_001000100111_100_1_000100010011;
      patterns[4413] = 29'b0_001000100111_101_1_100010001001;
      patterns[4414] = 29'b0_001000100111_110_0_001000100111;
      patterns[4415] = 29'b0_001000100111_111_0_001000100111;
      patterns[4416] = 29'b0_001000101000_000_0_001000101000;
      patterns[4417] = 29'b0_001000101000_001_0_101000001000;
      patterns[4418] = 29'b0_001000101000_010_0_010001010000;
      patterns[4419] = 29'b0_001000101000_011_0_100010100000;
      patterns[4420] = 29'b0_001000101000_100_0_000100010100;
      patterns[4421] = 29'b0_001000101000_101_0_000010001010;
      patterns[4422] = 29'b0_001000101000_110_0_001000101000;
      patterns[4423] = 29'b0_001000101000_111_0_001000101000;
      patterns[4424] = 29'b0_001000101001_000_0_001000101001;
      patterns[4425] = 29'b0_001000101001_001_0_101001001000;
      patterns[4426] = 29'b0_001000101001_010_0_010001010010;
      patterns[4427] = 29'b0_001000101001_011_0_100010100100;
      patterns[4428] = 29'b0_001000101001_100_1_000100010100;
      patterns[4429] = 29'b0_001000101001_101_0_100010001010;
      patterns[4430] = 29'b0_001000101001_110_0_001000101001;
      patterns[4431] = 29'b0_001000101001_111_0_001000101001;
      patterns[4432] = 29'b0_001000101010_000_0_001000101010;
      patterns[4433] = 29'b0_001000101010_001_0_101010001000;
      patterns[4434] = 29'b0_001000101010_010_0_010001010100;
      patterns[4435] = 29'b0_001000101010_011_0_100010101000;
      patterns[4436] = 29'b0_001000101010_100_0_000100010101;
      patterns[4437] = 29'b0_001000101010_101_1_000010001010;
      patterns[4438] = 29'b0_001000101010_110_0_001000101010;
      patterns[4439] = 29'b0_001000101010_111_0_001000101010;
      patterns[4440] = 29'b0_001000101011_000_0_001000101011;
      patterns[4441] = 29'b0_001000101011_001_0_101011001000;
      patterns[4442] = 29'b0_001000101011_010_0_010001010110;
      patterns[4443] = 29'b0_001000101011_011_0_100010101100;
      patterns[4444] = 29'b0_001000101011_100_1_000100010101;
      patterns[4445] = 29'b0_001000101011_101_1_100010001010;
      patterns[4446] = 29'b0_001000101011_110_0_001000101011;
      patterns[4447] = 29'b0_001000101011_111_0_001000101011;
      patterns[4448] = 29'b0_001000101100_000_0_001000101100;
      patterns[4449] = 29'b0_001000101100_001_0_101100001000;
      patterns[4450] = 29'b0_001000101100_010_0_010001011000;
      patterns[4451] = 29'b0_001000101100_011_0_100010110000;
      patterns[4452] = 29'b0_001000101100_100_0_000100010110;
      patterns[4453] = 29'b0_001000101100_101_0_000010001011;
      patterns[4454] = 29'b0_001000101100_110_0_001000101100;
      patterns[4455] = 29'b0_001000101100_111_0_001000101100;
      patterns[4456] = 29'b0_001000101101_000_0_001000101101;
      patterns[4457] = 29'b0_001000101101_001_0_101101001000;
      patterns[4458] = 29'b0_001000101101_010_0_010001011010;
      patterns[4459] = 29'b0_001000101101_011_0_100010110100;
      patterns[4460] = 29'b0_001000101101_100_1_000100010110;
      patterns[4461] = 29'b0_001000101101_101_0_100010001011;
      patterns[4462] = 29'b0_001000101101_110_0_001000101101;
      patterns[4463] = 29'b0_001000101101_111_0_001000101101;
      patterns[4464] = 29'b0_001000101110_000_0_001000101110;
      patterns[4465] = 29'b0_001000101110_001_0_101110001000;
      patterns[4466] = 29'b0_001000101110_010_0_010001011100;
      patterns[4467] = 29'b0_001000101110_011_0_100010111000;
      patterns[4468] = 29'b0_001000101110_100_0_000100010111;
      patterns[4469] = 29'b0_001000101110_101_1_000010001011;
      patterns[4470] = 29'b0_001000101110_110_0_001000101110;
      patterns[4471] = 29'b0_001000101110_111_0_001000101110;
      patterns[4472] = 29'b0_001000101111_000_0_001000101111;
      patterns[4473] = 29'b0_001000101111_001_0_101111001000;
      patterns[4474] = 29'b0_001000101111_010_0_010001011110;
      patterns[4475] = 29'b0_001000101111_011_0_100010111100;
      patterns[4476] = 29'b0_001000101111_100_1_000100010111;
      patterns[4477] = 29'b0_001000101111_101_1_100010001011;
      patterns[4478] = 29'b0_001000101111_110_0_001000101111;
      patterns[4479] = 29'b0_001000101111_111_0_001000101111;
      patterns[4480] = 29'b0_001000110000_000_0_001000110000;
      patterns[4481] = 29'b0_001000110000_001_0_110000001000;
      patterns[4482] = 29'b0_001000110000_010_0_010001100000;
      patterns[4483] = 29'b0_001000110000_011_0_100011000000;
      patterns[4484] = 29'b0_001000110000_100_0_000100011000;
      patterns[4485] = 29'b0_001000110000_101_0_000010001100;
      patterns[4486] = 29'b0_001000110000_110_0_001000110000;
      patterns[4487] = 29'b0_001000110000_111_0_001000110000;
      patterns[4488] = 29'b0_001000110001_000_0_001000110001;
      patterns[4489] = 29'b0_001000110001_001_0_110001001000;
      patterns[4490] = 29'b0_001000110001_010_0_010001100010;
      patterns[4491] = 29'b0_001000110001_011_0_100011000100;
      patterns[4492] = 29'b0_001000110001_100_1_000100011000;
      patterns[4493] = 29'b0_001000110001_101_0_100010001100;
      patterns[4494] = 29'b0_001000110001_110_0_001000110001;
      patterns[4495] = 29'b0_001000110001_111_0_001000110001;
      patterns[4496] = 29'b0_001000110010_000_0_001000110010;
      patterns[4497] = 29'b0_001000110010_001_0_110010001000;
      patterns[4498] = 29'b0_001000110010_010_0_010001100100;
      patterns[4499] = 29'b0_001000110010_011_0_100011001000;
      patterns[4500] = 29'b0_001000110010_100_0_000100011001;
      patterns[4501] = 29'b0_001000110010_101_1_000010001100;
      patterns[4502] = 29'b0_001000110010_110_0_001000110010;
      patterns[4503] = 29'b0_001000110010_111_0_001000110010;
      patterns[4504] = 29'b0_001000110011_000_0_001000110011;
      patterns[4505] = 29'b0_001000110011_001_0_110011001000;
      patterns[4506] = 29'b0_001000110011_010_0_010001100110;
      patterns[4507] = 29'b0_001000110011_011_0_100011001100;
      patterns[4508] = 29'b0_001000110011_100_1_000100011001;
      patterns[4509] = 29'b0_001000110011_101_1_100010001100;
      patterns[4510] = 29'b0_001000110011_110_0_001000110011;
      patterns[4511] = 29'b0_001000110011_111_0_001000110011;
      patterns[4512] = 29'b0_001000110100_000_0_001000110100;
      patterns[4513] = 29'b0_001000110100_001_0_110100001000;
      patterns[4514] = 29'b0_001000110100_010_0_010001101000;
      patterns[4515] = 29'b0_001000110100_011_0_100011010000;
      patterns[4516] = 29'b0_001000110100_100_0_000100011010;
      patterns[4517] = 29'b0_001000110100_101_0_000010001101;
      patterns[4518] = 29'b0_001000110100_110_0_001000110100;
      patterns[4519] = 29'b0_001000110100_111_0_001000110100;
      patterns[4520] = 29'b0_001000110101_000_0_001000110101;
      patterns[4521] = 29'b0_001000110101_001_0_110101001000;
      patterns[4522] = 29'b0_001000110101_010_0_010001101010;
      patterns[4523] = 29'b0_001000110101_011_0_100011010100;
      patterns[4524] = 29'b0_001000110101_100_1_000100011010;
      patterns[4525] = 29'b0_001000110101_101_0_100010001101;
      patterns[4526] = 29'b0_001000110101_110_0_001000110101;
      patterns[4527] = 29'b0_001000110101_111_0_001000110101;
      patterns[4528] = 29'b0_001000110110_000_0_001000110110;
      patterns[4529] = 29'b0_001000110110_001_0_110110001000;
      patterns[4530] = 29'b0_001000110110_010_0_010001101100;
      patterns[4531] = 29'b0_001000110110_011_0_100011011000;
      patterns[4532] = 29'b0_001000110110_100_0_000100011011;
      patterns[4533] = 29'b0_001000110110_101_1_000010001101;
      patterns[4534] = 29'b0_001000110110_110_0_001000110110;
      patterns[4535] = 29'b0_001000110110_111_0_001000110110;
      patterns[4536] = 29'b0_001000110111_000_0_001000110111;
      patterns[4537] = 29'b0_001000110111_001_0_110111001000;
      patterns[4538] = 29'b0_001000110111_010_0_010001101110;
      patterns[4539] = 29'b0_001000110111_011_0_100011011100;
      patterns[4540] = 29'b0_001000110111_100_1_000100011011;
      patterns[4541] = 29'b0_001000110111_101_1_100010001101;
      patterns[4542] = 29'b0_001000110111_110_0_001000110111;
      patterns[4543] = 29'b0_001000110111_111_0_001000110111;
      patterns[4544] = 29'b0_001000111000_000_0_001000111000;
      patterns[4545] = 29'b0_001000111000_001_0_111000001000;
      patterns[4546] = 29'b0_001000111000_010_0_010001110000;
      patterns[4547] = 29'b0_001000111000_011_0_100011100000;
      patterns[4548] = 29'b0_001000111000_100_0_000100011100;
      patterns[4549] = 29'b0_001000111000_101_0_000010001110;
      patterns[4550] = 29'b0_001000111000_110_0_001000111000;
      patterns[4551] = 29'b0_001000111000_111_0_001000111000;
      patterns[4552] = 29'b0_001000111001_000_0_001000111001;
      patterns[4553] = 29'b0_001000111001_001_0_111001001000;
      patterns[4554] = 29'b0_001000111001_010_0_010001110010;
      patterns[4555] = 29'b0_001000111001_011_0_100011100100;
      patterns[4556] = 29'b0_001000111001_100_1_000100011100;
      patterns[4557] = 29'b0_001000111001_101_0_100010001110;
      patterns[4558] = 29'b0_001000111001_110_0_001000111001;
      patterns[4559] = 29'b0_001000111001_111_0_001000111001;
      patterns[4560] = 29'b0_001000111010_000_0_001000111010;
      patterns[4561] = 29'b0_001000111010_001_0_111010001000;
      patterns[4562] = 29'b0_001000111010_010_0_010001110100;
      patterns[4563] = 29'b0_001000111010_011_0_100011101000;
      patterns[4564] = 29'b0_001000111010_100_0_000100011101;
      patterns[4565] = 29'b0_001000111010_101_1_000010001110;
      patterns[4566] = 29'b0_001000111010_110_0_001000111010;
      patterns[4567] = 29'b0_001000111010_111_0_001000111010;
      patterns[4568] = 29'b0_001000111011_000_0_001000111011;
      patterns[4569] = 29'b0_001000111011_001_0_111011001000;
      patterns[4570] = 29'b0_001000111011_010_0_010001110110;
      patterns[4571] = 29'b0_001000111011_011_0_100011101100;
      patterns[4572] = 29'b0_001000111011_100_1_000100011101;
      patterns[4573] = 29'b0_001000111011_101_1_100010001110;
      patterns[4574] = 29'b0_001000111011_110_0_001000111011;
      patterns[4575] = 29'b0_001000111011_111_0_001000111011;
      patterns[4576] = 29'b0_001000111100_000_0_001000111100;
      patterns[4577] = 29'b0_001000111100_001_0_111100001000;
      patterns[4578] = 29'b0_001000111100_010_0_010001111000;
      patterns[4579] = 29'b0_001000111100_011_0_100011110000;
      patterns[4580] = 29'b0_001000111100_100_0_000100011110;
      patterns[4581] = 29'b0_001000111100_101_0_000010001111;
      patterns[4582] = 29'b0_001000111100_110_0_001000111100;
      patterns[4583] = 29'b0_001000111100_111_0_001000111100;
      patterns[4584] = 29'b0_001000111101_000_0_001000111101;
      patterns[4585] = 29'b0_001000111101_001_0_111101001000;
      patterns[4586] = 29'b0_001000111101_010_0_010001111010;
      patterns[4587] = 29'b0_001000111101_011_0_100011110100;
      patterns[4588] = 29'b0_001000111101_100_1_000100011110;
      patterns[4589] = 29'b0_001000111101_101_0_100010001111;
      patterns[4590] = 29'b0_001000111101_110_0_001000111101;
      patterns[4591] = 29'b0_001000111101_111_0_001000111101;
      patterns[4592] = 29'b0_001000111110_000_0_001000111110;
      patterns[4593] = 29'b0_001000111110_001_0_111110001000;
      patterns[4594] = 29'b0_001000111110_010_0_010001111100;
      patterns[4595] = 29'b0_001000111110_011_0_100011111000;
      patterns[4596] = 29'b0_001000111110_100_0_000100011111;
      patterns[4597] = 29'b0_001000111110_101_1_000010001111;
      patterns[4598] = 29'b0_001000111110_110_0_001000111110;
      patterns[4599] = 29'b0_001000111110_111_0_001000111110;
      patterns[4600] = 29'b0_001000111111_000_0_001000111111;
      patterns[4601] = 29'b0_001000111111_001_0_111111001000;
      patterns[4602] = 29'b0_001000111111_010_0_010001111110;
      patterns[4603] = 29'b0_001000111111_011_0_100011111100;
      patterns[4604] = 29'b0_001000111111_100_1_000100011111;
      patterns[4605] = 29'b0_001000111111_101_1_100010001111;
      patterns[4606] = 29'b0_001000111111_110_0_001000111111;
      patterns[4607] = 29'b0_001000111111_111_0_001000111111;
      patterns[4608] = 29'b0_001001000000_000_0_001001000000;
      patterns[4609] = 29'b0_001001000000_001_0_000000001001;
      patterns[4610] = 29'b0_001001000000_010_0_010010000000;
      patterns[4611] = 29'b0_001001000000_011_0_100100000000;
      patterns[4612] = 29'b0_001001000000_100_0_000100100000;
      patterns[4613] = 29'b0_001001000000_101_0_000010010000;
      patterns[4614] = 29'b0_001001000000_110_0_001001000000;
      patterns[4615] = 29'b0_001001000000_111_0_001001000000;
      patterns[4616] = 29'b0_001001000001_000_0_001001000001;
      patterns[4617] = 29'b0_001001000001_001_0_000001001001;
      patterns[4618] = 29'b0_001001000001_010_0_010010000010;
      patterns[4619] = 29'b0_001001000001_011_0_100100000100;
      patterns[4620] = 29'b0_001001000001_100_1_000100100000;
      patterns[4621] = 29'b0_001001000001_101_0_100010010000;
      patterns[4622] = 29'b0_001001000001_110_0_001001000001;
      patterns[4623] = 29'b0_001001000001_111_0_001001000001;
      patterns[4624] = 29'b0_001001000010_000_0_001001000010;
      patterns[4625] = 29'b0_001001000010_001_0_000010001001;
      patterns[4626] = 29'b0_001001000010_010_0_010010000100;
      patterns[4627] = 29'b0_001001000010_011_0_100100001000;
      patterns[4628] = 29'b0_001001000010_100_0_000100100001;
      patterns[4629] = 29'b0_001001000010_101_1_000010010000;
      patterns[4630] = 29'b0_001001000010_110_0_001001000010;
      patterns[4631] = 29'b0_001001000010_111_0_001001000010;
      patterns[4632] = 29'b0_001001000011_000_0_001001000011;
      patterns[4633] = 29'b0_001001000011_001_0_000011001001;
      patterns[4634] = 29'b0_001001000011_010_0_010010000110;
      patterns[4635] = 29'b0_001001000011_011_0_100100001100;
      patterns[4636] = 29'b0_001001000011_100_1_000100100001;
      patterns[4637] = 29'b0_001001000011_101_1_100010010000;
      patterns[4638] = 29'b0_001001000011_110_0_001001000011;
      patterns[4639] = 29'b0_001001000011_111_0_001001000011;
      patterns[4640] = 29'b0_001001000100_000_0_001001000100;
      patterns[4641] = 29'b0_001001000100_001_0_000100001001;
      patterns[4642] = 29'b0_001001000100_010_0_010010001000;
      patterns[4643] = 29'b0_001001000100_011_0_100100010000;
      patterns[4644] = 29'b0_001001000100_100_0_000100100010;
      patterns[4645] = 29'b0_001001000100_101_0_000010010001;
      patterns[4646] = 29'b0_001001000100_110_0_001001000100;
      patterns[4647] = 29'b0_001001000100_111_0_001001000100;
      patterns[4648] = 29'b0_001001000101_000_0_001001000101;
      patterns[4649] = 29'b0_001001000101_001_0_000101001001;
      patterns[4650] = 29'b0_001001000101_010_0_010010001010;
      patterns[4651] = 29'b0_001001000101_011_0_100100010100;
      patterns[4652] = 29'b0_001001000101_100_1_000100100010;
      patterns[4653] = 29'b0_001001000101_101_0_100010010001;
      patterns[4654] = 29'b0_001001000101_110_0_001001000101;
      patterns[4655] = 29'b0_001001000101_111_0_001001000101;
      patterns[4656] = 29'b0_001001000110_000_0_001001000110;
      patterns[4657] = 29'b0_001001000110_001_0_000110001001;
      patterns[4658] = 29'b0_001001000110_010_0_010010001100;
      patterns[4659] = 29'b0_001001000110_011_0_100100011000;
      patterns[4660] = 29'b0_001001000110_100_0_000100100011;
      patterns[4661] = 29'b0_001001000110_101_1_000010010001;
      patterns[4662] = 29'b0_001001000110_110_0_001001000110;
      patterns[4663] = 29'b0_001001000110_111_0_001001000110;
      patterns[4664] = 29'b0_001001000111_000_0_001001000111;
      patterns[4665] = 29'b0_001001000111_001_0_000111001001;
      patterns[4666] = 29'b0_001001000111_010_0_010010001110;
      patterns[4667] = 29'b0_001001000111_011_0_100100011100;
      patterns[4668] = 29'b0_001001000111_100_1_000100100011;
      patterns[4669] = 29'b0_001001000111_101_1_100010010001;
      patterns[4670] = 29'b0_001001000111_110_0_001001000111;
      patterns[4671] = 29'b0_001001000111_111_0_001001000111;
      patterns[4672] = 29'b0_001001001000_000_0_001001001000;
      patterns[4673] = 29'b0_001001001000_001_0_001000001001;
      patterns[4674] = 29'b0_001001001000_010_0_010010010000;
      patterns[4675] = 29'b0_001001001000_011_0_100100100000;
      patterns[4676] = 29'b0_001001001000_100_0_000100100100;
      patterns[4677] = 29'b0_001001001000_101_0_000010010010;
      patterns[4678] = 29'b0_001001001000_110_0_001001001000;
      patterns[4679] = 29'b0_001001001000_111_0_001001001000;
      patterns[4680] = 29'b0_001001001001_000_0_001001001001;
      patterns[4681] = 29'b0_001001001001_001_0_001001001001;
      patterns[4682] = 29'b0_001001001001_010_0_010010010010;
      patterns[4683] = 29'b0_001001001001_011_0_100100100100;
      patterns[4684] = 29'b0_001001001001_100_1_000100100100;
      patterns[4685] = 29'b0_001001001001_101_0_100010010010;
      patterns[4686] = 29'b0_001001001001_110_0_001001001001;
      patterns[4687] = 29'b0_001001001001_111_0_001001001001;
      patterns[4688] = 29'b0_001001001010_000_0_001001001010;
      patterns[4689] = 29'b0_001001001010_001_0_001010001001;
      patterns[4690] = 29'b0_001001001010_010_0_010010010100;
      patterns[4691] = 29'b0_001001001010_011_0_100100101000;
      patterns[4692] = 29'b0_001001001010_100_0_000100100101;
      patterns[4693] = 29'b0_001001001010_101_1_000010010010;
      patterns[4694] = 29'b0_001001001010_110_0_001001001010;
      patterns[4695] = 29'b0_001001001010_111_0_001001001010;
      patterns[4696] = 29'b0_001001001011_000_0_001001001011;
      patterns[4697] = 29'b0_001001001011_001_0_001011001001;
      patterns[4698] = 29'b0_001001001011_010_0_010010010110;
      patterns[4699] = 29'b0_001001001011_011_0_100100101100;
      patterns[4700] = 29'b0_001001001011_100_1_000100100101;
      patterns[4701] = 29'b0_001001001011_101_1_100010010010;
      patterns[4702] = 29'b0_001001001011_110_0_001001001011;
      patterns[4703] = 29'b0_001001001011_111_0_001001001011;
      patterns[4704] = 29'b0_001001001100_000_0_001001001100;
      patterns[4705] = 29'b0_001001001100_001_0_001100001001;
      patterns[4706] = 29'b0_001001001100_010_0_010010011000;
      patterns[4707] = 29'b0_001001001100_011_0_100100110000;
      patterns[4708] = 29'b0_001001001100_100_0_000100100110;
      patterns[4709] = 29'b0_001001001100_101_0_000010010011;
      patterns[4710] = 29'b0_001001001100_110_0_001001001100;
      patterns[4711] = 29'b0_001001001100_111_0_001001001100;
      patterns[4712] = 29'b0_001001001101_000_0_001001001101;
      patterns[4713] = 29'b0_001001001101_001_0_001101001001;
      patterns[4714] = 29'b0_001001001101_010_0_010010011010;
      patterns[4715] = 29'b0_001001001101_011_0_100100110100;
      patterns[4716] = 29'b0_001001001101_100_1_000100100110;
      patterns[4717] = 29'b0_001001001101_101_0_100010010011;
      patterns[4718] = 29'b0_001001001101_110_0_001001001101;
      patterns[4719] = 29'b0_001001001101_111_0_001001001101;
      patterns[4720] = 29'b0_001001001110_000_0_001001001110;
      patterns[4721] = 29'b0_001001001110_001_0_001110001001;
      patterns[4722] = 29'b0_001001001110_010_0_010010011100;
      patterns[4723] = 29'b0_001001001110_011_0_100100111000;
      patterns[4724] = 29'b0_001001001110_100_0_000100100111;
      patterns[4725] = 29'b0_001001001110_101_1_000010010011;
      patterns[4726] = 29'b0_001001001110_110_0_001001001110;
      patterns[4727] = 29'b0_001001001110_111_0_001001001110;
      patterns[4728] = 29'b0_001001001111_000_0_001001001111;
      patterns[4729] = 29'b0_001001001111_001_0_001111001001;
      patterns[4730] = 29'b0_001001001111_010_0_010010011110;
      patterns[4731] = 29'b0_001001001111_011_0_100100111100;
      patterns[4732] = 29'b0_001001001111_100_1_000100100111;
      patterns[4733] = 29'b0_001001001111_101_1_100010010011;
      patterns[4734] = 29'b0_001001001111_110_0_001001001111;
      patterns[4735] = 29'b0_001001001111_111_0_001001001111;
      patterns[4736] = 29'b0_001001010000_000_0_001001010000;
      patterns[4737] = 29'b0_001001010000_001_0_010000001001;
      patterns[4738] = 29'b0_001001010000_010_0_010010100000;
      patterns[4739] = 29'b0_001001010000_011_0_100101000000;
      patterns[4740] = 29'b0_001001010000_100_0_000100101000;
      patterns[4741] = 29'b0_001001010000_101_0_000010010100;
      patterns[4742] = 29'b0_001001010000_110_0_001001010000;
      patterns[4743] = 29'b0_001001010000_111_0_001001010000;
      patterns[4744] = 29'b0_001001010001_000_0_001001010001;
      patterns[4745] = 29'b0_001001010001_001_0_010001001001;
      patterns[4746] = 29'b0_001001010001_010_0_010010100010;
      patterns[4747] = 29'b0_001001010001_011_0_100101000100;
      patterns[4748] = 29'b0_001001010001_100_1_000100101000;
      patterns[4749] = 29'b0_001001010001_101_0_100010010100;
      patterns[4750] = 29'b0_001001010001_110_0_001001010001;
      patterns[4751] = 29'b0_001001010001_111_0_001001010001;
      patterns[4752] = 29'b0_001001010010_000_0_001001010010;
      patterns[4753] = 29'b0_001001010010_001_0_010010001001;
      patterns[4754] = 29'b0_001001010010_010_0_010010100100;
      patterns[4755] = 29'b0_001001010010_011_0_100101001000;
      patterns[4756] = 29'b0_001001010010_100_0_000100101001;
      patterns[4757] = 29'b0_001001010010_101_1_000010010100;
      patterns[4758] = 29'b0_001001010010_110_0_001001010010;
      patterns[4759] = 29'b0_001001010010_111_0_001001010010;
      patterns[4760] = 29'b0_001001010011_000_0_001001010011;
      patterns[4761] = 29'b0_001001010011_001_0_010011001001;
      patterns[4762] = 29'b0_001001010011_010_0_010010100110;
      patterns[4763] = 29'b0_001001010011_011_0_100101001100;
      patterns[4764] = 29'b0_001001010011_100_1_000100101001;
      patterns[4765] = 29'b0_001001010011_101_1_100010010100;
      patterns[4766] = 29'b0_001001010011_110_0_001001010011;
      patterns[4767] = 29'b0_001001010011_111_0_001001010011;
      patterns[4768] = 29'b0_001001010100_000_0_001001010100;
      patterns[4769] = 29'b0_001001010100_001_0_010100001001;
      patterns[4770] = 29'b0_001001010100_010_0_010010101000;
      patterns[4771] = 29'b0_001001010100_011_0_100101010000;
      patterns[4772] = 29'b0_001001010100_100_0_000100101010;
      patterns[4773] = 29'b0_001001010100_101_0_000010010101;
      patterns[4774] = 29'b0_001001010100_110_0_001001010100;
      patterns[4775] = 29'b0_001001010100_111_0_001001010100;
      patterns[4776] = 29'b0_001001010101_000_0_001001010101;
      patterns[4777] = 29'b0_001001010101_001_0_010101001001;
      patterns[4778] = 29'b0_001001010101_010_0_010010101010;
      patterns[4779] = 29'b0_001001010101_011_0_100101010100;
      patterns[4780] = 29'b0_001001010101_100_1_000100101010;
      patterns[4781] = 29'b0_001001010101_101_0_100010010101;
      patterns[4782] = 29'b0_001001010101_110_0_001001010101;
      patterns[4783] = 29'b0_001001010101_111_0_001001010101;
      patterns[4784] = 29'b0_001001010110_000_0_001001010110;
      patterns[4785] = 29'b0_001001010110_001_0_010110001001;
      patterns[4786] = 29'b0_001001010110_010_0_010010101100;
      patterns[4787] = 29'b0_001001010110_011_0_100101011000;
      patterns[4788] = 29'b0_001001010110_100_0_000100101011;
      patterns[4789] = 29'b0_001001010110_101_1_000010010101;
      patterns[4790] = 29'b0_001001010110_110_0_001001010110;
      patterns[4791] = 29'b0_001001010110_111_0_001001010110;
      patterns[4792] = 29'b0_001001010111_000_0_001001010111;
      patterns[4793] = 29'b0_001001010111_001_0_010111001001;
      patterns[4794] = 29'b0_001001010111_010_0_010010101110;
      patterns[4795] = 29'b0_001001010111_011_0_100101011100;
      patterns[4796] = 29'b0_001001010111_100_1_000100101011;
      patterns[4797] = 29'b0_001001010111_101_1_100010010101;
      patterns[4798] = 29'b0_001001010111_110_0_001001010111;
      patterns[4799] = 29'b0_001001010111_111_0_001001010111;
      patterns[4800] = 29'b0_001001011000_000_0_001001011000;
      patterns[4801] = 29'b0_001001011000_001_0_011000001001;
      patterns[4802] = 29'b0_001001011000_010_0_010010110000;
      patterns[4803] = 29'b0_001001011000_011_0_100101100000;
      patterns[4804] = 29'b0_001001011000_100_0_000100101100;
      patterns[4805] = 29'b0_001001011000_101_0_000010010110;
      patterns[4806] = 29'b0_001001011000_110_0_001001011000;
      patterns[4807] = 29'b0_001001011000_111_0_001001011000;
      patterns[4808] = 29'b0_001001011001_000_0_001001011001;
      patterns[4809] = 29'b0_001001011001_001_0_011001001001;
      patterns[4810] = 29'b0_001001011001_010_0_010010110010;
      patterns[4811] = 29'b0_001001011001_011_0_100101100100;
      patterns[4812] = 29'b0_001001011001_100_1_000100101100;
      patterns[4813] = 29'b0_001001011001_101_0_100010010110;
      patterns[4814] = 29'b0_001001011001_110_0_001001011001;
      patterns[4815] = 29'b0_001001011001_111_0_001001011001;
      patterns[4816] = 29'b0_001001011010_000_0_001001011010;
      patterns[4817] = 29'b0_001001011010_001_0_011010001001;
      patterns[4818] = 29'b0_001001011010_010_0_010010110100;
      patterns[4819] = 29'b0_001001011010_011_0_100101101000;
      patterns[4820] = 29'b0_001001011010_100_0_000100101101;
      patterns[4821] = 29'b0_001001011010_101_1_000010010110;
      patterns[4822] = 29'b0_001001011010_110_0_001001011010;
      patterns[4823] = 29'b0_001001011010_111_0_001001011010;
      patterns[4824] = 29'b0_001001011011_000_0_001001011011;
      patterns[4825] = 29'b0_001001011011_001_0_011011001001;
      patterns[4826] = 29'b0_001001011011_010_0_010010110110;
      patterns[4827] = 29'b0_001001011011_011_0_100101101100;
      patterns[4828] = 29'b0_001001011011_100_1_000100101101;
      patterns[4829] = 29'b0_001001011011_101_1_100010010110;
      patterns[4830] = 29'b0_001001011011_110_0_001001011011;
      patterns[4831] = 29'b0_001001011011_111_0_001001011011;
      patterns[4832] = 29'b0_001001011100_000_0_001001011100;
      patterns[4833] = 29'b0_001001011100_001_0_011100001001;
      patterns[4834] = 29'b0_001001011100_010_0_010010111000;
      patterns[4835] = 29'b0_001001011100_011_0_100101110000;
      patterns[4836] = 29'b0_001001011100_100_0_000100101110;
      patterns[4837] = 29'b0_001001011100_101_0_000010010111;
      patterns[4838] = 29'b0_001001011100_110_0_001001011100;
      patterns[4839] = 29'b0_001001011100_111_0_001001011100;
      patterns[4840] = 29'b0_001001011101_000_0_001001011101;
      patterns[4841] = 29'b0_001001011101_001_0_011101001001;
      patterns[4842] = 29'b0_001001011101_010_0_010010111010;
      patterns[4843] = 29'b0_001001011101_011_0_100101110100;
      patterns[4844] = 29'b0_001001011101_100_1_000100101110;
      patterns[4845] = 29'b0_001001011101_101_0_100010010111;
      patterns[4846] = 29'b0_001001011101_110_0_001001011101;
      patterns[4847] = 29'b0_001001011101_111_0_001001011101;
      patterns[4848] = 29'b0_001001011110_000_0_001001011110;
      patterns[4849] = 29'b0_001001011110_001_0_011110001001;
      patterns[4850] = 29'b0_001001011110_010_0_010010111100;
      patterns[4851] = 29'b0_001001011110_011_0_100101111000;
      patterns[4852] = 29'b0_001001011110_100_0_000100101111;
      patterns[4853] = 29'b0_001001011110_101_1_000010010111;
      patterns[4854] = 29'b0_001001011110_110_0_001001011110;
      patterns[4855] = 29'b0_001001011110_111_0_001001011110;
      patterns[4856] = 29'b0_001001011111_000_0_001001011111;
      patterns[4857] = 29'b0_001001011111_001_0_011111001001;
      patterns[4858] = 29'b0_001001011111_010_0_010010111110;
      patterns[4859] = 29'b0_001001011111_011_0_100101111100;
      patterns[4860] = 29'b0_001001011111_100_1_000100101111;
      patterns[4861] = 29'b0_001001011111_101_1_100010010111;
      patterns[4862] = 29'b0_001001011111_110_0_001001011111;
      patterns[4863] = 29'b0_001001011111_111_0_001001011111;
      patterns[4864] = 29'b0_001001100000_000_0_001001100000;
      patterns[4865] = 29'b0_001001100000_001_0_100000001001;
      patterns[4866] = 29'b0_001001100000_010_0_010011000000;
      patterns[4867] = 29'b0_001001100000_011_0_100110000000;
      patterns[4868] = 29'b0_001001100000_100_0_000100110000;
      patterns[4869] = 29'b0_001001100000_101_0_000010011000;
      patterns[4870] = 29'b0_001001100000_110_0_001001100000;
      patterns[4871] = 29'b0_001001100000_111_0_001001100000;
      patterns[4872] = 29'b0_001001100001_000_0_001001100001;
      patterns[4873] = 29'b0_001001100001_001_0_100001001001;
      patterns[4874] = 29'b0_001001100001_010_0_010011000010;
      patterns[4875] = 29'b0_001001100001_011_0_100110000100;
      patterns[4876] = 29'b0_001001100001_100_1_000100110000;
      patterns[4877] = 29'b0_001001100001_101_0_100010011000;
      patterns[4878] = 29'b0_001001100001_110_0_001001100001;
      patterns[4879] = 29'b0_001001100001_111_0_001001100001;
      patterns[4880] = 29'b0_001001100010_000_0_001001100010;
      patterns[4881] = 29'b0_001001100010_001_0_100010001001;
      patterns[4882] = 29'b0_001001100010_010_0_010011000100;
      patterns[4883] = 29'b0_001001100010_011_0_100110001000;
      patterns[4884] = 29'b0_001001100010_100_0_000100110001;
      patterns[4885] = 29'b0_001001100010_101_1_000010011000;
      patterns[4886] = 29'b0_001001100010_110_0_001001100010;
      patterns[4887] = 29'b0_001001100010_111_0_001001100010;
      patterns[4888] = 29'b0_001001100011_000_0_001001100011;
      patterns[4889] = 29'b0_001001100011_001_0_100011001001;
      patterns[4890] = 29'b0_001001100011_010_0_010011000110;
      patterns[4891] = 29'b0_001001100011_011_0_100110001100;
      patterns[4892] = 29'b0_001001100011_100_1_000100110001;
      patterns[4893] = 29'b0_001001100011_101_1_100010011000;
      patterns[4894] = 29'b0_001001100011_110_0_001001100011;
      patterns[4895] = 29'b0_001001100011_111_0_001001100011;
      patterns[4896] = 29'b0_001001100100_000_0_001001100100;
      patterns[4897] = 29'b0_001001100100_001_0_100100001001;
      patterns[4898] = 29'b0_001001100100_010_0_010011001000;
      patterns[4899] = 29'b0_001001100100_011_0_100110010000;
      patterns[4900] = 29'b0_001001100100_100_0_000100110010;
      patterns[4901] = 29'b0_001001100100_101_0_000010011001;
      patterns[4902] = 29'b0_001001100100_110_0_001001100100;
      patterns[4903] = 29'b0_001001100100_111_0_001001100100;
      patterns[4904] = 29'b0_001001100101_000_0_001001100101;
      patterns[4905] = 29'b0_001001100101_001_0_100101001001;
      patterns[4906] = 29'b0_001001100101_010_0_010011001010;
      patterns[4907] = 29'b0_001001100101_011_0_100110010100;
      patterns[4908] = 29'b0_001001100101_100_1_000100110010;
      patterns[4909] = 29'b0_001001100101_101_0_100010011001;
      patterns[4910] = 29'b0_001001100101_110_0_001001100101;
      patterns[4911] = 29'b0_001001100101_111_0_001001100101;
      patterns[4912] = 29'b0_001001100110_000_0_001001100110;
      patterns[4913] = 29'b0_001001100110_001_0_100110001001;
      patterns[4914] = 29'b0_001001100110_010_0_010011001100;
      patterns[4915] = 29'b0_001001100110_011_0_100110011000;
      patterns[4916] = 29'b0_001001100110_100_0_000100110011;
      patterns[4917] = 29'b0_001001100110_101_1_000010011001;
      patterns[4918] = 29'b0_001001100110_110_0_001001100110;
      patterns[4919] = 29'b0_001001100110_111_0_001001100110;
      patterns[4920] = 29'b0_001001100111_000_0_001001100111;
      patterns[4921] = 29'b0_001001100111_001_0_100111001001;
      patterns[4922] = 29'b0_001001100111_010_0_010011001110;
      patterns[4923] = 29'b0_001001100111_011_0_100110011100;
      patterns[4924] = 29'b0_001001100111_100_1_000100110011;
      patterns[4925] = 29'b0_001001100111_101_1_100010011001;
      patterns[4926] = 29'b0_001001100111_110_0_001001100111;
      patterns[4927] = 29'b0_001001100111_111_0_001001100111;
      patterns[4928] = 29'b0_001001101000_000_0_001001101000;
      patterns[4929] = 29'b0_001001101000_001_0_101000001001;
      patterns[4930] = 29'b0_001001101000_010_0_010011010000;
      patterns[4931] = 29'b0_001001101000_011_0_100110100000;
      patterns[4932] = 29'b0_001001101000_100_0_000100110100;
      patterns[4933] = 29'b0_001001101000_101_0_000010011010;
      patterns[4934] = 29'b0_001001101000_110_0_001001101000;
      patterns[4935] = 29'b0_001001101000_111_0_001001101000;
      patterns[4936] = 29'b0_001001101001_000_0_001001101001;
      patterns[4937] = 29'b0_001001101001_001_0_101001001001;
      patterns[4938] = 29'b0_001001101001_010_0_010011010010;
      patterns[4939] = 29'b0_001001101001_011_0_100110100100;
      patterns[4940] = 29'b0_001001101001_100_1_000100110100;
      patterns[4941] = 29'b0_001001101001_101_0_100010011010;
      patterns[4942] = 29'b0_001001101001_110_0_001001101001;
      patterns[4943] = 29'b0_001001101001_111_0_001001101001;
      patterns[4944] = 29'b0_001001101010_000_0_001001101010;
      patterns[4945] = 29'b0_001001101010_001_0_101010001001;
      patterns[4946] = 29'b0_001001101010_010_0_010011010100;
      patterns[4947] = 29'b0_001001101010_011_0_100110101000;
      patterns[4948] = 29'b0_001001101010_100_0_000100110101;
      patterns[4949] = 29'b0_001001101010_101_1_000010011010;
      patterns[4950] = 29'b0_001001101010_110_0_001001101010;
      patterns[4951] = 29'b0_001001101010_111_0_001001101010;
      patterns[4952] = 29'b0_001001101011_000_0_001001101011;
      patterns[4953] = 29'b0_001001101011_001_0_101011001001;
      patterns[4954] = 29'b0_001001101011_010_0_010011010110;
      patterns[4955] = 29'b0_001001101011_011_0_100110101100;
      patterns[4956] = 29'b0_001001101011_100_1_000100110101;
      patterns[4957] = 29'b0_001001101011_101_1_100010011010;
      patterns[4958] = 29'b0_001001101011_110_0_001001101011;
      patterns[4959] = 29'b0_001001101011_111_0_001001101011;
      patterns[4960] = 29'b0_001001101100_000_0_001001101100;
      patterns[4961] = 29'b0_001001101100_001_0_101100001001;
      patterns[4962] = 29'b0_001001101100_010_0_010011011000;
      patterns[4963] = 29'b0_001001101100_011_0_100110110000;
      patterns[4964] = 29'b0_001001101100_100_0_000100110110;
      patterns[4965] = 29'b0_001001101100_101_0_000010011011;
      patterns[4966] = 29'b0_001001101100_110_0_001001101100;
      patterns[4967] = 29'b0_001001101100_111_0_001001101100;
      patterns[4968] = 29'b0_001001101101_000_0_001001101101;
      patterns[4969] = 29'b0_001001101101_001_0_101101001001;
      patterns[4970] = 29'b0_001001101101_010_0_010011011010;
      patterns[4971] = 29'b0_001001101101_011_0_100110110100;
      patterns[4972] = 29'b0_001001101101_100_1_000100110110;
      patterns[4973] = 29'b0_001001101101_101_0_100010011011;
      patterns[4974] = 29'b0_001001101101_110_0_001001101101;
      patterns[4975] = 29'b0_001001101101_111_0_001001101101;
      patterns[4976] = 29'b0_001001101110_000_0_001001101110;
      patterns[4977] = 29'b0_001001101110_001_0_101110001001;
      patterns[4978] = 29'b0_001001101110_010_0_010011011100;
      patterns[4979] = 29'b0_001001101110_011_0_100110111000;
      patterns[4980] = 29'b0_001001101110_100_0_000100110111;
      patterns[4981] = 29'b0_001001101110_101_1_000010011011;
      patterns[4982] = 29'b0_001001101110_110_0_001001101110;
      patterns[4983] = 29'b0_001001101110_111_0_001001101110;
      patterns[4984] = 29'b0_001001101111_000_0_001001101111;
      patterns[4985] = 29'b0_001001101111_001_0_101111001001;
      patterns[4986] = 29'b0_001001101111_010_0_010011011110;
      patterns[4987] = 29'b0_001001101111_011_0_100110111100;
      patterns[4988] = 29'b0_001001101111_100_1_000100110111;
      patterns[4989] = 29'b0_001001101111_101_1_100010011011;
      patterns[4990] = 29'b0_001001101111_110_0_001001101111;
      patterns[4991] = 29'b0_001001101111_111_0_001001101111;
      patterns[4992] = 29'b0_001001110000_000_0_001001110000;
      patterns[4993] = 29'b0_001001110000_001_0_110000001001;
      patterns[4994] = 29'b0_001001110000_010_0_010011100000;
      patterns[4995] = 29'b0_001001110000_011_0_100111000000;
      patterns[4996] = 29'b0_001001110000_100_0_000100111000;
      patterns[4997] = 29'b0_001001110000_101_0_000010011100;
      patterns[4998] = 29'b0_001001110000_110_0_001001110000;
      patterns[4999] = 29'b0_001001110000_111_0_001001110000;
      patterns[5000] = 29'b0_001001110001_000_0_001001110001;
      patterns[5001] = 29'b0_001001110001_001_0_110001001001;
      patterns[5002] = 29'b0_001001110001_010_0_010011100010;
      patterns[5003] = 29'b0_001001110001_011_0_100111000100;
      patterns[5004] = 29'b0_001001110001_100_1_000100111000;
      patterns[5005] = 29'b0_001001110001_101_0_100010011100;
      patterns[5006] = 29'b0_001001110001_110_0_001001110001;
      patterns[5007] = 29'b0_001001110001_111_0_001001110001;
      patterns[5008] = 29'b0_001001110010_000_0_001001110010;
      patterns[5009] = 29'b0_001001110010_001_0_110010001001;
      patterns[5010] = 29'b0_001001110010_010_0_010011100100;
      patterns[5011] = 29'b0_001001110010_011_0_100111001000;
      patterns[5012] = 29'b0_001001110010_100_0_000100111001;
      patterns[5013] = 29'b0_001001110010_101_1_000010011100;
      patterns[5014] = 29'b0_001001110010_110_0_001001110010;
      patterns[5015] = 29'b0_001001110010_111_0_001001110010;
      patterns[5016] = 29'b0_001001110011_000_0_001001110011;
      patterns[5017] = 29'b0_001001110011_001_0_110011001001;
      patterns[5018] = 29'b0_001001110011_010_0_010011100110;
      patterns[5019] = 29'b0_001001110011_011_0_100111001100;
      patterns[5020] = 29'b0_001001110011_100_1_000100111001;
      patterns[5021] = 29'b0_001001110011_101_1_100010011100;
      patterns[5022] = 29'b0_001001110011_110_0_001001110011;
      patterns[5023] = 29'b0_001001110011_111_0_001001110011;
      patterns[5024] = 29'b0_001001110100_000_0_001001110100;
      patterns[5025] = 29'b0_001001110100_001_0_110100001001;
      patterns[5026] = 29'b0_001001110100_010_0_010011101000;
      patterns[5027] = 29'b0_001001110100_011_0_100111010000;
      patterns[5028] = 29'b0_001001110100_100_0_000100111010;
      patterns[5029] = 29'b0_001001110100_101_0_000010011101;
      patterns[5030] = 29'b0_001001110100_110_0_001001110100;
      patterns[5031] = 29'b0_001001110100_111_0_001001110100;
      patterns[5032] = 29'b0_001001110101_000_0_001001110101;
      patterns[5033] = 29'b0_001001110101_001_0_110101001001;
      patterns[5034] = 29'b0_001001110101_010_0_010011101010;
      patterns[5035] = 29'b0_001001110101_011_0_100111010100;
      patterns[5036] = 29'b0_001001110101_100_1_000100111010;
      patterns[5037] = 29'b0_001001110101_101_0_100010011101;
      patterns[5038] = 29'b0_001001110101_110_0_001001110101;
      patterns[5039] = 29'b0_001001110101_111_0_001001110101;
      patterns[5040] = 29'b0_001001110110_000_0_001001110110;
      patterns[5041] = 29'b0_001001110110_001_0_110110001001;
      patterns[5042] = 29'b0_001001110110_010_0_010011101100;
      patterns[5043] = 29'b0_001001110110_011_0_100111011000;
      patterns[5044] = 29'b0_001001110110_100_0_000100111011;
      patterns[5045] = 29'b0_001001110110_101_1_000010011101;
      patterns[5046] = 29'b0_001001110110_110_0_001001110110;
      patterns[5047] = 29'b0_001001110110_111_0_001001110110;
      patterns[5048] = 29'b0_001001110111_000_0_001001110111;
      patterns[5049] = 29'b0_001001110111_001_0_110111001001;
      patterns[5050] = 29'b0_001001110111_010_0_010011101110;
      patterns[5051] = 29'b0_001001110111_011_0_100111011100;
      patterns[5052] = 29'b0_001001110111_100_1_000100111011;
      patterns[5053] = 29'b0_001001110111_101_1_100010011101;
      patterns[5054] = 29'b0_001001110111_110_0_001001110111;
      patterns[5055] = 29'b0_001001110111_111_0_001001110111;
      patterns[5056] = 29'b0_001001111000_000_0_001001111000;
      patterns[5057] = 29'b0_001001111000_001_0_111000001001;
      patterns[5058] = 29'b0_001001111000_010_0_010011110000;
      patterns[5059] = 29'b0_001001111000_011_0_100111100000;
      patterns[5060] = 29'b0_001001111000_100_0_000100111100;
      patterns[5061] = 29'b0_001001111000_101_0_000010011110;
      patterns[5062] = 29'b0_001001111000_110_0_001001111000;
      patterns[5063] = 29'b0_001001111000_111_0_001001111000;
      patterns[5064] = 29'b0_001001111001_000_0_001001111001;
      patterns[5065] = 29'b0_001001111001_001_0_111001001001;
      patterns[5066] = 29'b0_001001111001_010_0_010011110010;
      patterns[5067] = 29'b0_001001111001_011_0_100111100100;
      patterns[5068] = 29'b0_001001111001_100_1_000100111100;
      patterns[5069] = 29'b0_001001111001_101_0_100010011110;
      patterns[5070] = 29'b0_001001111001_110_0_001001111001;
      patterns[5071] = 29'b0_001001111001_111_0_001001111001;
      patterns[5072] = 29'b0_001001111010_000_0_001001111010;
      patterns[5073] = 29'b0_001001111010_001_0_111010001001;
      patterns[5074] = 29'b0_001001111010_010_0_010011110100;
      patterns[5075] = 29'b0_001001111010_011_0_100111101000;
      patterns[5076] = 29'b0_001001111010_100_0_000100111101;
      patterns[5077] = 29'b0_001001111010_101_1_000010011110;
      patterns[5078] = 29'b0_001001111010_110_0_001001111010;
      patterns[5079] = 29'b0_001001111010_111_0_001001111010;
      patterns[5080] = 29'b0_001001111011_000_0_001001111011;
      patterns[5081] = 29'b0_001001111011_001_0_111011001001;
      patterns[5082] = 29'b0_001001111011_010_0_010011110110;
      patterns[5083] = 29'b0_001001111011_011_0_100111101100;
      patterns[5084] = 29'b0_001001111011_100_1_000100111101;
      patterns[5085] = 29'b0_001001111011_101_1_100010011110;
      patterns[5086] = 29'b0_001001111011_110_0_001001111011;
      patterns[5087] = 29'b0_001001111011_111_0_001001111011;
      patterns[5088] = 29'b0_001001111100_000_0_001001111100;
      patterns[5089] = 29'b0_001001111100_001_0_111100001001;
      patterns[5090] = 29'b0_001001111100_010_0_010011111000;
      patterns[5091] = 29'b0_001001111100_011_0_100111110000;
      patterns[5092] = 29'b0_001001111100_100_0_000100111110;
      patterns[5093] = 29'b0_001001111100_101_0_000010011111;
      patterns[5094] = 29'b0_001001111100_110_0_001001111100;
      patterns[5095] = 29'b0_001001111100_111_0_001001111100;
      patterns[5096] = 29'b0_001001111101_000_0_001001111101;
      patterns[5097] = 29'b0_001001111101_001_0_111101001001;
      patterns[5098] = 29'b0_001001111101_010_0_010011111010;
      patterns[5099] = 29'b0_001001111101_011_0_100111110100;
      patterns[5100] = 29'b0_001001111101_100_1_000100111110;
      patterns[5101] = 29'b0_001001111101_101_0_100010011111;
      patterns[5102] = 29'b0_001001111101_110_0_001001111101;
      patterns[5103] = 29'b0_001001111101_111_0_001001111101;
      patterns[5104] = 29'b0_001001111110_000_0_001001111110;
      patterns[5105] = 29'b0_001001111110_001_0_111110001001;
      patterns[5106] = 29'b0_001001111110_010_0_010011111100;
      patterns[5107] = 29'b0_001001111110_011_0_100111111000;
      patterns[5108] = 29'b0_001001111110_100_0_000100111111;
      patterns[5109] = 29'b0_001001111110_101_1_000010011111;
      patterns[5110] = 29'b0_001001111110_110_0_001001111110;
      patterns[5111] = 29'b0_001001111110_111_0_001001111110;
      patterns[5112] = 29'b0_001001111111_000_0_001001111111;
      patterns[5113] = 29'b0_001001111111_001_0_111111001001;
      patterns[5114] = 29'b0_001001111111_010_0_010011111110;
      patterns[5115] = 29'b0_001001111111_011_0_100111111100;
      patterns[5116] = 29'b0_001001111111_100_1_000100111111;
      patterns[5117] = 29'b0_001001111111_101_1_100010011111;
      patterns[5118] = 29'b0_001001111111_110_0_001001111111;
      patterns[5119] = 29'b0_001001111111_111_0_001001111111;
      patterns[5120] = 29'b0_001010000000_000_0_001010000000;
      patterns[5121] = 29'b0_001010000000_001_0_000000001010;
      patterns[5122] = 29'b0_001010000000_010_0_010100000000;
      patterns[5123] = 29'b0_001010000000_011_0_101000000000;
      patterns[5124] = 29'b0_001010000000_100_0_000101000000;
      patterns[5125] = 29'b0_001010000000_101_0_000010100000;
      patterns[5126] = 29'b0_001010000000_110_0_001010000000;
      patterns[5127] = 29'b0_001010000000_111_0_001010000000;
      patterns[5128] = 29'b0_001010000001_000_0_001010000001;
      patterns[5129] = 29'b0_001010000001_001_0_000001001010;
      patterns[5130] = 29'b0_001010000001_010_0_010100000010;
      patterns[5131] = 29'b0_001010000001_011_0_101000000100;
      patterns[5132] = 29'b0_001010000001_100_1_000101000000;
      patterns[5133] = 29'b0_001010000001_101_0_100010100000;
      patterns[5134] = 29'b0_001010000001_110_0_001010000001;
      patterns[5135] = 29'b0_001010000001_111_0_001010000001;
      patterns[5136] = 29'b0_001010000010_000_0_001010000010;
      patterns[5137] = 29'b0_001010000010_001_0_000010001010;
      patterns[5138] = 29'b0_001010000010_010_0_010100000100;
      patterns[5139] = 29'b0_001010000010_011_0_101000001000;
      patterns[5140] = 29'b0_001010000010_100_0_000101000001;
      patterns[5141] = 29'b0_001010000010_101_1_000010100000;
      patterns[5142] = 29'b0_001010000010_110_0_001010000010;
      patterns[5143] = 29'b0_001010000010_111_0_001010000010;
      patterns[5144] = 29'b0_001010000011_000_0_001010000011;
      patterns[5145] = 29'b0_001010000011_001_0_000011001010;
      patterns[5146] = 29'b0_001010000011_010_0_010100000110;
      patterns[5147] = 29'b0_001010000011_011_0_101000001100;
      patterns[5148] = 29'b0_001010000011_100_1_000101000001;
      patterns[5149] = 29'b0_001010000011_101_1_100010100000;
      patterns[5150] = 29'b0_001010000011_110_0_001010000011;
      patterns[5151] = 29'b0_001010000011_111_0_001010000011;
      patterns[5152] = 29'b0_001010000100_000_0_001010000100;
      patterns[5153] = 29'b0_001010000100_001_0_000100001010;
      patterns[5154] = 29'b0_001010000100_010_0_010100001000;
      patterns[5155] = 29'b0_001010000100_011_0_101000010000;
      patterns[5156] = 29'b0_001010000100_100_0_000101000010;
      patterns[5157] = 29'b0_001010000100_101_0_000010100001;
      patterns[5158] = 29'b0_001010000100_110_0_001010000100;
      patterns[5159] = 29'b0_001010000100_111_0_001010000100;
      patterns[5160] = 29'b0_001010000101_000_0_001010000101;
      patterns[5161] = 29'b0_001010000101_001_0_000101001010;
      patterns[5162] = 29'b0_001010000101_010_0_010100001010;
      patterns[5163] = 29'b0_001010000101_011_0_101000010100;
      patterns[5164] = 29'b0_001010000101_100_1_000101000010;
      patterns[5165] = 29'b0_001010000101_101_0_100010100001;
      patterns[5166] = 29'b0_001010000101_110_0_001010000101;
      patterns[5167] = 29'b0_001010000101_111_0_001010000101;
      patterns[5168] = 29'b0_001010000110_000_0_001010000110;
      patterns[5169] = 29'b0_001010000110_001_0_000110001010;
      patterns[5170] = 29'b0_001010000110_010_0_010100001100;
      patterns[5171] = 29'b0_001010000110_011_0_101000011000;
      patterns[5172] = 29'b0_001010000110_100_0_000101000011;
      patterns[5173] = 29'b0_001010000110_101_1_000010100001;
      patterns[5174] = 29'b0_001010000110_110_0_001010000110;
      patterns[5175] = 29'b0_001010000110_111_0_001010000110;
      patterns[5176] = 29'b0_001010000111_000_0_001010000111;
      patterns[5177] = 29'b0_001010000111_001_0_000111001010;
      patterns[5178] = 29'b0_001010000111_010_0_010100001110;
      patterns[5179] = 29'b0_001010000111_011_0_101000011100;
      patterns[5180] = 29'b0_001010000111_100_1_000101000011;
      patterns[5181] = 29'b0_001010000111_101_1_100010100001;
      patterns[5182] = 29'b0_001010000111_110_0_001010000111;
      patterns[5183] = 29'b0_001010000111_111_0_001010000111;
      patterns[5184] = 29'b0_001010001000_000_0_001010001000;
      patterns[5185] = 29'b0_001010001000_001_0_001000001010;
      patterns[5186] = 29'b0_001010001000_010_0_010100010000;
      patterns[5187] = 29'b0_001010001000_011_0_101000100000;
      patterns[5188] = 29'b0_001010001000_100_0_000101000100;
      patterns[5189] = 29'b0_001010001000_101_0_000010100010;
      patterns[5190] = 29'b0_001010001000_110_0_001010001000;
      patterns[5191] = 29'b0_001010001000_111_0_001010001000;
      patterns[5192] = 29'b0_001010001001_000_0_001010001001;
      patterns[5193] = 29'b0_001010001001_001_0_001001001010;
      patterns[5194] = 29'b0_001010001001_010_0_010100010010;
      patterns[5195] = 29'b0_001010001001_011_0_101000100100;
      patterns[5196] = 29'b0_001010001001_100_1_000101000100;
      patterns[5197] = 29'b0_001010001001_101_0_100010100010;
      patterns[5198] = 29'b0_001010001001_110_0_001010001001;
      patterns[5199] = 29'b0_001010001001_111_0_001010001001;
      patterns[5200] = 29'b0_001010001010_000_0_001010001010;
      patterns[5201] = 29'b0_001010001010_001_0_001010001010;
      patterns[5202] = 29'b0_001010001010_010_0_010100010100;
      patterns[5203] = 29'b0_001010001010_011_0_101000101000;
      patterns[5204] = 29'b0_001010001010_100_0_000101000101;
      patterns[5205] = 29'b0_001010001010_101_1_000010100010;
      patterns[5206] = 29'b0_001010001010_110_0_001010001010;
      patterns[5207] = 29'b0_001010001010_111_0_001010001010;
      patterns[5208] = 29'b0_001010001011_000_0_001010001011;
      patterns[5209] = 29'b0_001010001011_001_0_001011001010;
      patterns[5210] = 29'b0_001010001011_010_0_010100010110;
      patterns[5211] = 29'b0_001010001011_011_0_101000101100;
      patterns[5212] = 29'b0_001010001011_100_1_000101000101;
      patterns[5213] = 29'b0_001010001011_101_1_100010100010;
      patterns[5214] = 29'b0_001010001011_110_0_001010001011;
      patterns[5215] = 29'b0_001010001011_111_0_001010001011;
      patterns[5216] = 29'b0_001010001100_000_0_001010001100;
      patterns[5217] = 29'b0_001010001100_001_0_001100001010;
      patterns[5218] = 29'b0_001010001100_010_0_010100011000;
      patterns[5219] = 29'b0_001010001100_011_0_101000110000;
      patterns[5220] = 29'b0_001010001100_100_0_000101000110;
      patterns[5221] = 29'b0_001010001100_101_0_000010100011;
      patterns[5222] = 29'b0_001010001100_110_0_001010001100;
      patterns[5223] = 29'b0_001010001100_111_0_001010001100;
      patterns[5224] = 29'b0_001010001101_000_0_001010001101;
      patterns[5225] = 29'b0_001010001101_001_0_001101001010;
      patterns[5226] = 29'b0_001010001101_010_0_010100011010;
      patterns[5227] = 29'b0_001010001101_011_0_101000110100;
      patterns[5228] = 29'b0_001010001101_100_1_000101000110;
      patterns[5229] = 29'b0_001010001101_101_0_100010100011;
      patterns[5230] = 29'b0_001010001101_110_0_001010001101;
      patterns[5231] = 29'b0_001010001101_111_0_001010001101;
      patterns[5232] = 29'b0_001010001110_000_0_001010001110;
      patterns[5233] = 29'b0_001010001110_001_0_001110001010;
      patterns[5234] = 29'b0_001010001110_010_0_010100011100;
      patterns[5235] = 29'b0_001010001110_011_0_101000111000;
      patterns[5236] = 29'b0_001010001110_100_0_000101000111;
      patterns[5237] = 29'b0_001010001110_101_1_000010100011;
      patterns[5238] = 29'b0_001010001110_110_0_001010001110;
      patterns[5239] = 29'b0_001010001110_111_0_001010001110;
      patterns[5240] = 29'b0_001010001111_000_0_001010001111;
      patterns[5241] = 29'b0_001010001111_001_0_001111001010;
      patterns[5242] = 29'b0_001010001111_010_0_010100011110;
      patterns[5243] = 29'b0_001010001111_011_0_101000111100;
      patterns[5244] = 29'b0_001010001111_100_1_000101000111;
      patterns[5245] = 29'b0_001010001111_101_1_100010100011;
      patterns[5246] = 29'b0_001010001111_110_0_001010001111;
      patterns[5247] = 29'b0_001010001111_111_0_001010001111;
      patterns[5248] = 29'b0_001010010000_000_0_001010010000;
      patterns[5249] = 29'b0_001010010000_001_0_010000001010;
      patterns[5250] = 29'b0_001010010000_010_0_010100100000;
      patterns[5251] = 29'b0_001010010000_011_0_101001000000;
      patterns[5252] = 29'b0_001010010000_100_0_000101001000;
      patterns[5253] = 29'b0_001010010000_101_0_000010100100;
      patterns[5254] = 29'b0_001010010000_110_0_001010010000;
      patterns[5255] = 29'b0_001010010000_111_0_001010010000;
      patterns[5256] = 29'b0_001010010001_000_0_001010010001;
      patterns[5257] = 29'b0_001010010001_001_0_010001001010;
      patterns[5258] = 29'b0_001010010001_010_0_010100100010;
      patterns[5259] = 29'b0_001010010001_011_0_101001000100;
      patterns[5260] = 29'b0_001010010001_100_1_000101001000;
      patterns[5261] = 29'b0_001010010001_101_0_100010100100;
      patterns[5262] = 29'b0_001010010001_110_0_001010010001;
      patterns[5263] = 29'b0_001010010001_111_0_001010010001;
      patterns[5264] = 29'b0_001010010010_000_0_001010010010;
      patterns[5265] = 29'b0_001010010010_001_0_010010001010;
      patterns[5266] = 29'b0_001010010010_010_0_010100100100;
      patterns[5267] = 29'b0_001010010010_011_0_101001001000;
      patterns[5268] = 29'b0_001010010010_100_0_000101001001;
      patterns[5269] = 29'b0_001010010010_101_1_000010100100;
      patterns[5270] = 29'b0_001010010010_110_0_001010010010;
      patterns[5271] = 29'b0_001010010010_111_0_001010010010;
      patterns[5272] = 29'b0_001010010011_000_0_001010010011;
      patterns[5273] = 29'b0_001010010011_001_0_010011001010;
      patterns[5274] = 29'b0_001010010011_010_0_010100100110;
      patterns[5275] = 29'b0_001010010011_011_0_101001001100;
      patterns[5276] = 29'b0_001010010011_100_1_000101001001;
      patterns[5277] = 29'b0_001010010011_101_1_100010100100;
      patterns[5278] = 29'b0_001010010011_110_0_001010010011;
      patterns[5279] = 29'b0_001010010011_111_0_001010010011;
      patterns[5280] = 29'b0_001010010100_000_0_001010010100;
      patterns[5281] = 29'b0_001010010100_001_0_010100001010;
      patterns[5282] = 29'b0_001010010100_010_0_010100101000;
      patterns[5283] = 29'b0_001010010100_011_0_101001010000;
      patterns[5284] = 29'b0_001010010100_100_0_000101001010;
      patterns[5285] = 29'b0_001010010100_101_0_000010100101;
      patterns[5286] = 29'b0_001010010100_110_0_001010010100;
      patterns[5287] = 29'b0_001010010100_111_0_001010010100;
      patterns[5288] = 29'b0_001010010101_000_0_001010010101;
      patterns[5289] = 29'b0_001010010101_001_0_010101001010;
      patterns[5290] = 29'b0_001010010101_010_0_010100101010;
      patterns[5291] = 29'b0_001010010101_011_0_101001010100;
      patterns[5292] = 29'b0_001010010101_100_1_000101001010;
      patterns[5293] = 29'b0_001010010101_101_0_100010100101;
      patterns[5294] = 29'b0_001010010101_110_0_001010010101;
      patterns[5295] = 29'b0_001010010101_111_0_001010010101;
      patterns[5296] = 29'b0_001010010110_000_0_001010010110;
      patterns[5297] = 29'b0_001010010110_001_0_010110001010;
      patterns[5298] = 29'b0_001010010110_010_0_010100101100;
      patterns[5299] = 29'b0_001010010110_011_0_101001011000;
      patterns[5300] = 29'b0_001010010110_100_0_000101001011;
      patterns[5301] = 29'b0_001010010110_101_1_000010100101;
      patterns[5302] = 29'b0_001010010110_110_0_001010010110;
      patterns[5303] = 29'b0_001010010110_111_0_001010010110;
      patterns[5304] = 29'b0_001010010111_000_0_001010010111;
      patterns[5305] = 29'b0_001010010111_001_0_010111001010;
      patterns[5306] = 29'b0_001010010111_010_0_010100101110;
      patterns[5307] = 29'b0_001010010111_011_0_101001011100;
      patterns[5308] = 29'b0_001010010111_100_1_000101001011;
      patterns[5309] = 29'b0_001010010111_101_1_100010100101;
      patterns[5310] = 29'b0_001010010111_110_0_001010010111;
      patterns[5311] = 29'b0_001010010111_111_0_001010010111;
      patterns[5312] = 29'b0_001010011000_000_0_001010011000;
      patterns[5313] = 29'b0_001010011000_001_0_011000001010;
      patterns[5314] = 29'b0_001010011000_010_0_010100110000;
      patterns[5315] = 29'b0_001010011000_011_0_101001100000;
      patterns[5316] = 29'b0_001010011000_100_0_000101001100;
      patterns[5317] = 29'b0_001010011000_101_0_000010100110;
      patterns[5318] = 29'b0_001010011000_110_0_001010011000;
      patterns[5319] = 29'b0_001010011000_111_0_001010011000;
      patterns[5320] = 29'b0_001010011001_000_0_001010011001;
      patterns[5321] = 29'b0_001010011001_001_0_011001001010;
      patterns[5322] = 29'b0_001010011001_010_0_010100110010;
      patterns[5323] = 29'b0_001010011001_011_0_101001100100;
      patterns[5324] = 29'b0_001010011001_100_1_000101001100;
      patterns[5325] = 29'b0_001010011001_101_0_100010100110;
      patterns[5326] = 29'b0_001010011001_110_0_001010011001;
      patterns[5327] = 29'b0_001010011001_111_0_001010011001;
      patterns[5328] = 29'b0_001010011010_000_0_001010011010;
      patterns[5329] = 29'b0_001010011010_001_0_011010001010;
      patterns[5330] = 29'b0_001010011010_010_0_010100110100;
      patterns[5331] = 29'b0_001010011010_011_0_101001101000;
      patterns[5332] = 29'b0_001010011010_100_0_000101001101;
      patterns[5333] = 29'b0_001010011010_101_1_000010100110;
      patterns[5334] = 29'b0_001010011010_110_0_001010011010;
      patterns[5335] = 29'b0_001010011010_111_0_001010011010;
      patterns[5336] = 29'b0_001010011011_000_0_001010011011;
      patterns[5337] = 29'b0_001010011011_001_0_011011001010;
      patterns[5338] = 29'b0_001010011011_010_0_010100110110;
      patterns[5339] = 29'b0_001010011011_011_0_101001101100;
      patterns[5340] = 29'b0_001010011011_100_1_000101001101;
      patterns[5341] = 29'b0_001010011011_101_1_100010100110;
      patterns[5342] = 29'b0_001010011011_110_0_001010011011;
      patterns[5343] = 29'b0_001010011011_111_0_001010011011;
      patterns[5344] = 29'b0_001010011100_000_0_001010011100;
      patterns[5345] = 29'b0_001010011100_001_0_011100001010;
      patterns[5346] = 29'b0_001010011100_010_0_010100111000;
      patterns[5347] = 29'b0_001010011100_011_0_101001110000;
      patterns[5348] = 29'b0_001010011100_100_0_000101001110;
      patterns[5349] = 29'b0_001010011100_101_0_000010100111;
      patterns[5350] = 29'b0_001010011100_110_0_001010011100;
      patterns[5351] = 29'b0_001010011100_111_0_001010011100;
      patterns[5352] = 29'b0_001010011101_000_0_001010011101;
      patterns[5353] = 29'b0_001010011101_001_0_011101001010;
      patterns[5354] = 29'b0_001010011101_010_0_010100111010;
      patterns[5355] = 29'b0_001010011101_011_0_101001110100;
      patterns[5356] = 29'b0_001010011101_100_1_000101001110;
      patterns[5357] = 29'b0_001010011101_101_0_100010100111;
      patterns[5358] = 29'b0_001010011101_110_0_001010011101;
      patterns[5359] = 29'b0_001010011101_111_0_001010011101;
      patterns[5360] = 29'b0_001010011110_000_0_001010011110;
      patterns[5361] = 29'b0_001010011110_001_0_011110001010;
      patterns[5362] = 29'b0_001010011110_010_0_010100111100;
      patterns[5363] = 29'b0_001010011110_011_0_101001111000;
      patterns[5364] = 29'b0_001010011110_100_0_000101001111;
      patterns[5365] = 29'b0_001010011110_101_1_000010100111;
      patterns[5366] = 29'b0_001010011110_110_0_001010011110;
      patterns[5367] = 29'b0_001010011110_111_0_001010011110;
      patterns[5368] = 29'b0_001010011111_000_0_001010011111;
      patterns[5369] = 29'b0_001010011111_001_0_011111001010;
      patterns[5370] = 29'b0_001010011111_010_0_010100111110;
      patterns[5371] = 29'b0_001010011111_011_0_101001111100;
      patterns[5372] = 29'b0_001010011111_100_1_000101001111;
      patterns[5373] = 29'b0_001010011111_101_1_100010100111;
      patterns[5374] = 29'b0_001010011111_110_0_001010011111;
      patterns[5375] = 29'b0_001010011111_111_0_001010011111;
      patterns[5376] = 29'b0_001010100000_000_0_001010100000;
      patterns[5377] = 29'b0_001010100000_001_0_100000001010;
      patterns[5378] = 29'b0_001010100000_010_0_010101000000;
      patterns[5379] = 29'b0_001010100000_011_0_101010000000;
      patterns[5380] = 29'b0_001010100000_100_0_000101010000;
      patterns[5381] = 29'b0_001010100000_101_0_000010101000;
      patterns[5382] = 29'b0_001010100000_110_0_001010100000;
      patterns[5383] = 29'b0_001010100000_111_0_001010100000;
      patterns[5384] = 29'b0_001010100001_000_0_001010100001;
      patterns[5385] = 29'b0_001010100001_001_0_100001001010;
      patterns[5386] = 29'b0_001010100001_010_0_010101000010;
      patterns[5387] = 29'b0_001010100001_011_0_101010000100;
      patterns[5388] = 29'b0_001010100001_100_1_000101010000;
      patterns[5389] = 29'b0_001010100001_101_0_100010101000;
      patterns[5390] = 29'b0_001010100001_110_0_001010100001;
      patterns[5391] = 29'b0_001010100001_111_0_001010100001;
      patterns[5392] = 29'b0_001010100010_000_0_001010100010;
      patterns[5393] = 29'b0_001010100010_001_0_100010001010;
      patterns[5394] = 29'b0_001010100010_010_0_010101000100;
      patterns[5395] = 29'b0_001010100010_011_0_101010001000;
      patterns[5396] = 29'b0_001010100010_100_0_000101010001;
      patterns[5397] = 29'b0_001010100010_101_1_000010101000;
      patterns[5398] = 29'b0_001010100010_110_0_001010100010;
      patterns[5399] = 29'b0_001010100010_111_0_001010100010;
      patterns[5400] = 29'b0_001010100011_000_0_001010100011;
      patterns[5401] = 29'b0_001010100011_001_0_100011001010;
      patterns[5402] = 29'b0_001010100011_010_0_010101000110;
      patterns[5403] = 29'b0_001010100011_011_0_101010001100;
      patterns[5404] = 29'b0_001010100011_100_1_000101010001;
      patterns[5405] = 29'b0_001010100011_101_1_100010101000;
      patterns[5406] = 29'b0_001010100011_110_0_001010100011;
      patterns[5407] = 29'b0_001010100011_111_0_001010100011;
      patterns[5408] = 29'b0_001010100100_000_0_001010100100;
      patterns[5409] = 29'b0_001010100100_001_0_100100001010;
      patterns[5410] = 29'b0_001010100100_010_0_010101001000;
      patterns[5411] = 29'b0_001010100100_011_0_101010010000;
      patterns[5412] = 29'b0_001010100100_100_0_000101010010;
      patterns[5413] = 29'b0_001010100100_101_0_000010101001;
      patterns[5414] = 29'b0_001010100100_110_0_001010100100;
      patterns[5415] = 29'b0_001010100100_111_0_001010100100;
      patterns[5416] = 29'b0_001010100101_000_0_001010100101;
      patterns[5417] = 29'b0_001010100101_001_0_100101001010;
      patterns[5418] = 29'b0_001010100101_010_0_010101001010;
      patterns[5419] = 29'b0_001010100101_011_0_101010010100;
      patterns[5420] = 29'b0_001010100101_100_1_000101010010;
      patterns[5421] = 29'b0_001010100101_101_0_100010101001;
      patterns[5422] = 29'b0_001010100101_110_0_001010100101;
      patterns[5423] = 29'b0_001010100101_111_0_001010100101;
      patterns[5424] = 29'b0_001010100110_000_0_001010100110;
      patterns[5425] = 29'b0_001010100110_001_0_100110001010;
      patterns[5426] = 29'b0_001010100110_010_0_010101001100;
      patterns[5427] = 29'b0_001010100110_011_0_101010011000;
      patterns[5428] = 29'b0_001010100110_100_0_000101010011;
      patterns[5429] = 29'b0_001010100110_101_1_000010101001;
      patterns[5430] = 29'b0_001010100110_110_0_001010100110;
      patterns[5431] = 29'b0_001010100110_111_0_001010100110;
      patterns[5432] = 29'b0_001010100111_000_0_001010100111;
      patterns[5433] = 29'b0_001010100111_001_0_100111001010;
      patterns[5434] = 29'b0_001010100111_010_0_010101001110;
      patterns[5435] = 29'b0_001010100111_011_0_101010011100;
      patterns[5436] = 29'b0_001010100111_100_1_000101010011;
      patterns[5437] = 29'b0_001010100111_101_1_100010101001;
      patterns[5438] = 29'b0_001010100111_110_0_001010100111;
      patterns[5439] = 29'b0_001010100111_111_0_001010100111;
      patterns[5440] = 29'b0_001010101000_000_0_001010101000;
      patterns[5441] = 29'b0_001010101000_001_0_101000001010;
      patterns[5442] = 29'b0_001010101000_010_0_010101010000;
      patterns[5443] = 29'b0_001010101000_011_0_101010100000;
      patterns[5444] = 29'b0_001010101000_100_0_000101010100;
      patterns[5445] = 29'b0_001010101000_101_0_000010101010;
      patterns[5446] = 29'b0_001010101000_110_0_001010101000;
      patterns[5447] = 29'b0_001010101000_111_0_001010101000;
      patterns[5448] = 29'b0_001010101001_000_0_001010101001;
      patterns[5449] = 29'b0_001010101001_001_0_101001001010;
      patterns[5450] = 29'b0_001010101001_010_0_010101010010;
      patterns[5451] = 29'b0_001010101001_011_0_101010100100;
      patterns[5452] = 29'b0_001010101001_100_1_000101010100;
      patterns[5453] = 29'b0_001010101001_101_0_100010101010;
      patterns[5454] = 29'b0_001010101001_110_0_001010101001;
      patterns[5455] = 29'b0_001010101001_111_0_001010101001;
      patterns[5456] = 29'b0_001010101010_000_0_001010101010;
      patterns[5457] = 29'b0_001010101010_001_0_101010001010;
      patterns[5458] = 29'b0_001010101010_010_0_010101010100;
      patterns[5459] = 29'b0_001010101010_011_0_101010101000;
      patterns[5460] = 29'b0_001010101010_100_0_000101010101;
      patterns[5461] = 29'b0_001010101010_101_1_000010101010;
      patterns[5462] = 29'b0_001010101010_110_0_001010101010;
      patterns[5463] = 29'b0_001010101010_111_0_001010101010;
      patterns[5464] = 29'b0_001010101011_000_0_001010101011;
      patterns[5465] = 29'b0_001010101011_001_0_101011001010;
      patterns[5466] = 29'b0_001010101011_010_0_010101010110;
      patterns[5467] = 29'b0_001010101011_011_0_101010101100;
      patterns[5468] = 29'b0_001010101011_100_1_000101010101;
      patterns[5469] = 29'b0_001010101011_101_1_100010101010;
      patterns[5470] = 29'b0_001010101011_110_0_001010101011;
      patterns[5471] = 29'b0_001010101011_111_0_001010101011;
      patterns[5472] = 29'b0_001010101100_000_0_001010101100;
      patterns[5473] = 29'b0_001010101100_001_0_101100001010;
      patterns[5474] = 29'b0_001010101100_010_0_010101011000;
      patterns[5475] = 29'b0_001010101100_011_0_101010110000;
      patterns[5476] = 29'b0_001010101100_100_0_000101010110;
      patterns[5477] = 29'b0_001010101100_101_0_000010101011;
      patterns[5478] = 29'b0_001010101100_110_0_001010101100;
      patterns[5479] = 29'b0_001010101100_111_0_001010101100;
      patterns[5480] = 29'b0_001010101101_000_0_001010101101;
      patterns[5481] = 29'b0_001010101101_001_0_101101001010;
      patterns[5482] = 29'b0_001010101101_010_0_010101011010;
      patterns[5483] = 29'b0_001010101101_011_0_101010110100;
      patterns[5484] = 29'b0_001010101101_100_1_000101010110;
      patterns[5485] = 29'b0_001010101101_101_0_100010101011;
      patterns[5486] = 29'b0_001010101101_110_0_001010101101;
      patterns[5487] = 29'b0_001010101101_111_0_001010101101;
      patterns[5488] = 29'b0_001010101110_000_0_001010101110;
      patterns[5489] = 29'b0_001010101110_001_0_101110001010;
      patterns[5490] = 29'b0_001010101110_010_0_010101011100;
      patterns[5491] = 29'b0_001010101110_011_0_101010111000;
      patterns[5492] = 29'b0_001010101110_100_0_000101010111;
      patterns[5493] = 29'b0_001010101110_101_1_000010101011;
      patterns[5494] = 29'b0_001010101110_110_0_001010101110;
      patterns[5495] = 29'b0_001010101110_111_0_001010101110;
      patterns[5496] = 29'b0_001010101111_000_0_001010101111;
      patterns[5497] = 29'b0_001010101111_001_0_101111001010;
      patterns[5498] = 29'b0_001010101111_010_0_010101011110;
      patterns[5499] = 29'b0_001010101111_011_0_101010111100;
      patterns[5500] = 29'b0_001010101111_100_1_000101010111;
      patterns[5501] = 29'b0_001010101111_101_1_100010101011;
      patterns[5502] = 29'b0_001010101111_110_0_001010101111;
      patterns[5503] = 29'b0_001010101111_111_0_001010101111;
      patterns[5504] = 29'b0_001010110000_000_0_001010110000;
      patterns[5505] = 29'b0_001010110000_001_0_110000001010;
      patterns[5506] = 29'b0_001010110000_010_0_010101100000;
      patterns[5507] = 29'b0_001010110000_011_0_101011000000;
      patterns[5508] = 29'b0_001010110000_100_0_000101011000;
      patterns[5509] = 29'b0_001010110000_101_0_000010101100;
      patterns[5510] = 29'b0_001010110000_110_0_001010110000;
      patterns[5511] = 29'b0_001010110000_111_0_001010110000;
      patterns[5512] = 29'b0_001010110001_000_0_001010110001;
      patterns[5513] = 29'b0_001010110001_001_0_110001001010;
      patterns[5514] = 29'b0_001010110001_010_0_010101100010;
      patterns[5515] = 29'b0_001010110001_011_0_101011000100;
      patterns[5516] = 29'b0_001010110001_100_1_000101011000;
      patterns[5517] = 29'b0_001010110001_101_0_100010101100;
      patterns[5518] = 29'b0_001010110001_110_0_001010110001;
      patterns[5519] = 29'b0_001010110001_111_0_001010110001;
      patterns[5520] = 29'b0_001010110010_000_0_001010110010;
      patterns[5521] = 29'b0_001010110010_001_0_110010001010;
      patterns[5522] = 29'b0_001010110010_010_0_010101100100;
      patterns[5523] = 29'b0_001010110010_011_0_101011001000;
      patterns[5524] = 29'b0_001010110010_100_0_000101011001;
      patterns[5525] = 29'b0_001010110010_101_1_000010101100;
      patterns[5526] = 29'b0_001010110010_110_0_001010110010;
      patterns[5527] = 29'b0_001010110010_111_0_001010110010;
      patterns[5528] = 29'b0_001010110011_000_0_001010110011;
      patterns[5529] = 29'b0_001010110011_001_0_110011001010;
      patterns[5530] = 29'b0_001010110011_010_0_010101100110;
      patterns[5531] = 29'b0_001010110011_011_0_101011001100;
      patterns[5532] = 29'b0_001010110011_100_1_000101011001;
      patterns[5533] = 29'b0_001010110011_101_1_100010101100;
      patterns[5534] = 29'b0_001010110011_110_0_001010110011;
      patterns[5535] = 29'b0_001010110011_111_0_001010110011;
      patterns[5536] = 29'b0_001010110100_000_0_001010110100;
      patterns[5537] = 29'b0_001010110100_001_0_110100001010;
      patterns[5538] = 29'b0_001010110100_010_0_010101101000;
      patterns[5539] = 29'b0_001010110100_011_0_101011010000;
      patterns[5540] = 29'b0_001010110100_100_0_000101011010;
      patterns[5541] = 29'b0_001010110100_101_0_000010101101;
      patterns[5542] = 29'b0_001010110100_110_0_001010110100;
      patterns[5543] = 29'b0_001010110100_111_0_001010110100;
      patterns[5544] = 29'b0_001010110101_000_0_001010110101;
      patterns[5545] = 29'b0_001010110101_001_0_110101001010;
      patterns[5546] = 29'b0_001010110101_010_0_010101101010;
      patterns[5547] = 29'b0_001010110101_011_0_101011010100;
      patterns[5548] = 29'b0_001010110101_100_1_000101011010;
      patterns[5549] = 29'b0_001010110101_101_0_100010101101;
      patterns[5550] = 29'b0_001010110101_110_0_001010110101;
      patterns[5551] = 29'b0_001010110101_111_0_001010110101;
      patterns[5552] = 29'b0_001010110110_000_0_001010110110;
      patterns[5553] = 29'b0_001010110110_001_0_110110001010;
      patterns[5554] = 29'b0_001010110110_010_0_010101101100;
      patterns[5555] = 29'b0_001010110110_011_0_101011011000;
      patterns[5556] = 29'b0_001010110110_100_0_000101011011;
      patterns[5557] = 29'b0_001010110110_101_1_000010101101;
      patterns[5558] = 29'b0_001010110110_110_0_001010110110;
      patterns[5559] = 29'b0_001010110110_111_0_001010110110;
      patterns[5560] = 29'b0_001010110111_000_0_001010110111;
      patterns[5561] = 29'b0_001010110111_001_0_110111001010;
      patterns[5562] = 29'b0_001010110111_010_0_010101101110;
      patterns[5563] = 29'b0_001010110111_011_0_101011011100;
      patterns[5564] = 29'b0_001010110111_100_1_000101011011;
      patterns[5565] = 29'b0_001010110111_101_1_100010101101;
      patterns[5566] = 29'b0_001010110111_110_0_001010110111;
      patterns[5567] = 29'b0_001010110111_111_0_001010110111;
      patterns[5568] = 29'b0_001010111000_000_0_001010111000;
      patterns[5569] = 29'b0_001010111000_001_0_111000001010;
      patterns[5570] = 29'b0_001010111000_010_0_010101110000;
      patterns[5571] = 29'b0_001010111000_011_0_101011100000;
      patterns[5572] = 29'b0_001010111000_100_0_000101011100;
      patterns[5573] = 29'b0_001010111000_101_0_000010101110;
      patterns[5574] = 29'b0_001010111000_110_0_001010111000;
      patterns[5575] = 29'b0_001010111000_111_0_001010111000;
      patterns[5576] = 29'b0_001010111001_000_0_001010111001;
      patterns[5577] = 29'b0_001010111001_001_0_111001001010;
      patterns[5578] = 29'b0_001010111001_010_0_010101110010;
      patterns[5579] = 29'b0_001010111001_011_0_101011100100;
      patterns[5580] = 29'b0_001010111001_100_1_000101011100;
      patterns[5581] = 29'b0_001010111001_101_0_100010101110;
      patterns[5582] = 29'b0_001010111001_110_0_001010111001;
      patterns[5583] = 29'b0_001010111001_111_0_001010111001;
      patterns[5584] = 29'b0_001010111010_000_0_001010111010;
      patterns[5585] = 29'b0_001010111010_001_0_111010001010;
      patterns[5586] = 29'b0_001010111010_010_0_010101110100;
      patterns[5587] = 29'b0_001010111010_011_0_101011101000;
      patterns[5588] = 29'b0_001010111010_100_0_000101011101;
      patterns[5589] = 29'b0_001010111010_101_1_000010101110;
      patterns[5590] = 29'b0_001010111010_110_0_001010111010;
      patterns[5591] = 29'b0_001010111010_111_0_001010111010;
      patterns[5592] = 29'b0_001010111011_000_0_001010111011;
      patterns[5593] = 29'b0_001010111011_001_0_111011001010;
      patterns[5594] = 29'b0_001010111011_010_0_010101110110;
      patterns[5595] = 29'b0_001010111011_011_0_101011101100;
      patterns[5596] = 29'b0_001010111011_100_1_000101011101;
      patterns[5597] = 29'b0_001010111011_101_1_100010101110;
      patterns[5598] = 29'b0_001010111011_110_0_001010111011;
      patterns[5599] = 29'b0_001010111011_111_0_001010111011;
      patterns[5600] = 29'b0_001010111100_000_0_001010111100;
      patterns[5601] = 29'b0_001010111100_001_0_111100001010;
      patterns[5602] = 29'b0_001010111100_010_0_010101111000;
      patterns[5603] = 29'b0_001010111100_011_0_101011110000;
      patterns[5604] = 29'b0_001010111100_100_0_000101011110;
      patterns[5605] = 29'b0_001010111100_101_0_000010101111;
      patterns[5606] = 29'b0_001010111100_110_0_001010111100;
      patterns[5607] = 29'b0_001010111100_111_0_001010111100;
      patterns[5608] = 29'b0_001010111101_000_0_001010111101;
      patterns[5609] = 29'b0_001010111101_001_0_111101001010;
      patterns[5610] = 29'b0_001010111101_010_0_010101111010;
      patterns[5611] = 29'b0_001010111101_011_0_101011110100;
      patterns[5612] = 29'b0_001010111101_100_1_000101011110;
      patterns[5613] = 29'b0_001010111101_101_0_100010101111;
      patterns[5614] = 29'b0_001010111101_110_0_001010111101;
      patterns[5615] = 29'b0_001010111101_111_0_001010111101;
      patterns[5616] = 29'b0_001010111110_000_0_001010111110;
      patterns[5617] = 29'b0_001010111110_001_0_111110001010;
      patterns[5618] = 29'b0_001010111110_010_0_010101111100;
      patterns[5619] = 29'b0_001010111110_011_0_101011111000;
      patterns[5620] = 29'b0_001010111110_100_0_000101011111;
      patterns[5621] = 29'b0_001010111110_101_1_000010101111;
      patterns[5622] = 29'b0_001010111110_110_0_001010111110;
      patterns[5623] = 29'b0_001010111110_111_0_001010111110;
      patterns[5624] = 29'b0_001010111111_000_0_001010111111;
      patterns[5625] = 29'b0_001010111111_001_0_111111001010;
      patterns[5626] = 29'b0_001010111111_010_0_010101111110;
      patterns[5627] = 29'b0_001010111111_011_0_101011111100;
      patterns[5628] = 29'b0_001010111111_100_1_000101011111;
      patterns[5629] = 29'b0_001010111111_101_1_100010101111;
      patterns[5630] = 29'b0_001010111111_110_0_001010111111;
      patterns[5631] = 29'b0_001010111111_111_0_001010111111;
      patterns[5632] = 29'b0_001011000000_000_0_001011000000;
      patterns[5633] = 29'b0_001011000000_001_0_000000001011;
      patterns[5634] = 29'b0_001011000000_010_0_010110000000;
      patterns[5635] = 29'b0_001011000000_011_0_101100000000;
      patterns[5636] = 29'b0_001011000000_100_0_000101100000;
      patterns[5637] = 29'b0_001011000000_101_0_000010110000;
      patterns[5638] = 29'b0_001011000000_110_0_001011000000;
      patterns[5639] = 29'b0_001011000000_111_0_001011000000;
      patterns[5640] = 29'b0_001011000001_000_0_001011000001;
      patterns[5641] = 29'b0_001011000001_001_0_000001001011;
      patterns[5642] = 29'b0_001011000001_010_0_010110000010;
      patterns[5643] = 29'b0_001011000001_011_0_101100000100;
      patterns[5644] = 29'b0_001011000001_100_1_000101100000;
      patterns[5645] = 29'b0_001011000001_101_0_100010110000;
      patterns[5646] = 29'b0_001011000001_110_0_001011000001;
      patterns[5647] = 29'b0_001011000001_111_0_001011000001;
      patterns[5648] = 29'b0_001011000010_000_0_001011000010;
      patterns[5649] = 29'b0_001011000010_001_0_000010001011;
      patterns[5650] = 29'b0_001011000010_010_0_010110000100;
      patterns[5651] = 29'b0_001011000010_011_0_101100001000;
      patterns[5652] = 29'b0_001011000010_100_0_000101100001;
      patterns[5653] = 29'b0_001011000010_101_1_000010110000;
      patterns[5654] = 29'b0_001011000010_110_0_001011000010;
      patterns[5655] = 29'b0_001011000010_111_0_001011000010;
      patterns[5656] = 29'b0_001011000011_000_0_001011000011;
      patterns[5657] = 29'b0_001011000011_001_0_000011001011;
      patterns[5658] = 29'b0_001011000011_010_0_010110000110;
      patterns[5659] = 29'b0_001011000011_011_0_101100001100;
      patterns[5660] = 29'b0_001011000011_100_1_000101100001;
      patterns[5661] = 29'b0_001011000011_101_1_100010110000;
      patterns[5662] = 29'b0_001011000011_110_0_001011000011;
      patterns[5663] = 29'b0_001011000011_111_0_001011000011;
      patterns[5664] = 29'b0_001011000100_000_0_001011000100;
      patterns[5665] = 29'b0_001011000100_001_0_000100001011;
      patterns[5666] = 29'b0_001011000100_010_0_010110001000;
      patterns[5667] = 29'b0_001011000100_011_0_101100010000;
      patterns[5668] = 29'b0_001011000100_100_0_000101100010;
      patterns[5669] = 29'b0_001011000100_101_0_000010110001;
      patterns[5670] = 29'b0_001011000100_110_0_001011000100;
      patterns[5671] = 29'b0_001011000100_111_0_001011000100;
      patterns[5672] = 29'b0_001011000101_000_0_001011000101;
      patterns[5673] = 29'b0_001011000101_001_0_000101001011;
      patterns[5674] = 29'b0_001011000101_010_0_010110001010;
      patterns[5675] = 29'b0_001011000101_011_0_101100010100;
      patterns[5676] = 29'b0_001011000101_100_1_000101100010;
      patterns[5677] = 29'b0_001011000101_101_0_100010110001;
      patterns[5678] = 29'b0_001011000101_110_0_001011000101;
      patterns[5679] = 29'b0_001011000101_111_0_001011000101;
      patterns[5680] = 29'b0_001011000110_000_0_001011000110;
      patterns[5681] = 29'b0_001011000110_001_0_000110001011;
      patterns[5682] = 29'b0_001011000110_010_0_010110001100;
      patterns[5683] = 29'b0_001011000110_011_0_101100011000;
      patterns[5684] = 29'b0_001011000110_100_0_000101100011;
      patterns[5685] = 29'b0_001011000110_101_1_000010110001;
      patterns[5686] = 29'b0_001011000110_110_0_001011000110;
      patterns[5687] = 29'b0_001011000110_111_0_001011000110;
      patterns[5688] = 29'b0_001011000111_000_0_001011000111;
      patterns[5689] = 29'b0_001011000111_001_0_000111001011;
      patterns[5690] = 29'b0_001011000111_010_0_010110001110;
      patterns[5691] = 29'b0_001011000111_011_0_101100011100;
      patterns[5692] = 29'b0_001011000111_100_1_000101100011;
      patterns[5693] = 29'b0_001011000111_101_1_100010110001;
      patterns[5694] = 29'b0_001011000111_110_0_001011000111;
      patterns[5695] = 29'b0_001011000111_111_0_001011000111;
      patterns[5696] = 29'b0_001011001000_000_0_001011001000;
      patterns[5697] = 29'b0_001011001000_001_0_001000001011;
      patterns[5698] = 29'b0_001011001000_010_0_010110010000;
      patterns[5699] = 29'b0_001011001000_011_0_101100100000;
      patterns[5700] = 29'b0_001011001000_100_0_000101100100;
      patterns[5701] = 29'b0_001011001000_101_0_000010110010;
      patterns[5702] = 29'b0_001011001000_110_0_001011001000;
      patterns[5703] = 29'b0_001011001000_111_0_001011001000;
      patterns[5704] = 29'b0_001011001001_000_0_001011001001;
      patterns[5705] = 29'b0_001011001001_001_0_001001001011;
      patterns[5706] = 29'b0_001011001001_010_0_010110010010;
      patterns[5707] = 29'b0_001011001001_011_0_101100100100;
      patterns[5708] = 29'b0_001011001001_100_1_000101100100;
      patterns[5709] = 29'b0_001011001001_101_0_100010110010;
      patterns[5710] = 29'b0_001011001001_110_0_001011001001;
      patterns[5711] = 29'b0_001011001001_111_0_001011001001;
      patterns[5712] = 29'b0_001011001010_000_0_001011001010;
      patterns[5713] = 29'b0_001011001010_001_0_001010001011;
      patterns[5714] = 29'b0_001011001010_010_0_010110010100;
      patterns[5715] = 29'b0_001011001010_011_0_101100101000;
      patterns[5716] = 29'b0_001011001010_100_0_000101100101;
      patterns[5717] = 29'b0_001011001010_101_1_000010110010;
      patterns[5718] = 29'b0_001011001010_110_0_001011001010;
      patterns[5719] = 29'b0_001011001010_111_0_001011001010;
      patterns[5720] = 29'b0_001011001011_000_0_001011001011;
      patterns[5721] = 29'b0_001011001011_001_0_001011001011;
      patterns[5722] = 29'b0_001011001011_010_0_010110010110;
      patterns[5723] = 29'b0_001011001011_011_0_101100101100;
      patterns[5724] = 29'b0_001011001011_100_1_000101100101;
      patterns[5725] = 29'b0_001011001011_101_1_100010110010;
      patterns[5726] = 29'b0_001011001011_110_0_001011001011;
      patterns[5727] = 29'b0_001011001011_111_0_001011001011;
      patterns[5728] = 29'b0_001011001100_000_0_001011001100;
      patterns[5729] = 29'b0_001011001100_001_0_001100001011;
      patterns[5730] = 29'b0_001011001100_010_0_010110011000;
      patterns[5731] = 29'b0_001011001100_011_0_101100110000;
      patterns[5732] = 29'b0_001011001100_100_0_000101100110;
      patterns[5733] = 29'b0_001011001100_101_0_000010110011;
      patterns[5734] = 29'b0_001011001100_110_0_001011001100;
      patterns[5735] = 29'b0_001011001100_111_0_001011001100;
      patterns[5736] = 29'b0_001011001101_000_0_001011001101;
      patterns[5737] = 29'b0_001011001101_001_0_001101001011;
      patterns[5738] = 29'b0_001011001101_010_0_010110011010;
      patterns[5739] = 29'b0_001011001101_011_0_101100110100;
      patterns[5740] = 29'b0_001011001101_100_1_000101100110;
      patterns[5741] = 29'b0_001011001101_101_0_100010110011;
      patterns[5742] = 29'b0_001011001101_110_0_001011001101;
      patterns[5743] = 29'b0_001011001101_111_0_001011001101;
      patterns[5744] = 29'b0_001011001110_000_0_001011001110;
      patterns[5745] = 29'b0_001011001110_001_0_001110001011;
      patterns[5746] = 29'b0_001011001110_010_0_010110011100;
      patterns[5747] = 29'b0_001011001110_011_0_101100111000;
      patterns[5748] = 29'b0_001011001110_100_0_000101100111;
      patterns[5749] = 29'b0_001011001110_101_1_000010110011;
      patterns[5750] = 29'b0_001011001110_110_0_001011001110;
      patterns[5751] = 29'b0_001011001110_111_0_001011001110;
      patterns[5752] = 29'b0_001011001111_000_0_001011001111;
      patterns[5753] = 29'b0_001011001111_001_0_001111001011;
      patterns[5754] = 29'b0_001011001111_010_0_010110011110;
      patterns[5755] = 29'b0_001011001111_011_0_101100111100;
      patterns[5756] = 29'b0_001011001111_100_1_000101100111;
      patterns[5757] = 29'b0_001011001111_101_1_100010110011;
      patterns[5758] = 29'b0_001011001111_110_0_001011001111;
      patterns[5759] = 29'b0_001011001111_111_0_001011001111;
      patterns[5760] = 29'b0_001011010000_000_0_001011010000;
      patterns[5761] = 29'b0_001011010000_001_0_010000001011;
      patterns[5762] = 29'b0_001011010000_010_0_010110100000;
      patterns[5763] = 29'b0_001011010000_011_0_101101000000;
      patterns[5764] = 29'b0_001011010000_100_0_000101101000;
      patterns[5765] = 29'b0_001011010000_101_0_000010110100;
      patterns[5766] = 29'b0_001011010000_110_0_001011010000;
      patterns[5767] = 29'b0_001011010000_111_0_001011010000;
      patterns[5768] = 29'b0_001011010001_000_0_001011010001;
      patterns[5769] = 29'b0_001011010001_001_0_010001001011;
      patterns[5770] = 29'b0_001011010001_010_0_010110100010;
      patterns[5771] = 29'b0_001011010001_011_0_101101000100;
      patterns[5772] = 29'b0_001011010001_100_1_000101101000;
      patterns[5773] = 29'b0_001011010001_101_0_100010110100;
      patterns[5774] = 29'b0_001011010001_110_0_001011010001;
      patterns[5775] = 29'b0_001011010001_111_0_001011010001;
      patterns[5776] = 29'b0_001011010010_000_0_001011010010;
      patterns[5777] = 29'b0_001011010010_001_0_010010001011;
      patterns[5778] = 29'b0_001011010010_010_0_010110100100;
      patterns[5779] = 29'b0_001011010010_011_0_101101001000;
      patterns[5780] = 29'b0_001011010010_100_0_000101101001;
      patterns[5781] = 29'b0_001011010010_101_1_000010110100;
      patterns[5782] = 29'b0_001011010010_110_0_001011010010;
      patterns[5783] = 29'b0_001011010010_111_0_001011010010;
      patterns[5784] = 29'b0_001011010011_000_0_001011010011;
      patterns[5785] = 29'b0_001011010011_001_0_010011001011;
      patterns[5786] = 29'b0_001011010011_010_0_010110100110;
      patterns[5787] = 29'b0_001011010011_011_0_101101001100;
      patterns[5788] = 29'b0_001011010011_100_1_000101101001;
      patterns[5789] = 29'b0_001011010011_101_1_100010110100;
      patterns[5790] = 29'b0_001011010011_110_0_001011010011;
      patterns[5791] = 29'b0_001011010011_111_0_001011010011;
      patterns[5792] = 29'b0_001011010100_000_0_001011010100;
      patterns[5793] = 29'b0_001011010100_001_0_010100001011;
      patterns[5794] = 29'b0_001011010100_010_0_010110101000;
      patterns[5795] = 29'b0_001011010100_011_0_101101010000;
      patterns[5796] = 29'b0_001011010100_100_0_000101101010;
      patterns[5797] = 29'b0_001011010100_101_0_000010110101;
      patterns[5798] = 29'b0_001011010100_110_0_001011010100;
      patterns[5799] = 29'b0_001011010100_111_0_001011010100;
      patterns[5800] = 29'b0_001011010101_000_0_001011010101;
      patterns[5801] = 29'b0_001011010101_001_0_010101001011;
      patterns[5802] = 29'b0_001011010101_010_0_010110101010;
      patterns[5803] = 29'b0_001011010101_011_0_101101010100;
      patterns[5804] = 29'b0_001011010101_100_1_000101101010;
      patterns[5805] = 29'b0_001011010101_101_0_100010110101;
      patterns[5806] = 29'b0_001011010101_110_0_001011010101;
      patterns[5807] = 29'b0_001011010101_111_0_001011010101;
      patterns[5808] = 29'b0_001011010110_000_0_001011010110;
      patterns[5809] = 29'b0_001011010110_001_0_010110001011;
      patterns[5810] = 29'b0_001011010110_010_0_010110101100;
      patterns[5811] = 29'b0_001011010110_011_0_101101011000;
      patterns[5812] = 29'b0_001011010110_100_0_000101101011;
      patterns[5813] = 29'b0_001011010110_101_1_000010110101;
      patterns[5814] = 29'b0_001011010110_110_0_001011010110;
      patterns[5815] = 29'b0_001011010110_111_0_001011010110;
      patterns[5816] = 29'b0_001011010111_000_0_001011010111;
      patterns[5817] = 29'b0_001011010111_001_0_010111001011;
      patterns[5818] = 29'b0_001011010111_010_0_010110101110;
      patterns[5819] = 29'b0_001011010111_011_0_101101011100;
      patterns[5820] = 29'b0_001011010111_100_1_000101101011;
      patterns[5821] = 29'b0_001011010111_101_1_100010110101;
      patterns[5822] = 29'b0_001011010111_110_0_001011010111;
      patterns[5823] = 29'b0_001011010111_111_0_001011010111;
      patterns[5824] = 29'b0_001011011000_000_0_001011011000;
      patterns[5825] = 29'b0_001011011000_001_0_011000001011;
      patterns[5826] = 29'b0_001011011000_010_0_010110110000;
      patterns[5827] = 29'b0_001011011000_011_0_101101100000;
      patterns[5828] = 29'b0_001011011000_100_0_000101101100;
      patterns[5829] = 29'b0_001011011000_101_0_000010110110;
      patterns[5830] = 29'b0_001011011000_110_0_001011011000;
      patterns[5831] = 29'b0_001011011000_111_0_001011011000;
      patterns[5832] = 29'b0_001011011001_000_0_001011011001;
      patterns[5833] = 29'b0_001011011001_001_0_011001001011;
      patterns[5834] = 29'b0_001011011001_010_0_010110110010;
      patterns[5835] = 29'b0_001011011001_011_0_101101100100;
      patterns[5836] = 29'b0_001011011001_100_1_000101101100;
      patterns[5837] = 29'b0_001011011001_101_0_100010110110;
      patterns[5838] = 29'b0_001011011001_110_0_001011011001;
      patterns[5839] = 29'b0_001011011001_111_0_001011011001;
      patterns[5840] = 29'b0_001011011010_000_0_001011011010;
      patterns[5841] = 29'b0_001011011010_001_0_011010001011;
      patterns[5842] = 29'b0_001011011010_010_0_010110110100;
      patterns[5843] = 29'b0_001011011010_011_0_101101101000;
      patterns[5844] = 29'b0_001011011010_100_0_000101101101;
      patterns[5845] = 29'b0_001011011010_101_1_000010110110;
      patterns[5846] = 29'b0_001011011010_110_0_001011011010;
      patterns[5847] = 29'b0_001011011010_111_0_001011011010;
      patterns[5848] = 29'b0_001011011011_000_0_001011011011;
      patterns[5849] = 29'b0_001011011011_001_0_011011001011;
      patterns[5850] = 29'b0_001011011011_010_0_010110110110;
      patterns[5851] = 29'b0_001011011011_011_0_101101101100;
      patterns[5852] = 29'b0_001011011011_100_1_000101101101;
      patterns[5853] = 29'b0_001011011011_101_1_100010110110;
      patterns[5854] = 29'b0_001011011011_110_0_001011011011;
      patterns[5855] = 29'b0_001011011011_111_0_001011011011;
      patterns[5856] = 29'b0_001011011100_000_0_001011011100;
      patterns[5857] = 29'b0_001011011100_001_0_011100001011;
      patterns[5858] = 29'b0_001011011100_010_0_010110111000;
      patterns[5859] = 29'b0_001011011100_011_0_101101110000;
      patterns[5860] = 29'b0_001011011100_100_0_000101101110;
      patterns[5861] = 29'b0_001011011100_101_0_000010110111;
      patterns[5862] = 29'b0_001011011100_110_0_001011011100;
      patterns[5863] = 29'b0_001011011100_111_0_001011011100;
      patterns[5864] = 29'b0_001011011101_000_0_001011011101;
      patterns[5865] = 29'b0_001011011101_001_0_011101001011;
      patterns[5866] = 29'b0_001011011101_010_0_010110111010;
      patterns[5867] = 29'b0_001011011101_011_0_101101110100;
      patterns[5868] = 29'b0_001011011101_100_1_000101101110;
      patterns[5869] = 29'b0_001011011101_101_0_100010110111;
      patterns[5870] = 29'b0_001011011101_110_0_001011011101;
      patterns[5871] = 29'b0_001011011101_111_0_001011011101;
      patterns[5872] = 29'b0_001011011110_000_0_001011011110;
      patterns[5873] = 29'b0_001011011110_001_0_011110001011;
      patterns[5874] = 29'b0_001011011110_010_0_010110111100;
      patterns[5875] = 29'b0_001011011110_011_0_101101111000;
      patterns[5876] = 29'b0_001011011110_100_0_000101101111;
      patterns[5877] = 29'b0_001011011110_101_1_000010110111;
      patterns[5878] = 29'b0_001011011110_110_0_001011011110;
      patterns[5879] = 29'b0_001011011110_111_0_001011011110;
      patterns[5880] = 29'b0_001011011111_000_0_001011011111;
      patterns[5881] = 29'b0_001011011111_001_0_011111001011;
      patterns[5882] = 29'b0_001011011111_010_0_010110111110;
      patterns[5883] = 29'b0_001011011111_011_0_101101111100;
      patterns[5884] = 29'b0_001011011111_100_1_000101101111;
      patterns[5885] = 29'b0_001011011111_101_1_100010110111;
      patterns[5886] = 29'b0_001011011111_110_0_001011011111;
      patterns[5887] = 29'b0_001011011111_111_0_001011011111;
      patterns[5888] = 29'b0_001011100000_000_0_001011100000;
      patterns[5889] = 29'b0_001011100000_001_0_100000001011;
      patterns[5890] = 29'b0_001011100000_010_0_010111000000;
      patterns[5891] = 29'b0_001011100000_011_0_101110000000;
      patterns[5892] = 29'b0_001011100000_100_0_000101110000;
      patterns[5893] = 29'b0_001011100000_101_0_000010111000;
      patterns[5894] = 29'b0_001011100000_110_0_001011100000;
      patterns[5895] = 29'b0_001011100000_111_0_001011100000;
      patterns[5896] = 29'b0_001011100001_000_0_001011100001;
      patterns[5897] = 29'b0_001011100001_001_0_100001001011;
      patterns[5898] = 29'b0_001011100001_010_0_010111000010;
      patterns[5899] = 29'b0_001011100001_011_0_101110000100;
      patterns[5900] = 29'b0_001011100001_100_1_000101110000;
      patterns[5901] = 29'b0_001011100001_101_0_100010111000;
      patterns[5902] = 29'b0_001011100001_110_0_001011100001;
      patterns[5903] = 29'b0_001011100001_111_0_001011100001;
      patterns[5904] = 29'b0_001011100010_000_0_001011100010;
      patterns[5905] = 29'b0_001011100010_001_0_100010001011;
      patterns[5906] = 29'b0_001011100010_010_0_010111000100;
      patterns[5907] = 29'b0_001011100010_011_0_101110001000;
      patterns[5908] = 29'b0_001011100010_100_0_000101110001;
      patterns[5909] = 29'b0_001011100010_101_1_000010111000;
      patterns[5910] = 29'b0_001011100010_110_0_001011100010;
      patterns[5911] = 29'b0_001011100010_111_0_001011100010;
      patterns[5912] = 29'b0_001011100011_000_0_001011100011;
      patterns[5913] = 29'b0_001011100011_001_0_100011001011;
      patterns[5914] = 29'b0_001011100011_010_0_010111000110;
      patterns[5915] = 29'b0_001011100011_011_0_101110001100;
      patterns[5916] = 29'b0_001011100011_100_1_000101110001;
      patterns[5917] = 29'b0_001011100011_101_1_100010111000;
      patterns[5918] = 29'b0_001011100011_110_0_001011100011;
      patterns[5919] = 29'b0_001011100011_111_0_001011100011;
      patterns[5920] = 29'b0_001011100100_000_0_001011100100;
      patterns[5921] = 29'b0_001011100100_001_0_100100001011;
      patterns[5922] = 29'b0_001011100100_010_0_010111001000;
      patterns[5923] = 29'b0_001011100100_011_0_101110010000;
      patterns[5924] = 29'b0_001011100100_100_0_000101110010;
      patterns[5925] = 29'b0_001011100100_101_0_000010111001;
      patterns[5926] = 29'b0_001011100100_110_0_001011100100;
      patterns[5927] = 29'b0_001011100100_111_0_001011100100;
      patterns[5928] = 29'b0_001011100101_000_0_001011100101;
      patterns[5929] = 29'b0_001011100101_001_0_100101001011;
      patterns[5930] = 29'b0_001011100101_010_0_010111001010;
      patterns[5931] = 29'b0_001011100101_011_0_101110010100;
      patterns[5932] = 29'b0_001011100101_100_1_000101110010;
      patterns[5933] = 29'b0_001011100101_101_0_100010111001;
      patterns[5934] = 29'b0_001011100101_110_0_001011100101;
      patterns[5935] = 29'b0_001011100101_111_0_001011100101;
      patterns[5936] = 29'b0_001011100110_000_0_001011100110;
      patterns[5937] = 29'b0_001011100110_001_0_100110001011;
      patterns[5938] = 29'b0_001011100110_010_0_010111001100;
      patterns[5939] = 29'b0_001011100110_011_0_101110011000;
      patterns[5940] = 29'b0_001011100110_100_0_000101110011;
      patterns[5941] = 29'b0_001011100110_101_1_000010111001;
      patterns[5942] = 29'b0_001011100110_110_0_001011100110;
      patterns[5943] = 29'b0_001011100110_111_0_001011100110;
      patterns[5944] = 29'b0_001011100111_000_0_001011100111;
      patterns[5945] = 29'b0_001011100111_001_0_100111001011;
      patterns[5946] = 29'b0_001011100111_010_0_010111001110;
      patterns[5947] = 29'b0_001011100111_011_0_101110011100;
      patterns[5948] = 29'b0_001011100111_100_1_000101110011;
      patterns[5949] = 29'b0_001011100111_101_1_100010111001;
      patterns[5950] = 29'b0_001011100111_110_0_001011100111;
      patterns[5951] = 29'b0_001011100111_111_0_001011100111;
      patterns[5952] = 29'b0_001011101000_000_0_001011101000;
      patterns[5953] = 29'b0_001011101000_001_0_101000001011;
      patterns[5954] = 29'b0_001011101000_010_0_010111010000;
      patterns[5955] = 29'b0_001011101000_011_0_101110100000;
      patterns[5956] = 29'b0_001011101000_100_0_000101110100;
      patterns[5957] = 29'b0_001011101000_101_0_000010111010;
      patterns[5958] = 29'b0_001011101000_110_0_001011101000;
      patterns[5959] = 29'b0_001011101000_111_0_001011101000;
      patterns[5960] = 29'b0_001011101001_000_0_001011101001;
      patterns[5961] = 29'b0_001011101001_001_0_101001001011;
      patterns[5962] = 29'b0_001011101001_010_0_010111010010;
      patterns[5963] = 29'b0_001011101001_011_0_101110100100;
      patterns[5964] = 29'b0_001011101001_100_1_000101110100;
      patterns[5965] = 29'b0_001011101001_101_0_100010111010;
      patterns[5966] = 29'b0_001011101001_110_0_001011101001;
      patterns[5967] = 29'b0_001011101001_111_0_001011101001;
      patterns[5968] = 29'b0_001011101010_000_0_001011101010;
      patterns[5969] = 29'b0_001011101010_001_0_101010001011;
      patterns[5970] = 29'b0_001011101010_010_0_010111010100;
      patterns[5971] = 29'b0_001011101010_011_0_101110101000;
      patterns[5972] = 29'b0_001011101010_100_0_000101110101;
      patterns[5973] = 29'b0_001011101010_101_1_000010111010;
      patterns[5974] = 29'b0_001011101010_110_0_001011101010;
      patterns[5975] = 29'b0_001011101010_111_0_001011101010;
      patterns[5976] = 29'b0_001011101011_000_0_001011101011;
      patterns[5977] = 29'b0_001011101011_001_0_101011001011;
      patterns[5978] = 29'b0_001011101011_010_0_010111010110;
      patterns[5979] = 29'b0_001011101011_011_0_101110101100;
      patterns[5980] = 29'b0_001011101011_100_1_000101110101;
      patterns[5981] = 29'b0_001011101011_101_1_100010111010;
      patterns[5982] = 29'b0_001011101011_110_0_001011101011;
      patterns[5983] = 29'b0_001011101011_111_0_001011101011;
      patterns[5984] = 29'b0_001011101100_000_0_001011101100;
      patterns[5985] = 29'b0_001011101100_001_0_101100001011;
      patterns[5986] = 29'b0_001011101100_010_0_010111011000;
      patterns[5987] = 29'b0_001011101100_011_0_101110110000;
      patterns[5988] = 29'b0_001011101100_100_0_000101110110;
      patterns[5989] = 29'b0_001011101100_101_0_000010111011;
      patterns[5990] = 29'b0_001011101100_110_0_001011101100;
      patterns[5991] = 29'b0_001011101100_111_0_001011101100;
      patterns[5992] = 29'b0_001011101101_000_0_001011101101;
      patterns[5993] = 29'b0_001011101101_001_0_101101001011;
      patterns[5994] = 29'b0_001011101101_010_0_010111011010;
      patterns[5995] = 29'b0_001011101101_011_0_101110110100;
      patterns[5996] = 29'b0_001011101101_100_1_000101110110;
      patterns[5997] = 29'b0_001011101101_101_0_100010111011;
      patterns[5998] = 29'b0_001011101101_110_0_001011101101;
      patterns[5999] = 29'b0_001011101101_111_0_001011101101;
      patterns[6000] = 29'b0_001011101110_000_0_001011101110;
      patterns[6001] = 29'b0_001011101110_001_0_101110001011;
      patterns[6002] = 29'b0_001011101110_010_0_010111011100;
      patterns[6003] = 29'b0_001011101110_011_0_101110111000;
      patterns[6004] = 29'b0_001011101110_100_0_000101110111;
      patterns[6005] = 29'b0_001011101110_101_1_000010111011;
      patterns[6006] = 29'b0_001011101110_110_0_001011101110;
      patterns[6007] = 29'b0_001011101110_111_0_001011101110;
      patterns[6008] = 29'b0_001011101111_000_0_001011101111;
      patterns[6009] = 29'b0_001011101111_001_0_101111001011;
      patterns[6010] = 29'b0_001011101111_010_0_010111011110;
      patterns[6011] = 29'b0_001011101111_011_0_101110111100;
      patterns[6012] = 29'b0_001011101111_100_1_000101110111;
      patterns[6013] = 29'b0_001011101111_101_1_100010111011;
      patterns[6014] = 29'b0_001011101111_110_0_001011101111;
      patterns[6015] = 29'b0_001011101111_111_0_001011101111;
      patterns[6016] = 29'b0_001011110000_000_0_001011110000;
      patterns[6017] = 29'b0_001011110000_001_0_110000001011;
      patterns[6018] = 29'b0_001011110000_010_0_010111100000;
      patterns[6019] = 29'b0_001011110000_011_0_101111000000;
      patterns[6020] = 29'b0_001011110000_100_0_000101111000;
      patterns[6021] = 29'b0_001011110000_101_0_000010111100;
      patterns[6022] = 29'b0_001011110000_110_0_001011110000;
      patterns[6023] = 29'b0_001011110000_111_0_001011110000;
      patterns[6024] = 29'b0_001011110001_000_0_001011110001;
      patterns[6025] = 29'b0_001011110001_001_0_110001001011;
      patterns[6026] = 29'b0_001011110001_010_0_010111100010;
      patterns[6027] = 29'b0_001011110001_011_0_101111000100;
      patterns[6028] = 29'b0_001011110001_100_1_000101111000;
      patterns[6029] = 29'b0_001011110001_101_0_100010111100;
      patterns[6030] = 29'b0_001011110001_110_0_001011110001;
      patterns[6031] = 29'b0_001011110001_111_0_001011110001;
      patterns[6032] = 29'b0_001011110010_000_0_001011110010;
      patterns[6033] = 29'b0_001011110010_001_0_110010001011;
      patterns[6034] = 29'b0_001011110010_010_0_010111100100;
      patterns[6035] = 29'b0_001011110010_011_0_101111001000;
      patterns[6036] = 29'b0_001011110010_100_0_000101111001;
      patterns[6037] = 29'b0_001011110010_101_1_000010111100;
      patterns[6038] = 29'b0_001011110010_110_0_001011110010;
      patterns[6039] = 29'b0_001011110010_111_0_001011110010;
      patterns[6040] = 29'b0_001011110011_000_0_001011110011;
      patterns[6041] = 29'b0_001011110011_001_0_110011001011;
      patterns[6042] = 29'b0_001011110011_010_0_010111100110;
      patterns[6043] = 29'b0_001011110011_011_0_101111001100;
      patterns[6044] = 29'b0_001011110011_100_1_000101111001;
      patterns[6045] = 29'b0_001011110011_101_1_100010111100;
      patterns[6046] = 29'b0_001011110011_110_0_001011110011;
      patterns[6047] = 29'b0_001011110011_111_0_001011110011;
      patterns[6048] = 29'b0_001011110100_000_0_001011110100;
      patterns[6049] = 29'b0_001011110100_001_0_110100001011;
      patterns[6050] = 29'b0_001011110100_010_0_010111101000;
      patterns[6051] = 29'b0_001011110100_011_0_101111010000;
      patterns[6052] = 29'b0_001011110100_100_0_000101111010;
      patterns[6053] = 29'b0_001011110100_101_0_000010111101;
      patterns[6054] = 29'b0_001011110100_110_0_001011110100;
      patterns[6055] = 29'b0_001011110100_111_0_001011110100;
      patterns[6056] = 29'b0_001011110101_000_0_001011110101;
      patterns[6057] = 29'b0_001011110101_001_0_110101001011;
      patterns[6058] = 29'b0_001011110101_010_0_010111101010;
      patterns[6059] = 29'b0_001011110101_011_0_101111010100;
      patterns[6060] = 29'b0_001011110101_100_1_000101111010;
      patterns[6061] = 29'b0_001011110101_101_0_100010111101;
      patterns[6062] = 29'b0_001011110101_110_0_001011110101;
      patterns[6063] = 29'b0_001011110101_111_0_001011110101;
      patterns[6064] = 29'b0_001011110110_000_0_001011110110;
      patterns[6065] = 29'b0_001011110110_001_0_110110001011;
      patterns[6066] = 29'b0_001011110110_010_0_010111101100;
      patterns[6067] = 29'b0_001011110110_011_0_101111011000;
      patterns[6068] = 29'b0_001011110110_100_0_000101111011;
      patterns[6069] = 29'b0_001011110110_101_1_000010111101;
      patterns[6070] = 29'b0_001011110110_110_0_001011110110;
      patterns[6071] = 29'b0_001011110110_111_0_001011110110;
      patterns[6072] = 29'b0_001011110111_000_0_001011110111;
      patterns[6073] = 29'b0_001011110111_001_0_110111001011;
      patterns[6074] = 29'b0_001011110111_010_0_010111101110;
      patterns[6075] = 29'b0_001011110111_011_0_101111011100;
      patterns[6076] = 29'b0_001011110111_100_1_000101111011;
      patterns[6077] = 29'b0_001011110111_101_1_100010111101;
      patterns[6078] = 29'b0_001011110111_110_0_001011110111;
      patterns[6079] = 29'b0_001011110111_111_0_001011110111;
      patterns[6080] = 29'b0_001011111000_000_0_001011111000;
      patterns[6081] = 29'b0_001011111000_001_0_111000001011;
      patterns[6082] = 29'b0_001011111000_010_0_010111110000;
      patterns[6083] = 29'b0_001011111000_011_0_101111100000;
      patterns[6084] = 29'b0_001011111000_100_0_000101111100;
      patterns[6085] = 29'b0_001011111000_101_0_000010111110;
      patterns[6086] = 29'b0_001011111000_110_0_001011111000;
      patterns[6087] = 29'b0_001011111000_111_0_001011111000;
      patterns[6088] = 29'b0_001011111001_000_0_001011111001;
      patterns[6089] = 29'b0_001011111001_001_0_111001001011;
      patterns[6090] = 29'b0_001011111001_010_0_010111110010;
      patterns[6091] = 29'b0_001011111001_011_0_101111100100;
      patterns[6092] = 29'b0_001011111001_100_1_000101111100;
      patterns[6093] = 29'b0_001011111001_101_0_100010111110;
      patterns[6094] = 29'b0_001011111001_110_0_001011111001;
      patterns[6095] = 29'b0_001011111001_111_0_001011111001;
      patterns[6096] = 29'b0_001011111010_000_0_001011111010;
      patterns[6097] = 29'b0_001011111010_001_0_111010001011;
      patterns[6098] = 29'b0_001011111010_010_0_010111110100;
      patterns[6099] = 29'b0_001011111010_011_0_101111101000;
      patterns[6100] = 29'b0_001011111010_100_0_000101111101;
      patterns[6101] = 29'b0_001011111010_101_1_000010111110;
      patterns[6102] = 29'b0_001011111010_110_0_001011111010;
      patterns[6103] = 29'b0_001011111010_111_0_001011111010;
      patterns[6104] = 29'b0_001011111011_000_0_001011111011;
      patterns[6105] = 29'b0_001011111011_001_0_111011001011;
      patterns[6106] = 29'b0_001011111011_010_0_010111110110;
      patterns[6107] = 29'b0_001011111011_011_0_101111101100;
      patterns[6108] = 29'b0_001011111011_100_1_000101111101;
      patterns[6109] = 29'b0_001011111011_101_1_100010111110;
      patterns[6110] = 29'b0_001011111011_110_0_001011111011;
      patterns[6111] = 29'b0_001011111011_111_0_001011111011;
      patterns[6112] = 29'b0_001011111100_000_0_001011111100;
      patterns[6113] = 29'b0_001011111100_001_0_111100001011;
      patterns[6114] = 29'b0_001011111100_010_0_010111111000;
      patterns[6115] = 29'b0_001011111100_011_0_101111110000;
      patterns[6116] = 29'b0_001011111100_100_0_000101111110;
      patterns[6117] = 29'b0_001011111100_101_0_000010111111;
      patterns[6118] = 29'b0_001011111100_110_0_001011111100;
      patterns[6119] = 29'b0_001011111100_111_0_001011111100;
      patterns[6120] = 29'b0_001011111101_000_0_001011111101;
      patterns[6121] = 29'b0_001011111101_001_0_111101001011;
      patterns[6122] = 29'b0_001011111101_010_0_010111111010;
      patterns[6123] = 29'b0_001011111101_011_0_101111110100;
      patterns[6124] = 29'b0_001011111101_100_1_000101111110;
      patterns[6125] = 29'b0_001011111101_101_0_100010111111;
      patterns[6126] = 29'b0_001011111101_110_0_001011111101;
      patterns[6127] = 29'b0_001011111101_111_0_001011111101;
      patterns[6128] = 29'b0_001011111110_000_0_001011111110;
      patterns[6129] = 29'b0_001011111110_001_0_111110001011;
      patterns[6130] = 29'b0_001011111110_010_0_010111111100;
      patterns[6131] = 29'b0_001011111110_011_0_101111111000;
      patterns[6132] = 29'b0_001011111110_100_0_000101111111;
      patterns[6133] = 29'b0_001011111110_101_1_000010111111;
      patterns[6134] = 29'b0_001011111110_110_0_001011111110;
      patterns[6135] = 29'b0_001011111110_111_0_001011111110;
      patterns[6136] = 29'b0_001011111111_000_0_001011111111;
      patterns[6137] = 29'b0_001011111111_001_0_111111001011;
      patterns[6138] = 29'b0_001011111111_010_0_010111111110;
      patterns[6139] = 29'b0_001011111111_011_0_101111111100;
      patterns[6140] = 29'b0_001011111111_100_1_000101111111;
      patterns[6141] = 29'b0_001011111111_101_1_100010111111;
      patterns[6142] = 29'b0_001011111111_110_0_001011111111;
      patterns[6143] = 29'b0_001011111111_111_0_001011111111;
      patterns[6144] = 29'b0_001100000000_000_0_001100000000;
      patterns[6145] = 29'b0_001100000000_001_0_000000001100;
      patterns[6146] = 29'b0_001100000000_010_0_011000000000;
      patterns[6147] = 29'b0_001100000000_011_0_110000000000;
      patterns[6148] = 29'b0_001100000000_100_0_000110000000;
      patterns[6149] = 29'b0_001100000000_101_0_000011000000;
      patterns[6150] = 29'b0_001100000000_110_0_001100000000;
      patterns[6151] = 29'b0_001100000000_111_0_001100000000;
      patterns[6152] = 29'b0_001100000001_000_0_001100000001;
      patterns[6153] = 29'b0_001100000001_001_0_000001001100;
      patterns[6154] = 29'b0_001100000001_010_0_011000000010;
      patterns[6155] = 29'b0_001100000001_011_0_110000000100;
      patterns[6156] = 29'b0_001100000001_100_1_000110000000;
      patterns[6157] = 29'b0_001100000001_101_0_100011000000;
      patterns[6158] = 29'b0_001100000001_110_0_001100000001;
      patterns[6159] = 29'b0_001100000001_111_0_001100000001;
      patterns[6160] = 29'b0_001100000010_000_0_001100000010;
      patterns[6161] = 29'b0_001100000010_001_0_000010001100;
      patterns[6162] = 29'b0_001100000010_010_0_011000000100;
      patterns[6163] = 29'b0_001100000010_011_0_110000001000;
      patterns[6164] = 29'b0_001100000010_100_0_000110000001;
      patterns[6165] = 29'b0_001100000010_101_1_000011000000;
      patterns[6166] = 29'b0_001100000010_110_0_001100000010;
      patterns[6167] = 29'b0_001100000010_111_0_001100000010;
      patterns[6168] = 29'b0_001100000011_000_0_001100000011;
      patterns[6169] = 29'b0_001100000011_001_0_000011001100;
      patterns[6170] = 29'b0_001100000011_010_0_011000000110;
      patterns[6171] = 29'b0_001100000011_011_0_110000001100;
      patterns[6172] = 29'b0_001100000011_100_1_000110000001;
      patterns[6173] = 29'b0_001100000011_101_1_100011000000;
      patterns[6174] = 29'b0_001100000011_110_0_001100000011;
      patterns[6175] = 29'b0_001100000011_111_0_001100000011;
      patterns[6176] = 29'b0_001100000100_000_0_001100000100;
      patterns[6177] = 29'b0_001100000100_001_0_000100001100;
      patterns[6178] = 29'b0_001100000100_010_0_011000001000;
      patterns[6179] = 29'b0_001100000100_011_0_110000010000;
      patterns[6180] = 29'b0_001100000100_100_0_000110000010;
      patterns[6181] = 29'b0_001100000100_101_0_000011000001;
      patterns[6182] = 29'b0_001100000100_110_0_001100000100;
      patterns[6183] = 29'b0_001100000100_111_0_001100000100;
      patterns[6184] = 29'b0_001100000101_000_0_001100000101;
      patterns[6185] = 29'b0_001100000101_001_0_000101001100;
      patterns[6186] = 29'b0_001100000101_010_0_011000001010;
      patterns[6187] = 29'b0_001100000101_011_0_110000010100;
      patterns[6188] = 29'b0_001100000101_100_1_000110000010;
      patterns[6189] = 29'b0_001100000101_101_0_100011000001;
      patterns[6190] = 29'b0_001100000101_110_0_001100000101;
      patterns[6191] = 29'b0_001100000101_111_0_001100000101;
      patterns[6192] = 29'b0_001100000110_000_0_001100000110;
      patterns[6193] = 29'b0_001100000110_001_0_000110001100;
      patterns[6194] = 29'b0_001100000110_010_0_011000001100;
      patterns[6195] = 29'b0_001100000110_011_0_110000011000;
      patterns[6196] = 29'b0_001100000110_100_0_000110000011;
      patterns[6197] = 29'b0_001100000110_101_1_000011000001;
      patterns[6198] = 29'b0_001100000110_110_0_001100000110;
      patterns[6199] = 29'b0_001100000110_111_0_001100000110;
      patterns[6200] = 29'b0_001100000111_000_0_001100000111;
      patterns[6201] = 29'b0_001100000111_001_0_000111001100;
      patterns[6202] = 29'b0_001100000111_010_0_011000001110;
      patterns[6203] = 29'b0_001100000111_011_0_110000011100;
      patterns[6204] = 29'b0_001100000111_100_1_000110000011;
      patterns[6205] = 29'b0_001100000111_101_1_100011000001;
      patterns[6206] = 29'b0_001100000111_110_0_001100000111;
      patterns[6207] = 29'b0_001100000111_111_0_001100000111;
      patterns[6208] = 29'b0_001100001000_000_0_001100001000;
      patterns[6209] = 29'b0_001100001000_001_0_001000001100;
      patterns[6210] = 29'b0_001100001000_010_0_011000010000;
      patterns[6211] = 29'b0_001100001000_011_0_110000100000;
      patterns[6212] = 29'b0_001100001000_100_0_000110000100;
      patterns[6213] = 29'b0_001100001000_101_0_000011000010;
      patterns[6214] = 29'b0_001100001000_110_0_001100001000;
      patterns[6215] = 29'b0_001100001000_111_0_001100001000;
      patterns[6216] = 29'b0_001100001001_000_0_001100001001;
      patterns[6217] = 29'b0_001100001001_001_0_001001001100;
      patterns[6218] = 29'b0_001100001001_010_0_011000010010;
      patterns[6219] = 29'b0_001100001001_011_0_110000100100;
      patterns[6220] = 29'b0_001100001001_100_1_000110000100;
      patterns[6221] = 29'b0_001100001001_101_0_100011000010;
      patterns[6222] = 29'b0_001100001001_110_0_001100001001;
      patterns[6223] = 29'b0_001100001001_111_0_001100001001;
      patterns[6224] = 29'b0_001100001010_000_0_001100001010;
      patterns[6225] = 29'b0_001100001010_001_0_001010001100;
      patterns[6226] = 29'b0_001100001010_010_0_011000010100;
      patterns[6227] = 29'b0_001100001010_011_0_110000101000;
      patterns[6228] = 29'b0_001100001010_100_0_000110000101;
      patterns[6229] = 29'b0_001100001010_101_1_000011000010;
      patterns[6230] = 29'b0_001100001010_110_0_001100001010;
      patterns[6231] = 29'b0_001100001010_111_0_001100001010;
      patterns[6232] = 29'b0_001100001011_000_0_001100001011;
      patterns[6233] = 29'b0_001100001011_001_0_001011001100;
      patterns[6234] = 29'b0_001100001011_010_0_011000010110;
      patterns[6235] = 29'b0_001100001011_011_0_110000101100;
      patterns[6236] = 29'b0_001100001011_100_1_000110000101;
      patterns[6237] = 29'b0_001100001011_101_1_100011000010;
      patterns[6238] = 29'b0_001100001011_110_0_001100001011;
      patterns[6239] = 29'b0_001100001011_111_0_001100001011;
      patterns[6240] = 29'b0_001100001100_000_0_001100001100;
      patterns[6241] = 29'b0_001100001100_001_0_001100001100;
      patterns[6242] = 29'b0_001100001100_010_0_011000011000;
      patterns[6243] = 29'b0_001100001100_011_0_110000110000;
      patterns[6244] = 29'b0_001100001100_100_0_000110000110;
      patterns[6245] = 29'b0_001100001100_101_0_000011000011;
      patterns[6246] = 29'b0_001100001100_110_0_001100001100;
      patterns[6247] = 29'b0_001100001100_111_0_001100001100;
      patterns[6248] = 29'b0_001100001101_000_0_001100001101;
      patterns[6249] = 29'b0_001100001101_001_0_001101001100;
      patterns[6250] = 29'b0_001100001101_010_0_011000011010;
      patterns[6251] = 29'b0_001100001101_011_0_110000110100;
      patterns[6252] = 29'b0_001100001101_100_1_000110000110;
      patterns[6253] = 29'b0_001100001101_101_0_100011000011;
      patterns[6254] = 29'b0_001100001101_110_0_001100001101;
      patterns[6255] = 29'b0_001100001101_111_0_001100001101;
      patterns[6256] = 29'b0_001100001110_000_0_001100001110;
      patterns[6257] = 29'b0_001100001110_001_0_001110001100;
      patterns[6258] = 29'b0_001100001110_010_0_011000011100;
      patterns[6259] = 29'b0_001100001110_011_0_110000111000;
      patterns[6260] = 29'b0_001100001110_100_0_000110000111;
      patterns[6261] = 29'b0_001100001110_101_1_000011000011;
      patterns[6262] = 29'b0_001100001110_110_0_001100001110;
      patterns[6263] = 29'b0_001100001110_111_0_001100001110;
      patterns[6264] = 29'b0_001100001111_000_0_001100001111;
      patterns[6265] = 29'b0_001100001111_001_0_001111001100;
      patterns[6266] = 29'b0_001100001111_010_0_011000011110;
      patterns[6267] = 29'b0_001100001111_011_0_110000111100;
      patterns[6268] = 29'b0_001100001111_100_1_000110000111;
      patterns[6269] = 29'b0_001100001111_101_1_100011000011;
      patterns[6270] = 29'b0_001100001111_110_0_001100001111;
      patterns[6271] = 29'b0_001100001111_111_0_001100001111;
      patterns[6272] = 29'b0_001100010000_000_0_001100010000;
      patterns[6273] = 29'b0_001100010000_001_0_010000001100;
      patterns[6274] = 29'b0_001100010000_010_0_011000100000;
      patterns[6275] = 29'b0_001100010000_011_0_110001000000;
      patterns[6276] = 29'b0_001100010000_100_0_000110001000;
      patterns[6277] = 29'b0_001100010000_101_0_000011000100;
      patterns[6278] = 29'b0_001100010000_110_0_001100010000;
      patterns[6279] = 29'b0_001100010000_111_0_001100010000;
      patterns[6280] = 29'b0_001100010001_000_0_001100010001;
      patterns[6281] = 29'b0_001100010001_001_0_010001001100;
      patterns[6282] = 29'b0_001100010001_010_0_011000100010;
      patterns[6283] = 29'b0_001100010001_011_0_110001000100;
      patterns[6284] = 29'b0_001100010001_100_1_000110001000;
      patterns[6285] = 29'b0_001100010001_101_0_100011000100;
      patterns[6286] = 29'b0_001100010001_110_0_001100010001;
      patterns[6287] = 29'b0_001100010001_111_0_001100010001;
      patterns[6288] = 29'b0_001100010010_000_0_001100010010;
      patterns[6289] = 29'b0_001100010010_001_0_010010001100;
      patterns[6290] = 29'b0_001100010010_010_0_011000100100;
      patterns[6291] = 29'b0_001100010010_011_0_110001001000;
      patterns[6292] = 29'b0_001100010010_100_0_000110001001;
      patterns[6293] = 29'b0_001100010010_101_1_000011000100;
      patterns[6294] = 29'b0_001100010010_110_0_001100010010;
      patterns[6295] = 29'b0_001100010010_111_0_001100010010;
      patterns[6296] = 29'b0_001100010011_000_0_001100010011;
      patterns[6297] = 29'b0_001100010011_001_0_010011001100;
      patterns[6298] = 29'b0_001100010011_010_0_011000100110;
      patterns[6299] = 29'b0_001100010011_011_0_110001001100;
      patterns[6300] = 29'b0_001100010011_100_1_000110001001;
      patterns[6301] = 29'b0_001100010011_101_1_100011000100;
      patterns[6302] = 29'b0_001100010011_110_0_001100010011;
      patterns[6303] = 29'b0_001100010011_111_0_001100010011;
      patterns[6304] = 29'b0_001100010100_000_0_001100010100;
      patterns[6305] = 29'b0_001100010100_001_0_010100001100;
      patterns[6306] = 29'b0_001100010100_010_0_011000101000;
      patterns[6307] = 29'b0_001100010100_011_0_110001010000;
      patterns[6308] = 29'b0_001100010100_100_0_000110001010;
      patterns[6309] = 29'b0_001100010100_101_0_000011000101;
      patterns[6310] = 29'b0_001100010100_110_0_001100010100;
      patterns[6311] = 29'b0_001100010100_111_0_001100010100;
      patterns[6312] = 29'b0_001100010101_000_0_001100010101;
      patterns[6313] = 29'b0_001100010101_001_0_010101001100;
      patterns[6314] = 29'b0_001100010101_010_0_011000101010;
      patterns[6315] = 29'b0_001100010101_011_0_110001010100;
      patterns[6316] = 29'b0_001100010101_100_1_000110001010;
      patterns[6317] = 29'b0_001100010101_101_0_100011000101;
      patterns[6318] = 29'b0_001100010101_110_0_001100010101;
      patterns[6319] = 29'b0_001100010101_111_0_001100010101;
      patterns[6320] = 29'b0_001100010110_000_0_001100010110;
      patterns[6321] = 29'b0_001100010110_001_0_010110001100;
      patterns[6322] = 29'b0_001100010110_010_0_011000101100;
      patterns[6323] = 29'b0_001100010110_011_0_110001011000;
      patterns[6324] = 29'b0_001100010110_100_0_000110001011;
      patterns[6325] = 29'b0_001100010110_101_1_000011000101;
      patterns[6326] = 29'b0_001100010110_110_0_001100010110;
      patterns[6327] = 29'b0_001100010110_111_0_001100010110;
      patterns[6328] = 29'b0_001100010111_000_0_001100010111;
      patterns[6329] = 29'b0_001100010111_001_0_010111001100;
      patterns[6330] = 29'b0_001100010111_010_0_011000101110;
      patterns[6331] = 29'b0_001100010111_011_0_110001011100;
      patterns[6332] = 29'b0_001100010111_100_1_000110001011;
      patterns[6333] = 29'b0_001100010111_101_1_100011000101;
      patterns[6334] = 29'b0_001100010111_110_0_001100010111;
      patterns[6335] = 29'b0_001100010111_111_0_001100010111;
      patterns[6336] = 29'b0_001100011000_000_0_001100011000;
      patterns[6337] = 29'b0_001100011000_001_0_011000001100;
      patterns[6338] = 29'b0_001100011000_010_0_011000110000;
      patterns[6339] = 29'b0_001100011000_011_0_110001100000;
      patterns[6340] = 29'b0_001100011000_100_0_000110001100;
      patterns[6341] = 29'b0_001100011000_101_0_000011000110;
      patterns[6342] = 29'b0_001100011000_110_0_001100011000;
      patterns[6343] = 29'b0_001100011000_111_0_001100011000;
      patterns[6344] = 29'b0_001100011001_000_0_001100011001;
      patterns[6345] = 29'b0_001100011001_001_0_011001001100;
      patterns[6346] = 29'b0_001100011001_010_0_011000110010;
      patterns[6347] = 29'b0_001100011001_011_0_110001100100;
      patterns[6348] = 29'b0_001100011001_100_1_000110001100;
      patterns[6349] = 29'b0_001100011001_101_0_100011000110;
      patterns[6350] = 29'b0_001100011001_110_0_001100011001;
      patterns[6351] = 29'b0_001100011001_111_0_001100011001;
      patterns[6352] = 29'b0_001100011010_000_0_001100011010;
      patterns[6353] = 29'b0_001100011010_001_0_011010001100;
      patterns[6354] = 29'b0_001100011010_010_0_011000110100;
      patterns[6355] = 29'b0_001100011010_011_0_110001101000;
      patterns[6356] = 29'b0_001100011010_100_0_000110001101;
      patterns[6357] = 29'b0_001100011010_101_1_000011000110;
      patterns[6358] = 29'b0_001100011010_110_0_001100011010;
      patterns[6359] = 29'b0_001100011010_111_0_001100011010;
      patterns[6360] = 29'b0_001100011011_000_0_001100011011;
      patterns[6361] = 29'b0_001100011011_001_0_011011001100;
      patterns[6362] = 29'b0_001100011011_010_0_011000110110;
      patterns[6363] = 29'b0_001100011011_011_0_110001101100;
      patterns[6364] = 29'b0_001100011011_100_1_000110001101;
      patterns[6365] = 29'b0_001100011011_101_1_100011000110;
      patterns[6366] = 29'b0_001100011011_110_0_001100011011;
      patterns[6367] = 29'b0_001100011011_111_0_001100011011;
      patterns[6368] = 29'b0_001100011100_000_0_001100011100;
      patterns[6369] = 29'b0_001100011100_001_0_011100001100;
      patterns[6370] = 29'b0_001100011100_010_0_011000111000;
      patterns[6371] = 29'b0_001100011100_011_0_110001110000;
      patterns[6372] = 29'b0_001100011100_100_0_000110001110;
      patterns[6373] = 29'b0_001100011100_101_0_000011000111;
      patterns[6374] = 29'b0_001100011100_110_0_001100011100;
      patterns[6375] = 29'b0_001100011100_111_0_001100011100;
      patterns[6376] = 29'b0_001100011101_000_0_001100011101;
      patterns[6377] = 29'b0_001100011101_001_0_011101001100;
      patterns[6378] = 29'b0_001100011101_010_0_011000111010;
      patterns[6379] = 29'b0_001100011101_011_0_110001110100;
      patterns[6380] = 29'b0_001100011101_100_1_000110001110;
      patterns[6381] = 29'b0_001100011101_101_0_100011000111;
      patterns[6382] = 29'b0_001100011101_110_0_001100011101;
      patterns[6383] = 29'b0_001100011101_111_0_001100011101;
      patterns[6384] = 29'b0_001100011110_000_0_001100011110;
      patterns[6385] = 29'b0_001100011110_001_0_011110001100;
      patterns[6386] = 29'b0_001100011110_010_0_011000111100;
      patterns[6387] = 29'b0_001100011110_011_0_110001111000;
      patterns[6388] = 29'b0_001100011110_100_0_000110001111;
      patterns[6389] = 29'b0_001100011110_101_1_000011000111;
      patterns[6390] = 29'b0_001100011110_110_0_001100011110;
      patterns[6391] = 29'b0_001100011110_111_0_001100011110;
      patterns[6392] = 29'b0_001100011111_000_0_001100011111;
      patterns[6393] = 29'b0_001100011111_001_0_011111001100;
      patterns[6394] = 29'b0_001100011111_010_0_011000111110;
      patterns[6395] = 29'b0_001100011111_011_0_110001111100;
      patterns[6396] = 29'b0_001100011111_100_1_000110001111;
      patterns[6397] = 29'b0_001100011111_101_1_100011000111;
      patterns[6398] = 29'b0_001100011111_110_0_001100011111;
      patterns[6399] = 29'b0_001100011111_111_0_001100011111;
      patterns[6400] = 29'b0_001100100000_000_0_001100100000;
      patterns[6401] = 29'b0_001100100000_001_0_100000001100;
      patterns[6402] = 29'b0_001100100000_010_0_011001000000;
      patterns[6403] = 29'b0_001100100000_011_0_110010000000;
      patterns[6404] = 29'b0_001100100000_100_0_000110010000;
      patterns[6405] = 29'b0_001100100000_101_0_000011001000;
      patterns[6406] = 29'b0_001100100000_110_0_001100100000;
      patterns[6407] = 29'b0_001100100000_111_0_001100100000;
      patterns[6408] = 29'b0_001100100001_000_0_001100100001;
      patterns[6409] = 29'b0_001100100001_001_0_100001001100;
      patterns[6410] = 29'b0_001100100001_010_0_011001000010;
      patterns[6411] = 29'b0_001100100001_011_0_110010000100;
      patterns[6412] = 29'b0_001100100001_100_1_000110010000;
      patterns[6413] = 29'b0_001100100001_101_0_100011001000;
      patterns[6414] = 29'b0_001100100001_110_0_001100100001;
      patterns[6415] = 29'b0_001100100001_111_0_001100100001;
      patterns[6416] = 29'b0_001100100010_000_0_001100100010;
      patterns[6417] = 29'b0_001100100010_001_0_100010001100;
      patterns[6418] = 29'b0_001100100010_010_0_011001000100;
      patterns[6419] = 29'b0_001100100010_011_0_110010001000;
      patterns[6420] = 29'b0_001100100010_100_0_000110010001;
      patterns[6421] = 29'b0_001100100010_101_1_000011001000;
      patterns[6422] = 29'b0_001100100010_110_0_001100100010;
      patterns[6423] = 29'b0_001100100010_111_0_001100100010;
      patterns[6424] = 29'b0_001100100011_000_0_001100100011;
      patterns[6425] = 29'b0_001100100011_001_0_100011001100;
      patterns[6426] = 29'b0_001100100011_010_0_011001000110;
      patterns[6427] = 29'b0_001100100011_011_0_110010001100;
      patterns[6428] = 29'b0_001100100011_100_1_000110010001;
      patterns[6429] = 29'b0_001100100011_101_1_100011001000;
      patterns[6430] = 29'b0_001100100011_110_0_001100100011;
      patterns[6431] = 29'b0_001100100011_111_0_001100100011;
      patterns[6432] = 29'b0_001100100100_000_0_001100100100;
      patterns[6433] = 29'b0_001100100100_001_0_100100001100;
      patterns[6434] = 29'b0_001100100100_010_0_011001001000;
      patterns[6435] = 29'b0_001100100100_011_0_110010010000;
      patterns[6436] = 29'b0_001100100100_100_0_000110010010;
      patterns[6437] = 29'b0_001100100100_101_0_000011001001;
      patterns[6438] = 29'b0_001100100100_110_0_001100100100;
      patterns[6439] = 29'b0_001100100100_111_0_001100100100;
      patterns[6440] = 29'b0_001100100101_000_0_001100100101;
      patterns[6441] = 29'b0_001100100101_001_0_100101001100;
      patterns[6442] = 29'b0_001100100101_010_0_011001001010;
      patterns[6443] = 29'b0_001100100101_011_0_110010010100;
      patterns[6444] = 29'b0_001100100101_100_1_000110010010;
      patterns[6445] = 29'b0_001100100101_101_0_100011001001;
      patterns[6446] = 29'b0_001100100101_110_0_001100100101;
      patterns[6447] = 29'b0_001100100101_111_0_001100100101;
      patterns[6448] = 29'b0_001100100110_000_0_001100100110;
      patterns[6449] = 29'b0_001100100110_001_0_100110001100;
      patterns[6450] = 29'b0_001100100110_010_0_011001001100;
      patterns[6451] = 29'b0_001100100110_011_0_110010011000;
      patterns[6452] = 29'b0_001100100110_100_0_000110010011;
      patterns[6453] = 29'b0_001100100110_101_1_000011001001;
      patterns[6454] = 29'b0_001100100110_110_0_001100100110;
      patterns[6455] = 29'b0_001100100110_111_0_001100100110;
      patterns[6456] = 29'b0_001100100111_000_0_001100100111;
      patterns[6457] = 29'b0_001100100111_001_0_100111001100;
      patterns[6458] = 29'b0_001100100111_010_0_011001001110;
      patterns[6459] = 29'b0_001100100111_011_0_110010011100;
      patterns[6460] = 29'b0_001100100111_100_1_000110010011;
      patterns[6461] = 29'b0_001100100111_101_1_100011001001;
      patterns[6462] = 29'b0_001100100111_110_0_001100100111;
      patterns[6463] = 29'b0_001100100111_111_0_001100100111;
      patterns[6464] = 29'b0_001100101000_000_0_001100101000;
      patterns[6465] = 29'b0_001100101000_001_0_101000001100;
      patterns[6466] = 29'b0_001100101000_010_0_011001010000;
      patterns[6467] = 29'b0_001100101000_011_0_110010100000;
      patterns[6468] = 29'b0_001100101000_100_0_000110010100;
      patterns[6469] = 29'b0_001100101000_101_0_000011001010;
      patterns[6470] = 29'b0_001100101000_110_0_001100101000;
      patterns[6471] = 29'b0_001100101000_111_0_001100101000;
      patterns[6472] = 29'b0_001100101001_000_0_001100101001;
      patterns[6473] = 29'b0_001100101001_001_0_101001001100;
      patterns[6474] = 29'b0_001100101001_010_0_011001010010;
      patterns[6475] = 29'b0_001100101001_011_0_110010100100;
      patterns[6476] = 29'b0_001100101001_100_1_000110010100;
      patterns[6477] = 29'b0_001100101001_101_0_100011001010;
      patterns[6478] = 29'b0_001100101001_110_0_001100101001;
      patterns[6479] = 29'b0_001100101001_111_0_001100101001;
      patterns[6480] = 29'b0_001100101010_000_0_001100101010;
      patterns[6481] = 29'b0_001100101010_001_0_101010001100;
      patterns[6482] = 29'b0_001100101010_010_0_011001010100;
      patterns[6483] = 29'b0_001100101010_011_0_110010101000;
      patterns[6484] = 29'b0_001100101010_100_0_000110010101;
      patterns[6485] = 29'b0_001100101010_101_1_000011001010;
      patterns[6486] = 29'b0_001100101010_110_0_001100101010;
      patterns[6487] = 29'b0_001100101010_111_0_001100101010;
      patterns[6488] = 29'b0_001100101011_000_0_001100101011;
      patterns[6489] = 29'b0_001100101011_001_0_101011001100;
      patterns[6490] = 29'b0_001100101011_010_0_011001010110;
      patterns[6491] = 29'b0_001100101011_011_0_110010101100;
      patterns[6492] = 29'b0_001100101011_100_1_000110010101;
      patterns[6493] = 29'b0_001100101011_101_1_100011001010;
      patterns[6494] = 29'b0_001100101011_110_0_001100101011;
      patterns[6495] = 29'b0_001100101011_111_0_001100101011;
      patterns[6496] = 29'b0_001100101100_000_0_001100101100;
      patterns[6497] = 29'b0_001100101100_001_0_101100001100;
      patterns[6498] = 29'b0_001100101100_010_0_011001011000;
      patterns[6499] = 29'b0_001100101100_011_0_110010110000;
      patterns[6500] = 29'b0_001100101100_100_0_000110010110;
      patterns[6501] = 29'b0_001100101100_101_0_000011001011;
      patterns[6502] = 29'b0_001100101100_110_0_001100101100;
      patterns[6503] = 29'b0_001100101100_111_0_001100101100;
      patterns[6504] = 29'b0_001100101101_000_0_001100101101;
      patterns[6505] = 29'b0_001100101101_001_0_101101001100;
      patterns[6506] = 29'b0_001100101101_010_0_011001011010;
      patterns[6507] = 29'b0_001100101101_011_0_110010110100;
      patterns[6508] = 29'b0_001100101101_100_1_000110010110;
      patterns[6509] = 29'b0_001100101101_101_0_100011001011;
      patterns[6510] = 29'b0_001100101101_110_0_001100101101;
      patterns[6511] = 29'b0_001100101101_111_0_001100101101;
      patterns[6512] = 29'b0_001100101110_000_0_001100101110;
      patterns[6513] = 29'b0_001100101110_001_0_101110001100;
      patterns[6514] = 29'b0_001100101110_010_0_011001011100;
      patterns[6515] = 29'b0_001100101110_011_0_110010111000;
      patterns[6516] = 29'b0_001100101110_100_0_000110010111;
      patterns[6517] = 29'b0_001100101110_101_1_000011001011;
      patterns[6518] = 29'b0_001100101110_110_0_001100101110;
      patterns[6519] = 29'b0_001100101110_111_0_001100101110;
      patterns[6520] = 29'b0_001100101111_000_0_001100101111;
      patterns[6521] = 29'b0_001100101111_001_0_101111001100;
      patterns[6522] = 29'b0_001100101111_010_0_011001011110;
      patterns[6523] = 29'b0_001100101111_011_0_110010111100;
      patterns[6524] = 29'b0_001100101111_100_1_000110010111;
      patterns[6525] = 29'b0_001100101111_101_1_100011001011;
      patterns[6526] = 29'b0_001100101111_110_0_001100101111;
      patterns[6527] = 29'b0_001100101111_111_0_001100101111;
      patterns[6528] = 29'b0_001100110000_000_0_001100110000;
      patterns[6529] = 29'b0_001100110000_001_0_110000001100;
      patterns[6530] = 29'b0_001100110000_010_0_011001100000;
      patterns[6531] = 29'b0_001100110000_011_0_110011000000;
      patterns[6532] = 29'b0_001100110000_100_0_000110011000;
      patterns[6533] = 29'b0_001100110000_101_0_000011001100;
      patterns[6534] = 29'b0_001100110000_110_0_001100110000;
      patterns[6535] = 29'b0_001100110000_111_0_001100110000;
      patterns[6536] = 29'b0_001100110001_000_0_001100110001;
      patterns[6537] = 29'b0_001100110001_001_0_110001001100;
      patterns[6538] = 29'b0_001100110001_010_0_011001100010;
      patterns[6539] = 29'b0_001100110001_011_0_110011000100;
      patterns[6540] = 29'b0_001100110001_100_1_000110011000;
      patterns[6541] = 29'b0_001100110001_101_0_100011001100;
      patterns[6542] = 29'b0_001100110001_110_0_001100110001;
      patterns[6543] = 29'b0_001100110001_111_0_001100110001;
      patterns[6544] = 29'b0_001100110010_000_0_001100110010;
      patterns[6545] = 29'b0_001100110010_001_0_110010001100;
      patterns[6546] = 29'b0_001100110010_010_0_011001100100;
      patterns[6547] = 29'b0_001100110010_011_0_110011001000;
      patterns[6548] = 29'b0_001100110010_100_0_000110011001;
      patterns[6549] = 29'b0_001100110010_101_1_000011001100;
      patterns[6550] = 29'b0_001100110010_110_0_001100110010;
      patterns[6551] = 29'b0_001100110010_111_0_001100110010;
      patterns[6552] = 29'b0_001100110011_000_0_001100110011;
      patterns[6553] = 29'b0_001100110011_001_0_110011001100;
      patterns[6554] = 29'b0_001100110011_010_0_011001100110;
      patterns[6555] = 29'b0_001100110011_011_0_110011001100;
      patterns[6556] = 29'b0_001100110011_100_1_000110011001;
      patterns[6557] = 29'b0_001100110011_101_1_100011001100;
      patterns[6558] = 29'b0_001100110011_110_0_001100110011;
      patterns[6559] = 29'b0_001100110011_111_0_001100110011;
      patterns[6560] = 29'b0_001100110100_000_0_001100110100;
      patterns[6561] = 29'b0_001100110100_001_0_110100001100;
      patterns[6562] = 29'b0_001100110100_010_0_011001101000;
      patterns[6563] = 29'b0_001100110100_011_0_110011010000;
      patterns[6564] = 29'b0_001100110100_100_0_000110011010;
      patterns[6565] = 29'b0_001100110100_101_0_000011001101;
      patterns[6566] = 29'b0_001100110100_110_0_001100110100;
      patterns[6567] = 29'b0_001100110100_111_0_001100110100;
      patterns[6568] = 29'b0_001100110101_000_0_001100110101;
      patterns[6569] = 29'b0_001100110101_001_0_110101001100;
      patterns[6570] = 29'b0_001100110101_010_0_011001101010;
      patterns[6571] = 29'b0_001100110101_011_0_110011010100;
      patterns[6572] = 29'b0_001100110101_100_1_000110011010;
      patterns[6573] = 29'b0_001100110101_101_0_100011001101;
      patterns[6574] = 29'b0_001100110101_110_0_001100110101;
      patterns[6575] = 29'b0_001100110101_111_0_001100110101;
      patterns[6576] = 29'b0_001100110110_000_0_001100110110;
      patterns[6577] = 29'b0_001100110110_001_0_110110001100;
      patterns[6578] = 29'b0_001100110110_010_0_011001101100;
      patterns[6579] = 29'b0_001100110110_011_0_110011011000;
      patterns[6580] = 29'b0_001100110110_100_0_000110011011;
      patterns[6581] = 29'b0_001100110110_101_1_000011001101;
      patterns[6582] = 29'b0_001100110110_110_0_001100110110;
      patterns[6583] = 29'b0_001100110110_111_0_001100110110;
      patterns[6584] = 29'b0_001100110111_000_0_001100110111;
      patterns[6585] = 29'b0_001100110111_001_0_110111001100;
      patterns[6586] = 29'b0_001100110111_010_0_011001101110;
      patterns[6587] = 29'b0_001100110111_011_0_110011011100;
      patterns[6588] = 29'b0_001100110111_100_1_000110011011;
      patterns[6589] = 29'b0_001100110111_101_1_100011001101;
      patterns[6590] = 29'b0_001100110111_110_0_001100110111;
      patterns[6591] = 29'b0_001100110111_111_0_001100110111;
      patterns[6592] = 29'b0_001100111000_000_0_001100111000;
      patterns[6593] = 29'b0_001100111000_001_0_111000001100;
      patterns[6594] = 29'b0_001100111000_010_0_011001110000;
      patterns[6595] = 29'b0_001100111000_011_0_110011100000;
      patterns[6596] = 29'b0_001100111000_100_0_000110011100;
      patterns[6597] = 29'b0_001100111000_101_0_000011001110;
      patterns[6598] = 29'b0_001100111000_110_0_001100111000;
      patterns[6599] = 29'b0_001100111000_111_0_001100111000;
      patterns[6600] = 29'b0_001100111001_000_0_001100111001;
      patterns[6601] = 29'b0_001100111001_001_0_111001001100;
      patterns[6602] = 29'b0_001100111001_010_0_011001110010;
      patterns[6603] = 29'b0_001100111001_011_0_110011100100;
      patterns[6604] = 29'b0_001100111001_100_1_000110011100;
      patterns[6605] = 29'b0_001100111001_101_0_100011001110;
      patterns[6606] = 29'b0_001100111001_110_0_001100111001;
      patterns[6607] = 29'b0_001100111001_111_0_001100111001;
      patterns[6608] = 29'b0_001100111010_000_0_001100111010;
      patterns[6609] = 29'b0_001100111010_001_0_111010001100;
      patterns[6610] = 29'b0_001100111010_010_0_011001110100;
      patterns[6611] = 29'b0_001100111010_011_0_110011101000;
      patterns[6612] = 29'b0_001100111010_100_0_000110011101;
      patterns[6613] = 29'b0_001100111010_101_1_000011001110;
      patterns[6614] = 29'b0_001100111010_110_0_001100111010;
      patterns[6615] = 29'b0_001100111010_111_0_001100111010;
      patterns[6616] = 29'b0_001100111011_000_0_001100111011;
      patterns[6617] = 29'b0_001100111011_001_0_111011001100;
      patterns[6618] = 29'b0_001100111011_010_0_011001110110;
      patterns[6619] = 29'b0_001100111011_011_0_110011101100;
      patterns[6620] = 29'b0_001100111011_100_1_000110011101;
      patterns[6621] = 29'b0_001100111011_101_1_100011001110;
      patterns[6622] = 29'b0_001100111011_110_0_001100111011;
      patterns[6623] = 29'b0_001100111011_111_0_001100111011;
      patterns[6624] = 29'b0_001100111100_000_0_001100111100;
      patterns[6625] = 29'b0_001100111100_001_0_111100001100;
      patterns[6626] = 29'b0_001100111100_010_0_011001111000;
      patterns[6627] = 29'b0_001100111100_011_0_110011110000;
      patterns[6628] = 29'b0_001100111100_100_0_000110011110;
      patterns[6629] = 29'b0_001100111100_101_0_000011001111;
      patterns[6630] = 29'b0_001100111100_110_0_001100111100;
      patterns[6631] = 29'b0_001100111100_111_0_001100111100;
      patterns[6632] = 29'b0_001100111101_000_0_001100111101;
      patterns[6633] = 29'b0_001100111101_001_0_111101001100;
      patterns[6634] = 29'b0_001100111101_010_0_011001111010;
      patterns[6635] = 29'b0_001100111101_011_0_110011110100;
      patterns[6636] = 29'b0_001100111101_100_1_000110011110;
      patterns[6637] = 29'b0_001100111101_101_0_100011001111;
      patterns[6638] = 29'b0_001100111101_110_0_001100111101;
      patterns[6639] = 29'b0_001100111101_111_0_001100111101;
      patterns[6640] = 29'b0_001100111110_000_0_001100111110;
      patterns[6641] = 29'b0_001100111110_001_0_111110001100;
      patterns[6642] = 29'b0_001100111110_010_0_011001111100;
      patterns[6643] = 29'b0_001100111110_011_0_110011111000;
      patterns[6644] = 29'b0_001100111110_100_0_000110011111;
      patterns[6645] = 29'b0_001100111110_101_1_000011001111;
      patterns[6646] = 29'b0_001100111110_110_0_001100111110;
      patterns[6647] = 29'b0_001100111110_111_0_001100111110;
      patterns[6648] = 29'b0_001100111111_000_0_001100111111;
      patterns[6649] = 29'b0_001100111111_001_0_111111001100;
      patterns[6650] = 29'b0_001100111111_010_0_011001111110;
      patterns[6651] = 29'b0_001100111111_011_0_110011111100;
      patterns[6652] = 29'b0_001100111111_100_1_000110011111;
      patterns[6653] = 29'b0_001100111111_101_1_100011001111;
      patterns[6654] = 29'b0_001100111111_110_0_001100111111;
      patterns[6655] = 29'b0_001100111111_111_0_001100111111;
      patterns[6656] = 29'b0_001101000000_000_0_001101000000;
      patterns[6657] = 29'b0_001101000000_001_0_000000001101;
      patterns[6658] = 29'b0_001101000000_010_0_011010000000;
      patterns[6659] = 29'b0_001101000000_011_0_110100000000;
      patterns[6660] = 29'b0_001101000000_100_0_000110100000;
      patterns[6661] = 29'b0_001101000000_101_0_000011010000;
      patterns[6662] = 29'b0_001101000000_110_0_001101000000;
      patterns[6663] = 29'b0_001101000000_111_0_001101000000;
      patterns[6664] = 29'b0_001101000001_000_0_001101000001;
      patterns[6665] = 29'b0_001101000001_001_0_000001001101;
      patterns[6666] = 29'b0_001101000001_010_0_011010000010;
      patterns[6667] = 29'b0_001101000001_011_0_110100000100;
      patterns[6668] = 29'b0_001101000001_100_1_000110100000;
      patterns[6669] = 29'b0_001101000001_101_0_100011010000;
      patterns[6670] = 29'b0_001101000001_110_0_001101000001;
      patterns[6671] = 29'b0_001101000001_111_0_001101000001;
      patterns[6672] = 29'b0_001101000010_000_0_001101000010;
      patterns[6673] = 29'b0_001101000010_001_0_000010001101;
      patterns[6674] = 29'b0_001101000010_010_0_011010000100;
      patterns[6675] = 29'b0_001101000010_011_0_110100001000;
      patterns[6676] = 29'b0_001101000010_100_0_000110100001;
      patterns[6677] = 29'b0_001101000010_101_1_000011010000;
      patterns[6678] = 29'b0_001101000010_110_0_001101000010;
      patterns[6679] = 29'b0_001101000010_111_0_001101000010;
      patterns[6680] = 29'b0_001101000011_000_0_001101000011;
      patterns[6681] = 29'b0_001101000011_001_0_000011001101;
      patterns[6682] = 29'b0_001101000011_010_0_011010000110;
      patterns[6683] = 29'b0_001101000011_011_0_110100001100;
      patterns[6684] = 29'b0_001101000011_100_1_000110100001;
      patterns[6685] = 29'b0_001101000011_101_1_100011010000;
      patterns[6686] = 29'b0_001101000011_110_0_001101000011;
      patterns[6687] = 29'b0_001101000011_111_0_001101000011;
      patterns[6688] = 29'b0_001101000100_000_0_001101000100;
      patterns[6689] = 29'b0_001101000100_001_0_000100001101;
      patterns[6690] = 29'b0_001101000100_010_0_011010001000;
      patterns[6691] = 29'b0_001101000100_011_0_110100010000;
      patterns[6692] = 29'b0_001101000100_100_0_000110100010;
      patterns[6693] = 29'b0_001101000100_101_0_000011010001;
      patterns[6694] = 29'b0_001101000100_110_0_001101000100;
      patterns[6695] = 29'b0_001101000100_111_0_001101000100;
      patterns[6696] = 29'b0_001101000101_000_0_001101000101;
      patterns[6697] = 29'b0_001101000101_001_0_000101001101;
      patterns[6698] = 29'b0_001101000101_010_0_011010001010;
      patterns[6699] = 29'b0_001101000101_011_0_110100010100;
      patterns[6700] = 29'b0_001101000101_100_1_000110100010;
      patterns[6701] = 29'b0_001101000101_101_0_100011010001;
      patterns[6702] = 29'b0_001101000101_110_0_001101000101;
      patterns[6703] = 29'b0_001101000101_111_0_001101000101;
      patterns[6704] = 29'b0_001101000110_000_0_001101000110;
      patterns[6705] = 29'b0_001101000110_001_0_000110001101;
      patterns[6706] = 29'b0_001101000110_010_0_011010001100;
      patterns[6707] = 29'b0_001101000110_011_0_110100011000;
      patterns[6708] = 29'b0_001101000110_100_0_000110100011;
      patterns[6709] = 29'b0_001101000110_101_1_000011010001;
      patterns[6710] = 29'b0_001101000110_110_0_001101000110;
      patterns[6711] = 29'b0_001101000110_111_0_001101000110;
      patterns[6712] = 29'b0_001101000111_000_0_001101000111;
      patterns[6713] = 29'b0_001101000111_001_0_000111001101;
      patterns[6714] = 29'b0_001101000111_010_0_011010001110;
      patterns[6715] = 29'b0_001101000111_011_0_110100011100;
      patterns[6716] = 29'b0_001101000111_100_1_000110100011;
      patterns[6717] = 29'b0_001101000111_101_1_100011010001;
      patterns[6718] = 29'b0_001101000111_110_0_001101000111;
      patterns[6719] = 29'b0_001101000111_111_0_001101000111;
      patterns[6720] = 29'b0_001101001000_000_0_001101001000;
      patterns[6721] = 29'b0_001101001000_001_0_001000001101;
      patterns[6722] = 29'b0_001101001000_010_0_011010010000;
      patterns[6723] = 29'b0_001101001000_011_0_110100100000;
      patterns[6724] = 29'b0_001101001000_100_0_000110100100;
      patterns[6725] = 29'b0_001101001000_101_0_000011010010;
      patterns[6726] = 29'b0_001101001000_110_0_001101001000;
      patterns[6727] = 29'b0_001101001000_111_0_001101001000;
      patterns[6728] = 29'b0_001101001001_000_0_001101001001;
      patterns[6729] = 29'b0_001101001001_001_0_001001001101;
      patterns[6730] = 29'b0_001101001001_010_0_011010010010;
      patterns[6731] = 29'b0_001101001001_011_0_110100100100;
      patterns[6732] = 29'b0_001101001001_100_1_000110100100;
      patterns[6733] = 29'b0_001101001001_101_0_100011010010;
      patterns[6734] = 29'b0_001101001001_110_0_001101001001;
      patterns[6735] = 29'b0_001101001001_111_0_001101001001;
      patterns[6736] = 29'b0_001101001010_000_0_001101001010;
      patterns[6737] = 29'b0_001101001010_001_0_001010001101;
      patterns[6738] = 29'b0_001101001010_010_0_011010010100;
      patterns[6739] = 29'b0_001101001010_011_0_110100101000;
      patterns[6740] = 29'b0_001101001010_100_0_000110100101;
      patterns[6741] = 29'b0_001101001010_101_1_000011010010;
      patterns[6742] = 29'b0_001101001010_110_0_001101001010;
      patterns[6743] = 29'b0_001101001010_111_0_001101001010;
      patterns[6744] = 29'b0_001101001011_000_0_001101001011;
      patterns[6745] = 29'b0_001101001011_001_0_001011001101;
      patterns[6746] = 29'b0_001101001011_010_0_011010010110;
      patterns[6747] = 29'b0_001101001011_011_0_110100101100;
      patterns[6748] = 29'b0_001101001011_100_1_000110100101;
      patterns[6749] = 29'b0_001101001011_101_1_100011010010;
      patterns[6750] = 29'b0_001101001011_110_0_001101001011;
      patterns[6751] = 29'b0_001101001011_111_0_001101001011;
      patterns[6752] = 29'b0_001101001100_000_0_001101001100;
      patterns[6753] = 29'b0_001101001100_001_0_001100001101;
      patterns[6754] = 29'b0_001101001100_010_0_011010011000;
      patterns[6755] = 29'b0_001101001100_011_0_110100110000;
      patterns[6756] = 29'b0_001101001100_100_0_000110100110;
      patterns[6757] = 29'b0_001101001100_101_0_000011010011;
      patterns[6758] = 29'b0_001101001100_110_0_001101001100;
      patterns[6759] = 29'b0_001101001100_111_0_001101001100;
      patterns[6760] = 29'b0_001101001101_000_0_001101001101;
      patterns[6761] = 29'b0_001101001101_001_0_001101001101;
      patterns[6762] = 29'b0_001101001101_010_0_011010011010;
      patterns[6763] = 29'b0_001101001101_011_0_110100110100;
      patterns[6764] = 29'b0_001101001101_100_1_000110100110;
      patterns[6765] = 29'b0_001101001101_101_0_100011010011;
      patterns[6766] = 29'b0_001101001101_110_0_001101001101;
      patterns[6767] = 29'b0_001101001101_111_0_001101001101;
      patterns[6768] = 29'b0_001101001110_000_0_001101001110;
      patterns[6769] = 29'b0_001101001110_001_0_001110001101;
      patterns[6770] = 29'b0_001101001110_010_0_011010011100;
      patterns[6771] = 29'b0_001101001110_011_0_110100111000;
      patterns[6772] = 29'b0_001101001110_100_0_000110100111;
      patterns[6773] = 29'b0_001101001110_101_1_000011010011;
      patterns[6774] = 29'b0_001101001110_110_0_001101001110;
      patterns[6775] = 29'b0_001101001110_111_0_001101001110;
      patterns[6776] = 29'b0_001101001111_000_0_001101001111;
      patterns[6777] = 29'b0_001101001111_001_0_001111001101;
      patterns[6778] = 29'b0_001101001111_010_0_011010011110;
      patterns[6779] = 29'b0_001101001111_011_0_110100111100;
      patterns[6780] = 29'b0_001101001111_100_1_000110100111;
      patterns[6781] = 29'b0_001101001111_101_1_100011010011;
      patterns[6782] = 29'b0_001101001111_110_0_001101001111;
      patterns[6783] = 29'b0_001101001111_111_0_001101001111;
      patterns[6784] = 29'b0_001101010000_000_0_001101010000;
      patterns[6785] = 29'b0_001101010000_001_0_010000001101;
      patterns[6786] = 29'b0_001101010000_010_0_011010100000;
      patterns[6787] = 29'b0_001101010000_011_0_110101000000;
      patterns[6788] = 29'b0_001101010000_100_0_000110101000;
      patterns[6789] = 29'b0_001101010000_101_0_000011010100;
      patterns[6790] = 29'b0_001101010000_110_0_001101010000;
      patterns[6791] = 29'b0_001101010000_111_0_001101010000;
      patterns[6792] = 29'b0_001101010001_000_0_001101010001;
      patterns[6793] = 29'b0_001101010001_001_0_010001001101;
      patterns[6794] = 29'b0_001101010001_010_0_011010100010;
      patterns[6795] = 29'b0_001101010001_011_0_110101000100;
      patterns[6796] = 29'b0_001101010001_100_1_000110101000;
      patterns[6797] = 29'b0_001101010001_101_0_100011010100;
      patterns[6798] = 29'b0_001101010001_110_0_001101010001;
      patterns[6799] = 29'b0_001101010001_111_0_001101010001;
      patterns[6800] = 29'b0_001101010010_000_0_001101010010;
      patterns[6801] = 29'b0_001101010010_001_0_010010001101;
      patterns[6802] = 29'b0_001101010010_010_0_011010100100;
      patterns[6803] = 29'b0_001101010010_011_0_110101001000;
      patterns[6804] = 29'b0_001101010010_100_0_000110101001;
      patterns[6805] = 29'b0_001101010010_101_1_000011010100;
      patterns[6806] = 29'b0_001101010010_110_0_001101010010;
      patterns[6807] = 29'b0_001101010010_111_0_001101010010;
      patterns[6808] = 29'b0_001101010011_000_0_001101010011;
      patterns[6809] = 29'b0_001101010011_001_0_010011001101;
      patterns[6810] = 29'b0_001101010011_010_0_011010100110;
      patterns[6811] = 29'b0_001101010011_011_0_110101001100;
      patterns[6812] = 29'b0_001101010011_100_1_000110101001;
      patterns[6813] = 29'b0_001101010011_101_1_100011010100;
      patterns[6814] = 29'b0_001101010011_110_0_001101010011;
      patterns[6815] = 29'b0_001101010011_111_0_001101010011;
      patterns[6816] = 29'b0_001101010100_000_0_001101010100;
      patterns[6817] = 29'b0_001101010100_001_0_010100001101;
      patterns[6818] = 29'b0_001101010100_010_0_011010101000;
      patterns[6819] = 29'b0_001101010100_011_0_110101010000;
      patterns[6820] = 29'b0_001101010100_100_0_000110101010;
      patterns[6821] = 29'b0_001101010100_101_0_000011010101;
      patterns[6822] = 29'b0_001101010100_110_0_001101010100;
      patterns[6823] = 29'b0_001101010100_111_0_001101010100;
      patterns[6824] = 29'b0_001101010101_000_0_001101010101;
      patterns[6825] = 29'b0_001101010101_001_0_010101001101;
      patterns[6826] = 29'b0_001101010101_010_0_011010101010;
      patterns[6827] = 29'b0_001101010101_011_0_110101010100;
      patterns[6828] = 29'b0_001101010101_100_1_000110101010;
      patterns[6829] = 29'b0_001101010101_101_0_100011010101;
      patterns[6830] = 29'b0_001101010101_110_0_001101010101;
      patterns[6831] = 29'b0_001101010101_111_0_001101010101;
      patterns[6832] = 29'b0_001101010110_000_0_001101010110;
      patterns[6833] = 29'b0_001101010110_001_0_010110001101;
      patterns[6834] = 29'b0_001101010110_010_0_011010101100;
      patterns[6835] = 29'b0_001101010110_011_0_110101011000;
      patterns[6836] = 29'b0_001101010110_100_0_000110101011;
      patterns[6837] = 29'b0_001101010110_101_1_000011010101;
      patterns[6838] = 29'b0_001101010110_110_0_001101010110;
      patterns[6839] = 29'b0_001101010110_111_0_001101010110;
      patterns[6840] = 29'b0_001101010111_000_0_001101010111;
      patterns[6841] = 29'b0_001101010111_001_0_010111001101;
      patterns[6842] = 29'b0_001101010111_010_0_011010101110;
      patterns[6843] = 29'b0_001101010111_011_0_110101011100;
      patterns[6844] = 29'b0_001101010111_100_1_000110101011;
      patterns[6845] = 29'b0_001101010111_101_1_100011010101;
      patterns[6846] = 29'b0_001101010111_110_0_001101010111;
      patterns[6847] = 29'b0_001101010111_111_0_001101010111;
      patterns[6848] = 29'b0_001101011000_000_0_001101011000;
      patterns[6849] = 29'b0_001101011000_001_0_011000001101;
      patterns[6850] = 29'b0_001101011000_010_0_011010110000;
      patterns[6851] = 29'b0_001101011000_011_0_110101100000;
      patterns[6852] = 29'b0_001101011000_100_0_000110101100;
      patterns[6853] = 29'b0_001101011000_101_0_000011010110;
      patterns[6854] = 29'b0_001101011000_110_0_001101011000;
      patterns[6855] = 29'b0_001101011000_111_0_001101011000;
      patterns[6856] = 29'b0_001101011001_000_0_001101011001;
      patterns[6857] = 29'b0_001101011001_001_0_011001001101;
      patterns[6858] = 29'b0_001101011001_010_0_011010110010;
      patterns[6859] = 29'b0_001101011001_011_0_110101100100;
      patterns[6860] = 29'b0_001101011001_100_1_000110101100;
      patterns[6861] = 29'b0_001101011001_101_0_100011010110;
      patterns[6862] = 29'b0_001101011001_110_0_001101011001;
      patterns[6863] = 29'b0_001101011001_111_0_001101011001;
      patterns[6864] = 29'b0_001101011010_000_0_001101011010;
      patterns[6865] = 29'b0_001101011010_001_0_011010001101;
      patterns[6866] = 29'b0_001101011010_010_0_011010110100;
      patterns[6867] = 29'b0_001101011010_011_0_110101101000;
      patterns[6868] = 29'b0_001101011010_100_0_000110101101;
      patterns[6869] = 29'b0_001101011010_101_1_000011010110;
      patterns[6870] = 29'b0_001101011010_110_0_001101011010;
      patterns[6871] = 29'b0_001101011010_111_0_001101011010;
      patterns[6872] = 29'b0_001101011011_000_0_001101011011;
      patterns[6873] = 29'b0_001101011011_001_0_011011001101;
      patterns[6874] = 29'b0_001101011011_010_0_011010110110;
      patterns[6875] = 29'b0_001101011011_011_0_110101101100;
      patterns[6876] = 29'b0_001101011011_100_1_000110101101;
      patterns[6877] = 29'b0_001101011011_101_1_100011010110;
      patterns[6878] = 29'b0_001101011011_110_0_001101011011;
      patterns[6879] = 29'b0_001101011011_111_0_001101011011;
      patterns[6880] = 29'b0_001101011100_000_0_001101011100;
      patterns[6881] = 29'b0_001101011100_001_0_011100001101;
      patterns[6882] = 29'b0_001101011100_010_0_011010111000;
      patterns[6883] = 29'b0_001101011100_011_0_110101110000;
      patterns[6884] = 29'b0_001101011100_100_0_000110101110;
      patterns[6885] = 29'b0_001101011100_101_0_000011010111;
      patterns[6886] = 29'b0_001101011100_110_0_001101011100;
      patterns[6887] = 29'b0_001101011100_111_0_001101011100;
      patterns[6888] = 29'b0_001101011101_000_0_001101011101;
      patterns[6889] = 29'b0_001101011101_001_0_011101001101;
      patterns[6890] = 29'b0_001101011101_010_0_011010111010;
      patterns[6891] = 29'b0_001101011101_011_0_110101110100;
      patterns[6892] = 29'b0_001101011101_100_1_000110101110;
      patterns[6893] = 29'b0_001101011101_101_0_100011010111;
      patterns[6894] = 29'b0_001101011101_110_0_001101011101;
      patterns[6895] = 29'b0_001101011101_111_0_001101011101;
      patterns[6896] = 29'b0_001101011110_000_0_001101011110;
      patterns[6897] = 29'b0_001101011110_001_0_011110001101;
      patterns[6898] = 29'b0_001101011110_010_0_011010111100;
      patterns[6899] = 29'b0_001101011110_011_0_110101111000;
      patterns[6900] = 29'b0_001101011110_100_0_000110101111;
      patterns[6901] = 29'b0_001101011110_101_1_000011010111;
      patterns[6902] = 29'b0_001101011110_110_0_001101011110;
      patterns[6903] = 29'b0_001101011110_111_0_001101011110;
      patterns[6904] = 29'b0_001101011111_000_0_001101011111;
      patterns[6905] = 29'b0_001101011111_001_0_011111001101;
      patterns[6906] = 29'b0_001101011111_010_0_011010111110;
      patterns[6907] = 29'b0_001101011111_011_0_110101111100;
      patterns[6908] = 29'b0_001101011111_100_1_000110101111;
      patterns[6909] = 29'b0_001101011111_101_1_100011010111;
      patterns[6910] = 29'b0_001101011111_110_0_001101011111;
      patterns[6911] = 29'b0_001101011111_111_0_001101011111;
      patterns[6912] = 29'b0_001101100000_000_0_001101100000;
      patterns[6913] = 29'b0_001101100000_001_0_100000001101;
      patterns[6914] = 29'b0_001101100000_010_0_011011000000;
      patterns[6915] = 29'b0_001101100000_011_0_110110000000;
      patterns[6916] = 29'b0_001101100000_100_0_000110110000;
      patterns[6917] = 29'b0_001101100000_101_0_000011011000;
      patterns[6918] = 29'b0_001101100000_110_0_001101100000;
      patterns[6919] = 29'b0_001101100000_111_0_001101100000;
      patterns[6920] = 29'b0_001101100001_000_0_001101100001;
      patterns[6921] = 29'b0_001101100001_001_0_100001001101;
      patterns[6922] = 29'b0_001101100001_010_0_011011000010;
      patterns[6923] = 29'b0_001101100001_011_0_110110000100;
      patterns[6924] = 29'b0_001101100001_100_1_000110110000;
      patterns[6925] = 29'b0_001101100001_101_0_100011011000;
      patterns[6926] = 29'b0_001101100001_110_0_001101100001;
      patterns[6927] = 29'b0_001101100001_111_0_001101100001;
      patterns[6928] = 29'b0_001101100010_000_0_001101100010;
      patterns[6929] = 29'b0_001101100010_001_0_100010001101;
      patterns[6930] = 29'b0_001101100010_010_0_011011000100;
      patterns[6931] = 29'b0_001101100010_011_0_110110001000;
      patterns[6932] = 29'b0_001101100010_100_0_000110110001;
      patterns[6933] = 29'b0_001101100010_101_1_000011011000;
      patterns[6934] = 29'b0_001101100010_110_0_001101100010;
      patterns[6935] = 29'b0_001101100010_111_0_001101100010;
      patterns[6936] = 29'b0_001101100011_000_0_001101100011;
      patterns[6937] = 29'b0_001101100011_001_0_100011001101;
      patterns[6938] = 29'b0_001101100011_010_0_011011000110;
      patterns[6939] = 29'b0_001101100011_011_0_110110001100;
      patterns[6940] = 29'b0_001101100011_100_1_000110110001;
      patterns[6941] = 29'b0_001101100011_101_1_100011011000;
      patterns[6942] = 29'b0_001101100011_110_0_001101100011;
      patterns[6943] = 29'b0_001101100011_111_0_001101100011;
      patterns[6944] = 29'b0_001101100100_000_0_001101100100;
      patterns[6945] = 29'b0_001101100100_001_0_100100001101;
      patterns[6946] = 29'b0_001101100100_010_0_011011001000;
      patterns[6947] = 29'b0_001101100100_011_0_110110010000;
      patterns[6948] = 29'b0_001101100100_100_0_000110110010;
      patterns[6949] = 29'b0_001101100100_101_0_000011011001;
      patterns[6950] = 29'b0_001101100100_110_0_001101100100;
      patterns[6951] = 29'b0_001101100100_111_0_001101100100;
      patterns[6952] = 29'b0_001101100101_000_0_001101100101;
      patterns[6953] = 29'b0_001101100101_001_0_100101001101;
      patterns[6954] = 29'b0_001101100101_010_0_011011001010;
      patterns[6955] = 29'b0_001101100101_011_0_110110010100;
      patterns[6956] = 29'b0_001101100101_100_1_000110110010;
      patterns[6957] = 29'b0_001101100101_101_0_100011011001;
      patterns[6958] = 29'b0_001101100101_110_0_001101100101;
      patterns[6959] = 29'b0_001101100101_111_0_001101100101;
      patterns[6960] = 29'b0_001101100110_000_0_001101100110;
      patterns[6961] = 29'b0_001101100110_001_0_100110001101;
      patterns[6962] = 29'b0_001101100110_010_0_011011001100;
      patterns[6963] = 29'b0_001101100110_011_0_110110011000;
      patterns[6964] = 29'b0_001101100110_100_0_000110110011;
      patterns[6965] = 29'b0_001101100110_101_1_000011011001;
      patterns[6966] = 29'b0_001101100110_110_0_001101100110;
      patterns[6967] = 29'b0_001101100110_111_0_001101100110;
      patterns[6968] = 29'b0_001101100111_000_0_001101100111;
      patterns[6969] = 29'b0_001101100111_001_0_100111001101;
      patterns[6970] = 29'b0_001101100111_010_0_011011001110;
      patterns[6971] = 29'b0_001101100111_011_0_110110011100;
      patterns[6972] = 29'b0_001101100111_100_1_000110110011;
      patterns[6973] = 29'b0_001101100111_101_1_100011011001;
      patterns[6974] = 29'b0_001101100111_110_0_001101100111;
      patterns[6975] = 29'b0_001101100111_111_0_001101100111;
      patterns[6976] = 29'b0_001101101000_000_0_001101101000;
      patterns[6977] = 29'b0_001101101000_001_0_101000001101;
      patterns[6978] = 29'b0_001101101000_010_0_011011010000;
      patterns[6979] = 29'b0_001101101000_011_0_110110100000;
      patterns[6980] = 29'b0_001101101000_100_0_000110110100;
      patterns[6981] = 29'b0_001101101000_101_0_000011011010;
      patterns[6982] = 29'b0_001101101000_110_0_001101101000;
      patterns[6983] = 29'b0_001101101000_111_0_001101101000;
      patterns[6984] = 29'b0_001101101001_000_0_001101101001;
      patterns[6985] = 29'b0_001101101001_001_0_101001001101;
      patterns[6986] = 29'b0_001101101001_010_0_011011010010;
      patterns[6987] = 29'b0_001101101001_011_0_110110100100;
      patterns[6988] = 29'b0_001101101001_100_1_000110110100;
      patterns[6989] = 29'b0_001101101001_101_0_100011011010;
      patterns[6990] = 29'b0_001101101001_110_0_001101101001;
      patterns[6991] = 29'b0_001101101001_111_0_001101101001;
      patterns[6992] = 29'b0_001101101010_000_0_001101101010;
      patterns[6993] = 29'b0_001101101010_001_0_101010001101;
      patterns[6994] = 29'b0_001101101010_010_0_011011010100;
      patterns[6995] = 29'b0_001101101010_011_0_110110101000;
      patterns[6996] = 29'b0_001101101010_100_0_000110110101;
      patterns[6997] = 29'b0_001101101010_101_1_000011011010;
      patterns[6998] = 29'b0_001101101010_110_0_001101101010;
      patterns[6999] = 29'b0_001101101010_111_0_001101101010;
      patterns[7000] = 29'b0_001101101011_000_0_001101101011;
      patterns[7001] = 29'b0_001101101011_001_0_101011001101;
      patterns[7002] = 29'b0_001101101011_010_0_011011010110;
      patterns[7003] = 29'b0_001101101011_011_0_110110101100;
      patterns[7004] = 29'b0_001101101011_100_1_000110110101;
      patterns[7005] = 29'b0_001101101011_101_1_100011011010;
      patterns[7006] = 29'b0_001101101011_110_0_001101101011;
      patterns[7007] = 29'b0_001101101011_111_0_001101101011;
      patterns[7008] = 29'b0_001101101100_000_0_001101101100;
      patterns[7009] = 29'b0_001101101100_001_0_101100001101;
      patterns[7010] = 29'b0_001101101100_010_0_011011011000;
      patterns[7011] = 29'b0_001101101100_011_0_110110110000;
      patterns[7012] = 29'b0_001101101100_100_0_000110110110;
      patterns[7013] = 29'b0_001101101100_101_0_000011011011;
      patterns[7014] = 29'b0_001101101100_110_0_001101101100;
      patterns[7015] = 29'b0_001101101100_111_0_001101101100;
      patterns[7016] = 29'b0_001101101101_000_0_001101101101;
      patterns[7017] = 29'b0_001101101101_001_0_101101001101;
      patterns[7018] = 29'b0_001101101101_010_0_011011011010;
      patterns[7019] = 29'b0_001101101101_011_0_110110110100;
      patterns[7020] = 29'b0_001101101101_100_1_000110110110;
      patterns[7021] = 29'b0_001101101101_101_0_100011011011;
      patterns[7022] = 29'b0_001101101101_110_0_001101101101;
      patterns[7023] = 29'b0_001101101101_111_0_001101101101;
      patterns[7024] = 29'b0_001101101110_000_0_001101101110;
      patterns[7025] = 29'b0_001101101110_001_0_101110001101;
      patterns[7026] = 29'b0_001101101110_010_0_011011011100;
      patterns[7027] = 29'b0_001101101110_011_0_110110111000;
      patterns[7028] = 29'b0_001101101110_100_0_000110110111;
      patterns[7029] = 29'b0_001101101110_101_1_000011011011;
      patterns[7030] = 29'b0_001101101110_110_0_001101101110;
      patterns[7031] = 29'b0_001101101110_111_0_001101101110;
      patterns[7032] = 29'b0_001101101111_000_0_001101101111;
      patterns[7033] = 29'b0_001101101111_001_0_101111001101;
      patterns[7034] = 29'b0_001101101111_010_0_011011011110;
      patterns[7035] = 29'b0_001101101111_011_0_110110111100;
      patterns[7036] = 29'b0_001101101111_100_1_000110110111;
      patterns[7037] = 29'b0_001101101111_101_1_100011011011;
      patterns[7038] = 29'b0_001101101111_110_0_001101101111;
      patterns[7039] = 29'b0_001101101111_111_0_001101101111;
      patterns[7040] = 29'b0_001101110000_000_0_001101110000;
      patterns[7041] = 29'b0_001101110000_001_0_110000001101;
      patterns[7042] = 29'b0_001101110000_010_0_011011100000;
      patterns[7043] = 29'b0_001101110000_011_0_110111000000;
      patterns[7044] = 29'b0_001101110000_100_0_000110111000;
      patterns[7045] = 29'b0_001101110000_101_0_000011011100;
      patterns[7046] = 29'b0_001101110000_110_0_001101110000;
      patterns[7047] = 29'b0_001101110000_111_0_001101110000;
      patterns[7048] = 29'b0_001101110001_000_0_001101110001;
      patterns[7049] = 29'b0_001101110001_001_0_110001001101;
      patterns[7050] = 29'b0_001101110001_010_0_011011100010;
      patterns[7051] = 29'b0_001101110001_011_0_110111000100;
      patterns[7052] = 29'b0_001101110001_100_1_000110111000;
      patterns[7053] = 29'b0_001101110001_101_0_100011011100;
      patterns[7054] = 29'b0_001101110001_110_0_001101110001;
      patterns[7055] = 29'b0_001101110001_111_0_001101110001;
      patterns[7056] = 29'b0_001101110010_000_0_001101110010;
      patterns[7057] = 29'b0_001101110010_001_0_110010001101;
      patterns[7058] = 29'b0_001101110010_010_0_011011100100;
      patterns[7059] = 29'b0_001101110010_011_0_110111001000;
      patterns[7060] = 29'b0_001101110010_100_0_000110111001;
      patterns[7061] = 29'b0_001101110010_101_1_000011011100;
      patterns[7062] = 29'b0_001101110010_110_0_001101110010;
      patterns[7063] = 29'b0_001101110010_111_0_001101110010;
      patterns[7064] = 29'b0_001101110011_000_0_001101110011;
      patterns[7065] = 29'b0_001101110011_001_0_110011001101;
      patterns[7066] = 29'b0_001101110011_010_0_011011100110;
      patterns[7067] = 29'b0_001101110011_011_0_110111001100;
      patterns[7068] = 29'b0_001101110011_100_1_000110111001;
      patterns[7069] = 29'b0_001101110011_101_1_100011011100;
      patterns[7070] = 29'b0_001101110011_110_0_001101110011;
      patterns[7071] = 29'b0_001101110011_111_0_001101110011;
      patterns[7072] = 29'b0_001101110100_000_0_001101110100;
      patterns[7073] = 29'b0_001101110100_001_0_110100001101;
      patterns[7074] = 29'b0_001101110100_010_0_011011101000;
      patterns[7075] = 29'b0_001101110100_011_0_110111010000;
      patterns[7076] = 29'b0_001101110100_100_0_000110111010;
      patterns[7077] = 29'b0_001101110100_101_0_000011011101;
      patterns[7078] = 29'b0_001101110100_110_0_001101110100;
      patterns[7079] = 29'b0_001101110100_111_0_001101110100;
      patterns[7080] = 29'b0_001101110101_000_0_001101110101;
      patterns[7081] = 29'b0_001101110101_001_0_110101001101;
      patterns[7082] = 29'b0_001101110101_010_0_011011101010;
      patterns[7083] = 29'b0_001101110101_011_0_110111010100;
      patterns[7084] = 29'b0_001101110101_100_1_000110111010;
      patterns[7085] = 29'b0_001101110101_101_0_100011011101;
      patterns[7086] = 29'b0_001101110101_110_0_001101110101;
      patterns[7087] = 29'b0_001101110101_111_0_001101110101;
      patterns[7088] = 29'b0_001101110110_000_0_001101110110;
      patterns[7089] = 29'b0_001101110110_001_0_110110001101;
      patterns[7090] = 29'b0_001101110110_010_0_011011101100;
      patterns[7091] = 29'b0_001101110110_011_0_110111011000;
      patterns[7092] = 29'b0_001101110110_100_0_000110111011;
      patterns[7093] = 29'b0_001101110110_101_1_000011011101;
      patterns[7094] = 29'b0_001101110110_110_0_001101110110;
      patterns[7095] = 29'b0_001101110110_111_0_001101110110;
      patterns[7096] = 29'b0_001101110111_000_0_001101110111;
      patterns[7097] = 29'b0_001101110111_001_0_110111001101;
      patterns[7098] = 29'b0_001101110111_010_0_011011101110;
      patterns[7099] = 29'b0_001101110111_011_0_110111011100;
      patterns[7100] = 29'b0_001101110111_100_1_000110111011;
      patterns[7101] = 29'b0_001101110111_101_1_100011011101;
      patterns[7102] = 29'b0_001101110111_110_0_001101110111;
      patterns[7103] = 29'b0_001101110111_111_0_001101110111;
      patterns[7104] = 29'b0_001101111000_000_0_001101111000;
      patterns[7105] = 29'b0_001101111000_001_0_111000001101;
      patterns[7106] = 29'b0_001101111000_010_0_011011110000;
      patterns[7107] = 29'b0_001101111000_011_0_110111100000;
      patterns[7108] = 29'b0_001101111000_100_0_000110111100;
      patterns[7109] = 29'b0_001101111000_101_0_000011011110;
      patterns[7110] = 29'b0_001101111000_110_0_001101111000;
      patterns[7111] = 29'b0_001101111000_111_0_001101111000;
      patterns[7112] = 29'b0_001101111001_000_0_001101111001;
      patterns[7113] = 29'b0_001101111001_001_0_111001001101;
      patterns[7114] = 29'b0_001101111001_010_0_011011110010;
      patterns[7115] = 29'b0_001101111001_011_0_110111100100;
      patterns[7116] = 29'b0_001101111001_100_1_000110111100;
      patterns[7117] = 29'b0_001101111001_101_0_100011011110;
      patterns[7118] = 29'b0_001101111001_110_0_001101111001;
      patterns[7119] = 29'b0_001101111001_111_0_001101111001;
      patterns[7120] = 29'b0_001101111010_000_0_001101111010;
      patterns[7121] = 29'b0_001101111010_001_0_111010001101;
      patterns[7122] = 29'b0_001101111010_010_0_011011110100;
      patterns[7123] = 29'b0_001101111010_011_0_110111101000;
      patterns[7124] = 29'b0_001101111010_100_0_000110111101;
      patterns[7125] = 29'b0_001101111010_101_1_000011011110;
      patterns[7126] = 29'b0_001101111010_110_0_001101111010;
      patterns[7127] = 29'b0_001101111010_111_0_001101111010;
      patterns[7128] = 29'b0_001101111011_000_0_001101111011;
      patterns[7129] = 29'b0_001101111011_001_0_111011001101;
      patterns[7130] = 29'b0_001101111011_010_0_011011110110;
      patterns[7131] = 29'b0_001101111011_011_0_110111101100;
      patterns[7132] = 29'b0_001101111011_100_1_000110111101;
      patterns[7133] = 29'b0_001101111011_101_1_100011011110;
      patterns[7134] = 29'b0_001101111011_110_0_001101111011;
      patterns[7135] = 29'b0_001101111011_111_0_001101111011;
      patterns[7136] = 29'b0_001101111100_000_0_001101111100;
      patterns[7137] = 29'b0_001101111100_001_0_111100001101;
      patterns[7138] = 29'b0_001101111100_010_0_011011111000;
      patterns[7139] = 29'b0_001101111100_011_0_110111110000;
      patterns[7140] = 29'b0_001101111100_100_0_000110111110;
      patterns[7141] = 29'b0_001101111100_101_0_000011011111;
      patterns[7142] = 29'b0_001101111100_110_0_001101111100;
      patterns[7143] = 29'b0_001101111100_111_0_001101111100;
      patterns[7144] = 29'b0_001101111101_000_0_001101111101;
      patterns[7145] = 29'b0_001101111101_001_0_111101001101;
      patterns[7146] = 29'b0_001101111101_010_0_011011111010;
      patterns[7147] = 29'b0_001101111101_011_0_110111110100;
      patterns[7148] = 29'b0_001101111101_100_1_000110111110;
      patterns[7149] = 29'b0_001101111101_101_0_100011011111;
      patterns[7150] = 29'b0_001101111101_110_0_001101111101;
      patterns[7151] = 29'b0_001101111101_111_0_001101111101;
      patterns[7152] = 29'b0_001101111110_000_0_001101111110;
      patterns[7153] = 29'b0_001101111110_001_0_111110001101;
      patterns[7154] = 29'b0_001101111110_010_0_011011111100;
      patterns[7155] = 29'b0_001101111110_011_0_110111111000;
      patterns[7156] = 29'b0_001101111110_100_0_000110111111;
      patterns[7157] = 29'b0_001101111110_101_1_000011011111;
      patterns[7158] = 29'b0_001101111110_110_0_001101111110;
      patterns[7159] = 29'b0_001101111110_111_0_001101111110;
      patterns[7160] = 29'b0_001101111111_000_0_001101111111;
      patterns[7161] = 29'b0_001101111111_001_0_111111001101;
      patterns[7162] = 29'b0_001101111111_010_0_011011111110;
      patterns[7163] = 29'b0_001101111111_011_0_110111111100;
      patterns[7164] = 29'b0_001101111111_100_1_000110111111;
      patterns[7165] = 29'b0_001101111111_101_1_100011011111;
      patterns[7166] = 29'b0_001101111111_110_0_001101111111;
      patterns[7167] = 29'b0_001101111111_111_0_001101111111;
      patterns[7168] = 29'b0_001110000000_000_0_001110000000;
      patterns[7169] = 29'b0_001110000000_001_0_000000001110;
      patterns[7170] = 29'b0_001110000000_010_0_011100000000;
      patterns[7171] = 29'b0_001110000000_011_0_111000000000;
      patterns[7172] = 29'b0_001110000000_100_0_000111000000;
      patterns[7173] = 29'b0_001110000000_101_0_000011100000;
      patterns[7174] = 29'b0_001110000000_110_0_001110000000;
      patterns[7175] = 29'b0_001110000000_111_0_001110000000;
      patterns[7176] = 29'b0_001110000001_000_0_001110000001;
      patterns[7177] = 29'b0_001110000001_001_0_000001001110;
      patterns[7178] = 29'b0_001110000001_010_0_011100000010;
      patterns[7179] = 29'b0_001110000001_011_0_111000000100;
      patterns[7180] = 29'b0_001110000001_100_1_000111000000;
      patterns[7181] = 29'b0_001110000001_101_0_100011100000;
      patterns[7182] = 29'b0_001110000001_110_0_001110000001;
      patterns[7183] = 29'b0_001110000001_111_0_001110000001;
      patterns[7184] = 29'b0_001110000010_000_0_001110000010;
      patterns[7185] = 29'b0_001110000010_001_0_000010001110;
      patterns[7186] = 29'b0_001110000010_010_0_011100000100;
      patterns[7187] = 29'b0_001110000010_011_0_111000001000;
      patterns[7188] = 29'b0_001110000010_100_0_000111000001;
      patterns[7189] = 29'b0_001110000010_101_1_000011100000;
      patterns[7190] = 29'b0_001110000010_110_0_001110000010;
      patterns[7191] = 29'b0_001110000010_111_0_001110000010;
      patterns[7192] = 29'b0_001110000011_000_0_001110000011;
      patterns[7193] = 29'b0_001110000011_001_0_000011001110;
      patterns[7194] = 29'b0_001110000011_010_0_011100000110;
      patterns[7195] = 29'b0_001110000011_011_0_111000001100;
      patterns[7196] = 29'b0_001110000011_100_1_000111000001;
      patterns[7197] = 29'b0_001110000011_101_1_100011100000;
      patterns[7198] = 29'b0_001110000011_110_0_001110000011;
      patterns[7199] = 29'b0_001110000011_111_0_001110000011;
      patterns[7200] = 29'b0_001110000100_000_0_001110000100;
      patterns[7201] = 29'b0_001110000100_001_0_000100001110;
      patterns[7202] = 29'b0_001110000100_010_0_011100001000;
      patterns[7203] = 29'b0_001110000100_011_0_111000010000;
      patterns[7204] = 29'b0_001110000100_100_0_000111000010;
      patterns[7205] = 29'b0_001110000100_101_0_000011100001;
      patterns[7206] = 29'b0_001110000100_110_0_001110000100;
      patterns[7207] = 29'b0_001110000100_111_0_001110000100;
      patterns[7208] = 29'b0_001110000101_000_0_001110000101;
      patterns[7209] = 29'b0_001110000101_001_0_000101001110;
      patterns[7210] = 29'b0_001110000101_010_0_011100001010;
      patterns[7211] = 29'b0_001110000101_011_0_111000010100;
      patterns[7212] = 29'b0_001110000101_100_1_000111000010;
      patterns[7213] = 29'b0_001110000101_101_0_100011100001;
      patterns[7214] = 29'b0_001110000101_110_0_001110000101;
      patterns[7215] = 29'b0_001110000101_111_0_001110000101;
      patterns[7216] = 29'b0_001110000110_000_0_001110000110;
      patterns[7217] = 29'b0_001110000110_001_0_000110001110;
      patterns[7218] = 29'b0_001110000110_010_0_011100001100;
      patterns[7219] = 29'b0_001110000110_011_0_111000011000;
      patterns[7220] = 29'b0_001110000110_100_0_000111000011;
      patterns[7221] = 29'b0_001110000110_101_1_000011100001;
      patterns[7222] = 29'b0_001110000110_110_0_001110000110;
      patterns[7223] = 29'b0_001110000110_111_0_001110000110;
      patterns[7224] = 29'b0_001110000111_000_0_001110000111;
      patterns[7225] = 29'b0_001110000111_001_0_000111001110;
      patterns[7226] = 29'b0_001110000111_010_0_011100001110;
      patterns[7227] = 29'b0_001110000111_011_0_111000011100;
      patterns[7228] = 29'b0_001110000111_100_1_000111000011;
      patterns[7229] = 29'b0_001110000111_101_1_100011100001;
      patterns[7230] = 29'b0_001110000111_110_0_001110000111;
      patterns[7231] = 29'b0_001110000111_111_0_001110000111;
      patterns[7232] = 29'b0_001110001000_000_0_001110001000;
      patterns[7233] = 29'b0_001110001000_001_0_001000001110;
      patterns[7234] = 29'b0_001110001000_010_0_011100010000;
      patterns[7235] = 29'b0_001110001000_011_0_111000100000;
      patterns[7236] = 29'b0_001110001000_100_0_000111000100;
      patterns[7237] = 29'b0_001110001000_101_0_000011100010;
      patterns[7238] = 29'b0_001110001000_110_0_001110001000;
      patterns[7239] = 29'b0_001110001000_111_0_001110001000;
      patterns[7240] = 29'b0_001110001001_000_0_001110001001;
      patterns[7241] = 29'b0_001110001001_001_0_001001001110;
      patterns[7242] = 29'b0_001110001001_010_0_011100010010;
      patterns[7243] = 29'b0_001110001001_011_0_111000100100;
      patterns[7244] = 29'b0_001110001001_100_1_000111000100;
      patterns[7245] = 29'b0_001110001001_101_0_100011100010;
      patterns[7246] = 29'b0_001110001001_110_0_001110001001;
      patterns[7247] = 29'b0_001110001001_111_0_001110001001;
      patterns[7248] = 29'b0_001110001010_000_0_001110001010;
      patterns[7249] = 29'b0_001110001010_001_0_001010001110;
      patterns[7250] = 29'b0_001110001010_010_0_011100010100;
      patterns[7251] = 29'b0_001110001010_011_0_111000101000;
      patterns[7252] = 29'b0_001110001010_100_0_000111000101;
      patterns[7253] = 29'b0_001110001010_101_1_000011100010;
      patterns[7254] = 29'b0_001110001010_110_0_001110001010;
      patterns[7255] = 29'b0_001110001010_111_0_001110001010;
      patterns[7256] = 29'b0_001110001011_000_0_001110001011;
      patterns[7257] = 29'b0_001110001011_001_0_001011001110;
      patterns[7258] = 29'b0_001110001011_010_0_011100010110;
      patterns[7259] = 29'b0_001110001011_011_0_111000101100;
      patterns[7260] = 29'b0_001110001011_100_1_000111000101;
      patterns[7261] = 29'b0_001110001011_101_1_100011100010;
      patterns[7262] = 29'b0_001110001011_110_0_001110001011;
      patterns[7263] = 29'b0_001110001011_111_0_001110001011;
      patterns[7264] = 29'b0_001110001100_000_0_001110001100;
      patterns[7265] = 29'b0_001110001100_001_0_001100001110;
      patterns[7266] = 29'b0_001110001100_010_0_011100011000;
      patterns[7267] = 29'b0_001110001100_011_0_111000110000;
      patterns[7268] = 29'b0_001110001100_100_0_000111000110;
      patterns[7269] = 29'b0_001110001100_101_0_000011100011;
      patterns[7270] = 29'b0_001110001100_110_0_001110001100;
      patterns[7271] = 29'b0_001110001100_111_0_001110001100;
      patterns[7272] = 29'b0_001110001101_000_0_001110001101;
      patterns[7273] = 29'b0_001110001101_001_0_001101001110;
      patterns[7274] = 29'b0_001110001101_010_0_011100011010;
      patterns[7275] = 29'b0_001110001101_011_0_111000110100;
      patterns[7276] = 29'b0_001110001101_100_1_000111000110;
      patterns[7277] = 29'b0_001110001101_101_0_100011100011;
      patterns[7278] = 29'b0_001110001101_110_0_001110001101;
      patterns[7279] = 29'b0_001110001101_111_0_001110001101;
      patterns[7280] = 29'b0_001110001110_000_0_001110001110;
      patterns[7281] = 29'b0_001110001110_001_0_001110001110;
      patterns[7282] = 29'b0_001110001110_010_0_011100011100;
      patterns[7283] = 29'b0_001110001110_011_0_111000111000;
      patterns[7284] = 29'b0_001110001110_100_0_000111000111;
      patterns[7285] = 29'b0_001110001110_101_1_000011100011;
      patterns[7286] = 29'b0_001110001110_110_0_001110001110;
      patterns[7287] = 29'b0_001110001110_111_0_001110001110;
      patterns[7288] = 29'b0_001110001111_000_0_001110001111;
      patterns[7289] = 29'b0_001110001111_001_0_001111001110;
      patterns[7290] = 29'b0_001110001111_010_0_011100011110;
      patterns[7291] = 29'b0_001110001111_011_0_111000111100;
      patterns[7292] = 29'b0_001110001111_100_1_000111000111;
      patterns[7293] = 29'b0_001110001111_101_1_100011100011;
      patterns[7294] = 29'b0_001110001111_110_0_001110001111;
      patterns[7295] = 29'b0_001110001111_111_0_001110001111;
      patterns[7296] = 29'b0_001110010000_000_0_001110010000;
      patterns[7297] = 29'b0_001110010000_001_0_010000001110;
      patterns[7298] = 29'b0_001110010000_010_0_011100100000;
      patterns[7299] = 29'b0_001110010000_011_0_111001000000;
      patterns[7300] = 29'b0_001110010000_100_0_000111001000;
      patterns[7301] = 29'b0_001110010000_101_0_000011100100;
      patterns[7302] = 29'b0_001110010000_110_0_001110010000;
      patterns[7303] = 29'b0_001110010000_111_0_001110010000;
      patterns[7304] = 29'b0_001110010001_000_0_001110010001;
      patterns[7305] = 29'b0_001110010001_001_0_010001001110;
      patterns[7306] = 29'b0_001110010001_010_0_011100100010;
      patterns[7307] = 29'b0_001110010001_011_0_111001000100;
      patterns[7308] = 29'b0_001110010001_100_1_000111001000;
      patterns[7309] = 29'b0_001110010001_101_0_100011100100;
      patterns[7310] = 29'b0_001110010001_110_0_001110010001;
      patterns[7311] = 29'b0_001110010001_111_0_001110010001;
      patterns[7312] = 29'b0_001110010010_000_0_001110010010;
      patterns[7313] = 29'b0_001110010010_001_0_010010001110;
      patterns[7314] = 29'b0_001110010010_010_0_011100100100;
      patterns[7315] = 29'b0_001110010010_011_0_111001001000;
      patterns[7316] = 29'b0_001110010010_100_0_000111001001;
      patterns[7317] = 29'b0_001110010010_101_1_000011100100;
      patterns[7318] = 29'b0_001110010010_110_0_001110010010;
      patterns[7319] = 29'b0_001110010010_111_0_001110010010;
      patterns[7320] = 29'b0_001110010011_000_0_001110010011;
      patterns[7321] = 29'b0_001110010011_001_0_010011001110;
      patterns[7322] = 29'b0_001110010011_010_0_011100100110;
      patterns[7323] = 29'b0_001110010011_011_0_111001001100;
      patterns[7324] = 29'b0_001110010011_100_1_000111001001;
      patterns[7325] = 29'b0_001110010011_101_1_100011100100;
      patterns[7326] = 29'b0_001110010011_110_0_001110010011;
      patterns[7327] = 29'b0_001110010011_111_0_001110010011;
      patterns[7328] = 29'b0_001110010100_000_0_001110010100;
      patterns[7329] = 29'b0_001110010100_001_0_010100001110;
      patterns[7330] = 29'b0_001110010100_010_0_011100101000;
      patterns[7331] = 29'b0_001110010100_011_0_111001010000;
      patterns[7332] = 29'b0_001110010100_100_0_000111001010;
      patterns[7333] = 29'b0_001110010100_101_0_000011100101;
      patterns[7334] = 29'b0_001110010100_110_0_001110010100;
      patterns[7335] = 29'b0_001110010100_111_0_001110010100;
      patterns[7336] = 29'b0_001110010101_000_0_001110010101;
      patterns[7337] = 29'b0_001110010101_001_0_010101001110;
      patterns[7338] = 29'b0_001110010101_010_0_011100101010;
      patterns[7339] = 29'b0_001110010101_011_0_111001010100;
      patterns[7340] = 29'b0_001110010101_100_1_000111001010;
      patterns[7341] = 29'b0_001110010101_101_0_100011100101;
      patterns[7342] = 29'b0_001110010101_110_0_001110010101;
      patterns[7343] = 29'b0_001110010101_111_0_001110010101;
      patterns[7344] = 29'b0_001110010110_000_0_001110010110;
      patterns[7345] = 29'b0_001110010110_001_0_010110001110;
      patterns[7346] = 29'b0_001110010110_010_0_011100101100;
      patterns[7347] = 29'b0_001110010110_011_0_111001011000;
      patterns[7348] = 29'b0_001110010110_100_0_000111001011;
      patterns[7349] = 29'b0_001110010110_101_1_000011100101;
      patterns[7350] = 29'b0_001110010110_110_0_001110010110;
      patterns[7351] = 29'b0_001110010110_111_0_001110010110;
      patterns[7352] = 29'b0_001110010111_000_0_001110010111;
      patterns[7353] = 29'b0_001110010111_001_0_010111001110;
      patterns[7354] = 29'b0_001110010111_010_0_011100101110;
      patterns[7355] = 29'b0_001110010111_011_0_111001011100;
      patterns[7356] = 29'b0_001110010111_100_1_000111001011;
      patterns[7357] = 29'b0_001110010111_101_1_100011100101;
      patterns[7358] = 29'b0_001110010111_110_0_001110010111;
      patterns[7359] = 29'b0_001110010111_111_0_001110010111;
      patterns[7360] = 29'b0_001110011000_000_0_001110011000;
      patterns[7361] = 29'b0_001110011000_001_0_011000001110;
      patterns[7362] = 29'b0_001110011000_010_0_011100110000;
      patterns[7363] = 29'b0_001110011000_011_0_111001100000;
      patterns[7364] = 29'b0_001110011000_100_0_000111001100;
      patterns[7365] = 29'b0_001110011000_101_0_000011100110;
      patterns[7366] = 29'b0_001110011000_110_0_001110011000;
      patterns[7367] = 29'b0_001110011000_111_0_001110011000;
      patterns[7368] = 29'b0_001110011001_000_0_001110011001;
      patterns[7369] = 29'b0_001110011001_001_0_011001001110;
      patterns[7370] = 29'b0_001110011001_010_0_011100110010;
      patterns[7371] = 29'b0_001110011001_011_0_111001100100;
      patterns[7372] = 29'b0_001110011001_100_1_000111001100;
      patterns[7373] = 29'b0_001110011001_101_0_100011100110;
      patterns[7374] = 29'b0_001110011001_110_0_001110011001;
      patterns[7375] = 29'b0_001110011001_111_0_001110011001;
      patterns[7376] = 29'b0_001110011010_000_0_001110011010;
      patterns[7377] = 29'b0_001110011010_001_0_011010001110;
      patterns[7378] = 29'b0_001110011010_010_0_011100110100;
      patterns[7379] = 29'b0_001110011010_011_0_111001101000;
      patterns[7380] = 29'b0_001110011010_100_0_000111001101;
      patterns[7381] = 29'b0_001110011010_101_1_000011100110;
      patterns[7382] = 29'b0_001110011010_110_0_001110011010;
      patterns[7383] = 29'b0_001110011010_111_0_001110011010;
      patterns[7384] = 29'b0_001110011011_000_0_001110011011;
      patterns[7385] = 29'b0_001110011011_001_0_011011001110;
      patterns[7386] = 29'b0_001110011011_010_0_011100110110;
      patterns[7387] = 29'b0_001110011011_011_0_111001101100;
      patterns[7388] = 29'b0_001110011011_100_1_000111001101;
      patterns[7389] = 29'b0_001110011011_101_1_100011100110;
      patterns[7390] = 29'b0_001110011011_110_0_001110011011;
      patterns[7391] = 29'b0_001110011011_111_0_001110011011;
      patterns[7392] = 29'b0_001110011100_000_0_001110011100;
      patterns[7393] = 29'b0_001110011100_001_0_011100001110;
      patterns[7394] = 29'b0_001110011100_010_0_011100111000;
      patterns[7395] = 29'b0_001110011100_011_0_111001110000;
      patterns[7396] = 29'b0_001110011100_100_0_000111001110;
      patterns[7397] = 29'b0_001110011100_101_0_000011100111;
      patterns[7398] = 29'b0_001110011100_110_0_001110011100;
      patterns[7399] = 29'b0_001110011100_111_0_001110011100;
      patterns[7400] = 29'b0_001110011101_000_0_001110011101;
      patterns[7401] = 29'b0_001110011101_001_0_011101001110;
      patterns[7402] = 29'b0_001110011101_010_0_011100111010;
      patterns[7403] = 29'b0_001110011101_011_0_111001110100;
      patterns[7404] = 29'b0_001110011101_100_1_000111001110;
      patterns[7405] = 29'b0_001110011101_101_0_100011100111;
      patterns[7406] = 29'b0_001110011101_110_0_001110011101;
      patterns[7407] = 29'b0_001110011101_111_0_001110011101;
      patterns[7408] = 29'b0_001110011110_000_0_001110011110;
      patterns[7409] = 29'b0_001110011110_001_0_011110001110;
      patterns[7410] = 29'b0_001110011110_010_0_011100111100;
      patterns[7411] = 29'b0_001110011110_011_0_111001111000;
      patterns[7412] = 29'b0_001110011110_100_0_000111001111;
      patterns[7413] = 29'b0_001110011110_101_1_000011100111;
      patterns[7414] = 29'b0_001110011110_110_0_001110011110;
      patterns[7415] = 29'b0_001110011110_111_0_001110011110;
      patterns[7416] = 29'b0_001110011111_000_0_001110011111;
      patterns[7417] = 29'b0_001110011111_001_0_011111001110;
      patterns[7418] = 29'b0_001110011111_010_0_011100111110;
      patterns[7419] = 29'b0_001110011111_011_0_111001111100;
      patterns[7420] = 29'b0_001110011111_100_1_000111001111;
      patterns[7421] = 29'b0_001110011111_101_1_100011100111;
      patterns[7422] = 29'b0_001110011111_110_0_001110011111;
      patterns[7423] = 29'b0_001110011111_111_0_001110011111;
      patterns[7424] = 29'b0_001110100000_000_0_001110100000;
      patterns[7425] = 29'b0_001110100000_001_0_100000001110;
      patterns[7426] = 29'b0_001110100000_010_0_011101000000;
      patterns[7427] = 29'b0_001110100000_011_0_111010000000;
      patterns[7428] = 29'b0_001110100000_100_0_000111010000;
      patterns[7429] = 29'b0_001110100000_101_0_000011101000;
      patterns[7430] = 29'b0_001110100000_110_0_001110100000;
      patterns[7431] = 29'b0_001110100000_111_0_001110100000;
      patterns[7432] = 29'b0_001110100001_000_0_001110100001;
      patterns[7433] = 29'b0_001110100001_001_0_100001001110;
      patterns[7434] = 29'b0_001110100001_010_0_011101000010;
      patterns[7435] = 29'b0_001110100001_011_0_111010000100;
      patterns[7436] = 29'b0_001110100001_100_1_000111010000;
      patterns[7437] = 29'b0_001110100001_101_0_100011101000;
      patterns[7438] = 29'b0_001110100001_110_0_001110100001;
      patterns[7439] = 29'b0_001110100001_111_0_001110100001;
      patterns[7440] = 29'b0_001110100010_000_0_001110100010;
      patterns[7441] = 29'b0_001110100010_001_0_100010001110;
      patterns[7442] = 29'b0_001110100010_010_0_011101000100;
      patterns[7443] = 29'b0_001110100010_011_0_111010001000;
      patterns[7444] = 29'b0_001110100010_100_0_000111010001;
      patterns[7445] = 29'b0_001110100010_101_1_000011101000;
      patterns[7446] = 29'b0_001110100010_110_0_001110100010;
      patterns[7447] = 29'b0_001110100010_111_0_001110100010;
      patterns[7448] = 29'b0_001110100011_000_0_001110100011;
      patterns[7449] = 29'b0_001110100011_001_0_100011001110;
      patterns[7450] = 29'b0_001110100011_010_0_011101000110;
      patterns[7451] = 29'b0_001110100011_011_0_111010001100;
      patterns[7452] = 29'b0_001110100011_100_1_000111010001;
      patterns[7453] = 29'b0_001110100011_101_1_100011101000;
      patterns[7454] = 29'b0_001110100011_110_0_001110100011;
      patterns[7455] = 29'b0_001110100011_111_0_001110100011;
      patterns[7456] = 29'b0_001110100100_000_0_001110100100;
      patterns[7457] = 29'b0_001110100100_001_0_100100001110;
      patterns[7458] = 29'b0_001110100100_010_0_011101001000;
      patterns[7459] = 29'b0_001110100100_011_0_111010010000;
      patterns[7460] = 29'b0_001110100100_100_0_000111010010;
      patterns[7461] = 29'b0_001110100100_101_0_000011101001;
      patterns[7462] = 29'b0_001110100100_110_0_001110100100;
      patterns[7463] = 29'b0_001110100100_111_0_001110100100;
      patterns[7464] = 29'b0_001110100101_000_0_001110100101;
      patterns[7465] = 29'b0_001110100101_001_0_100101001110;
      patterns[7466] = 29'b0_001110100101_010_0_011101001010;
      patterns[7467] = 29'b0_001110100101_011_0_111010010100;
      patterns[7468] = 29'b0_001110100101_100_1_000111010010;
      patterns[7469] = 29'b0_001110100101_101_0_100011101001;
      patterns[7470] = 29'b0_001110100101_110_0_001110100101;
      patterns[7471] = 29'b0_001110100101_111_0_001110100101;
      patterns[7472] = 29'b0_001110100110_000_0_001110100110;
      patterns[7473] = 29'b0_001110100110_001_0_100110001110;
      patterns[7474] = 29'b0_001110100110_010_0_011101001100;
      patterns[7475] = 29'b0_001110100110_011_0_111010011000;
      patterns[7476] = 29'b0_001110100110_100_0_000111010011;
      patterns[7477] = 29'b0_001110100110_101_1_000011101001;
      patterns[7478] = 29'b0_001110100110_110_0_001110100110;
      patterns[7479] = 29'b0_001110100110_111_0_001110100110;
      patterns[7480] = 29'b0_001110100111_000_0_001110100111;
      patterns[7481] = 29'b0_001110100111_001_0_100111001110;
      patterns[7482] = 29'b0_001110100111_010_0_011101001110;
      patterns[7483] = 29'b0_001110100111_011_0_111010011100;
      patterns[7484] = 29'b0_001110100111_100_1_000111010011;
      patterns[7485] = 29'b0_001110100111_101_1_100011101001;
      patterns[7486] = 29'b0_001110100111_110_0_001110100111;
      patterns[7487] = 29'b0_001110100111_111_0_001110100111;
      patterns[7488] = 29'b0_001110101000_000_0_001110101000;
      patterns[7489] = 29'b0_001110101000_001_0_101000001110;
      patterns[7490] = 29'b0_001110101000_010_0_011101010000;
      patterns[7491] = 29'b0_001110101000_011_0_111010100000;
      patterns[7492] = 29'b0_001110101000_100_0_000111010100;
      patterns[7493] = 29'b0_001110101000_101_0_000011101010;
      patterns[7494] = 29'b0_001110101000_110_0_001110101000;
      patterns[7495] = 29'b0_001110101000_111_0_001110101000;
      patterns[7496] = 29'b0_001110101001_000_0_001110101001;
      patterns[7497] = 29'b0_001110101001_001_0_101001001110;
      patterns[7498] = 29'b0_001110101001_010_0_011101010010;
      patterns[7499] = 29'b0_001110101001_011_0_111010100100;
      patterns[7500] = 29'b0_001110101001_100_1_000111010100;
      patterns[7501] = 29'b0_001110101001_101_0_100011101010;
      patterns[7502] = 29'b0_001110101001_110_0_001110101001;
      patterns[7503] = 29'b0_001110101001_111_0_001110101001;
      patterns[7504] = 29'b0_001110101010_000_0_001110101010;
      patterns[7505] = 29'b0_001110101010_001_0_101010001110;
      patterns[7506] = 29'b0_001110101010_010_0_011101010100;
      patterns[7507] = 29'b0_001110101010_011_0_111010101000;
      patterns[7508] = 29'b0_001110101010_100_0_000111010101;
      patterns[7509] = 29'b0_001110101010_101_1_000011101010;
      patterns[7510] = 29'b0_001110101010_110_0_001110101010;
      patterns[7511] = 29'b0_001110101010_111_0_001110101010;
      patterns[7512] = 29'b0_001110101011_000_0_001110101011;
      patterns[7513] = 29'b0_001110101011_001_0_101011001110;
      patterns[7514] = 29'b0_001110101011_010_0_011101010110;
      patterns[7515] = 29'b0_001110101011_011_0_111010101100;
      patterns[7516] = 29'b0_001110101011_100_1_000111010101;
      patterns[7517] = 29'b0_001110101011_101_1_100011101010;
      patterns[7518] = 29'b0_001110101011_110_0_001110101011;
      patterns[7519] = 29'b0_001110101011_111_0_001110101011;
      patterns[7520] = 29'b0_001110101100_000_0_001110101100;
      patterns[7521] = 29'b0_001110101100_001_0_101100001110;
      patterns[7522] = 29'b0_001110101100_010_0_011101011000;
      patterns[7523] = 29'b0_001110101100_011_0_111010110000;
      patterns[7524] = 29'b0_001110101100_100_0_000111010110;
      patterns[7525] = 29'b0_001110101100_101_0_000011101011;
      patterns[7526] = 29'b0_001110101100_110_0_001110101100;
      patterns[7527] = 29'b0_001110101100_111_0_001110101100;
      patterns[7528] = 29'b0_001110101101_000_0_001110101101;
      patterns[7529] = 29'b0_001110101101_001_0_101101001110;
      patterns[7530] = 29'b0_001110101101_010_0_011101011010;
      patterns[7531] = 29'b0_001110101101_011_0_111010110100;
      patterns[7532] = 29'b0_001110101101_100_1_000111010110;
      patterns[7533] = 29'b0_001110101101_101_0_100011101011;
      patterns[7534] = 29'b0_001110101101_110_0_001110101101;
      patterns[7535] = 29'b0_001110101101_111_0_001110101101;
      patterns[7536] = 29'b0_001110101110_000_0_001110101110;
      patterns[7537] = 29'b0_001110101110_001_0_101110001110;
      patterns[7538] = 29'b0_001110101110_010_0_011101011100;
      patterns[7539] = 29'b0_001110101110_011_0_111010111000;
      patterns[7540] = 29'b0_001110101110_100_0_000111010111;
      patterns[7541] = 29'b0_001110101110_101_1_000011101011;
      patterns[7542] = 29'b0_001110101110_110_0_001110101110;
      patterns[7543] = 29'b0_001110101110_111_0_001110101110;
      patterns[7544] = 29'b0_001110101111_000_0_001110101111;
      patterns[7545] = 29'b0_001110101111_001_0_101111001110;
      patterns[7546] = 29'b0_001110101111_010_0_011101011110;
      patterns[7547] = 29'b0_001110101111_011_0_111010111100;
      patterns[7548] = 29'b0_001110101111_100_1_000111010111;
      patterns[7549] = 29'b0_001110101111_101_1_100011101011;
      patterns[7550] = 29'b0_001110101111_110_0_001110101111;
      patterns[7551] = 29'b0_001110101111_111_0_001110101111;
      patterns[7552] = 29'b0_001110110000_000_0_001110110000;
      patterns[7553] = 29'b0_001110110000_001_0_110000001110;
      patterns[7554] = 29'b0_001110110000_010_0_011101100000;
      patterns[7555] = 29'b0_001110110000_011_0_111011000000;
      patterns[7556] = 29'b0_001110110000_100_0_000111011000;
      patterns[7557] = 29'b0_001110110000_101_0_000011101100;
      patterns[7558] = 29'b0_001110110000_110_0_001110110000;
      patterns[7559] = 29'b0_001110110000_111_0_001110110000;
      patterns[7560] = 29'b0_001110110001_000_0_001110110001;
      patterns[7561] = 29'b0_001110110001_001_0_110001001110;
      patterns[7562] = 29'b0_001110110001_010_0_011101100010;
      patterns[7563] = 29'b0_001110110001_011_0_111011000100;
      patterns[7564] = 29'b0_001110110001_100_1_000111011000;
      patterns[7565] = 29'b0_001110110001_101_0_100011101100;
      patterns[7566] = 29'b0_001110110001_110_0_001110110001;
      patterns[7567] = 29'b0_001110110001_111_0_001110110001;
      patterns[7568] = 29'b0_001110110010_000_0_001110110010;
      patterns[7569] = 29'b0_001110110010_001_0_110010001110;
      patterns[7570] = 29'b0_001110110010_010_0_011101100100;
      patterns[7571] = 29'b0_001110110010_011_0_111011001000;
      patterns[7572] = 29'b0_001110110010_100_0_000111011001;
      patterns[7573] = 29'b0_001110110010_101_1_000011101100;
      patterns[7574] = 29'b0_001110110010_110_0_001110110010;
      patterns[7575] = 29'b0_001110110010_111_0_001110110010;
      patterns[7576] = 29'b0_001110110011_000_0_001110110011;
      patterns[7577] = 29'b0_001110110011_001_0_110011001110;
      patterns[7578] = 29'b0_001110110011_010_0_011101100110;
      patterns[7579] = 29'b0_001110110011_011_0_111011001100;
      patterns[7580] = 29'b0_001110110011_100_1_000111011001;
      patterns[7581] = 29'b0_001110110011_101_1_100011101100;
      patterns[7582] = 29'b0_001110110011_110_0_001110110011;
      patterns[7583] = 29'b0_001110110011_111_0_001110110011;
      patterns[7584] = 29'b0_001110110100_000_0_001110110100;
      patterns[7585] = 29'b0_001110110100_001_0_110100001110;
      patterns[7586] = 29'b0_001110110100_010_0_011101101000;
      patterns[7587] = 29'b0_001110110100_011_0_111011010000;
      patterns[7588] = 29'b0_001110110100_100_0_000111011010;
      patterns[7589] = 29'b0_001110110100_101_0_000011101101;
      patterns[7590] = 29'b0_001110110100_110_0_001110110100;
      patterns[7591] = 29'b0_001110110100_111_0_001110110100;
      patterns[7592] = 29'b0_001110110101_000_0_001110110101;
      patterns[7593] = 29'b0_001110110101_001_0_110101001110;
      patterns[7594] = 29'b0_001110110101_010_0_011101101010;
      patterns[7595] = 29'b0_001110110101_011_0_111011010100;
      patterns[7596] = 29'b0_001110110101_100_1_000111011010;
      patterns[7597] = 29'b0_001110110101_101_0_100011101101;
      patterns[7598] = 29'b0_001110110101_110_0_001110110101;
      patterns[7599] = 29'b0_001110110101_111_0_001110110101;
      patterns[7600] = 29'b0_001110110110_000_0_001110110110;
      patterns[7601] = 29'b0_001110110110_001_0_110110001110;
      patterns[7602] = 29'b0_001110110110_010_0_011101101100;
      patterns[7603] = 29'b0_001110110110_011_0_111011011000;
      patterns[7604] = 29'b0_001110110110_100_0_000111011011;
      patterns[7605] = 29'b0_001110110110_101_1_000011101101;
      patterns[7606] = 29'b0_001110110110_110_0_001110110110;
      patterns[7607] = 29'b0_001110110110_111_0_001110110110;
      patterns[7608] = 29'b0_001110110111_000_0_001110110111;
      patterns[7609] = 29'b0_001110110111_001_0_110111001110;
      patterns[7610] = 29'b0_001110110111_010_0_011101101110;
      patterns[7611] = 29'b0_001110110111_011_0_111011011100;
      patterns[7612] = 29'b0_001110110111_100_1_000111011011;
      patterns[7613] = 29'b0_001110110111_101_1_100011101101;
      patterns[7614] = 29'b0_001110110111_110_0_001110110111;
      patterns[7615] = 29'b0_001110110111_111_0_001110110111;
      patterns[7616] = 29'b0_001110111000_000_0_001110111000;
      patterns[7617] = 29'b0_001110111000_001_0_111000001110;
      patterns[7618] = 29'b0_001110111000_010_0_011101110000;
      patterns[7619] = 29'b0_001110111000_011_0_111011100000;
      patterns[7620] = 29'b0_001110111000_100_0_000111011100;
      patterns[7621] = 29'b0_001110111000_101_0_000011101110;
      patterns[7622] = 29'b0_001110111000_110_0_001110111000;
      patterns[7623] = 29'b0_001110111000_111_0_001110111000;
      patterns[7624] = 29'b0_001110111001_000_0_001110111001;
      patterns[7625] = 29'b0_001110111001_001_0_111001001110;
      patterns[7626] = 29'b0_001110111001_010_0_011101110010;
      patterns[7627] = 29'b0_001110111001_011_0_111011100100;
      patterns[7628] = 29'b0_001110111001_100_1_000111011100;
      patterns[7629] = 29'b0_001110111001_101_0_100011101110;
      patterns[7630] = 29'b0_001110111001_110_0_001110111001;
      patterns[7631] = 29'b0_001110111001_111_0_001110111001;
      patterns[7632] = 29'b0_001110111010_000_0_001110111010;
      patterns[7633] = 29'b0_001110111010_001_0_111010001110;
      patterns[7634] = 29'b0_001110111010_010_0_011101110100;
      patterns[7635] = 29'b0_001110111010_011_0_111011101000;
      patterns[7636] = 29'b0_001110111010_100_0_000111011101;
      patterns[7637] = 29'b0_001110111010_101_1_000011101110;
      patterns[7638] = 29'b0_001110111010_110_0_001110111010;
      patterns[7639] = 29'b0_001110111010_111_0_001110111010;
      patterns[7640] = 29'b0_001110111011_000_0_001110111011;
      patterns[7641] = 29'b0_001110111011_001_0_111011001110;
      patterns[7642] = 29'b0_001110111011_010_0_011101110110;
      patterns[7643] = 29'b0_001110111011_011_0_111011101100;
      patterns[7644] = 29'b0_001110111011_100_1_000111011101;
      patterns[7645] = 29'b0_001110111011_101_1_100011101110;
      patterns[7646] = 29'b0_001110111011_110_0_001110111011;
      patterns[7647] = 29'b0_001110111011_111_0_001110111011;
      patterns[7648] = 29'b0_001110111100_000_0_001110111100;
      patterns[7649] = 29'b0_001110111100_001_0_111100001110;
      patterns[7650] = 29'b0_001110111100_010_0_011101111000;
      patterns[7651] = 29'b0_001110111100_011_0_111011110000;
      patterns[7652] = 29'b0_001110111100_100_0_000111011110;
      patterns[7653] = 29'b0_001110111100_101_0_000011101111;
      patterns[7654] = 29'b0_001110111100_110_0_001110111100;
      patterns[7655] = 29'b0_001110111100_111_0_001110111100;
      patterns[7656] = 29'b0_001110111101_000_0_001110111101;
      patterns[7657] = 29'b0_001110111101_001_0_111101001110;
      patterns[7658] = 29'b0_001110111101_010_0_011101111010;
      patterns[7659] = 29'b0_001110111101_011_0_111011110100;
      patterns[7660] = 29'b0_001110111101_100_1_000111011110;
      patterns[7661] = 29'b0_001110111101_101_0_100011101111;
      patterns[7662] = 29'b0_001110111101_110_0_001110111101;
      patterns[7663] = 29'b0_001110111101_111_0_001110111101;
      patterns[7664] = 29'b0_001110111110_000_0_001110111110;
      patterns[7665] = 29'b0_001110111110_001_0_111110001110;
      patterns[7666] = 29'b0_001110111110_010_0_011101111100;
      patterns[7667] = 29'b0_001110111110_011_0_111011111000;
      patterns[7668] = 29'b0_001110111110_100_0_000111011111;
      patterns[7669] = 29'b0_001110111110_101_1_000011101111;
      patterns[7670] = 29'b0_001110111110_110_0_001110111110;
      patterns[7671] = 29'b0_001110111110_111_0_001110111110;
      patterns[7672] = 29'b0_001110111111_000_0_001110111111;
      patterns[7673] = 29'b0_001110111111_001_0_111111001110;
      patterns[7674] = 29'b0_001110111111_010_0_011101111110;
      patterns[7675] = 29'b0_001110111111_011_0_111011111100;
      patterns[7676] = 29'b0_001110111111_100_1_000111011111;
      patterns[7677] = 29'b0_001110111111_101_1_100011101111;
      patterns[7678] = 29'b0_001110111111_110_0_001110111111;
      patterns[7679] = 29'b0_001110111111_111_0_001110111111;
      patterns[7680] = 29'b0_001111000000_000_0_001111000000;
      patterns[7681] = 29'b0_001111000000_001_0_000000001111;
      patterns[7682] = 29'b0_001111000000_010_0_011110000000;
      patterns[7683] = 29'b0_001111000000_011_0_111100000000;
      patterns[7684] = 29'b0_001111000000_100_0_000111100000;
      patterns[7685] = 29'b0_001111000000_101_0_000011110000;
      patterns[7686] = 29'b0_001111000000_110_0_001111000000;
      patterns[7687] = 29'b0_001111000000_111_0_001111000000;
      patterns[7688] = 29'b0_001111000001_000_0_001111000001;
      patterns[7689] = 29'b0_001111000001_001_0_000001001111;
      patterns[7690] = 29'b0_001111000001_010_0_011110000010;
      patterns[7691] = 29'b0_001111000001_011_0_111100000100;
      patterns[7692] = 29'b0_001111000001_100_1_000111100000;
      patterns[7693] = 29'b0_001111000001_101_0_100011110000;
      patterns[7694] = 29'b0_001111000001_110_0_001111000001;
      patterns[7695] = 29'b0_001111000001_111_0_001111000001;
      patterns[7696] = 29'b0_001111000010_000_0_001111000010;
      patterns[7697] = 29'b0_001111000010_001_0_000010001111;
      patterns[7698] = 29'b0_001111000010_010_0_011110000100;
      patterns[7699] = 29'b0_001111000010_011_0_111100001000;
      patterns[7700] = 29'b0_001111000010_100_0_000111100001;
      patterns[7701] = 29'b0_001111000010_101_1_000011110000;
      patterns[7702] = 29'b0_001111000010_110_0_001111000010;
      patterns[7703] = 29'b0_001111000010_111_0_001111000010;
      patterns[7704] = 29'b0_001111000011_000_0_001111000011;
      patterns[7705] = 29'b0_001111000011_001_0_000011001111;
      patterns[7706] = 29'b0_001111000011_010_0_011110000110;
      patterns[7707] = 29'b0_001111000011_011_0_111100001100;
      patterns[7708] = 29'b0_001111000011_100_1_000111100001;
      patterns[7709] = 29'b0_001111000011_101_1_100011110000;
      patterns[7710] = 29'b0_001111000011_110_0_001111000011;
      patterns[7711] = 29'b0_001111000011_111_0_001111000011;
      patterns[7712] = 29'b0_001111000100_000_0_001111000100;
      patterns[7713] = 29'b0_001111000100_001_0_000100001111;
      patterns[7714] = 29'b0_001111000100_010_0_011110001000;
      patterns[7715] = 29'b0_001111000100_011_0_111100010000;
      patterns[7716] = 29'b0_001111000100_100_0_000111100010;
      patterns[7717] = 29'b0_001111000100_101_0_000011110001;
      patterns[7718] = 29'b0_001111000100_110_0_001111000100;
      patterns[7719] = 29'b0_001111000100_111_0_001111000100;
      patterns[7720] = 29'b0_001111000101_000_0_001111000101;
      patterns[7721] = 29'b0_001111000101_001_0_000101001111;
      patterns[7722] = 29'b0_001111000101_010_0_011110001010;
      patterns[7723] = 29'b0_001111000101_011_0_111100010100;
      patterns[7724] = 29'b0_001111000101_100_1_000111100010;
      patterns[7725] = 29'b0_001111000101_101_0_100011110001;
      patterns[7726] = 29'b0_001111000101_110_0_001111000101;
      patterns[7727] = 29'b0_001111000101_111_0_001111000101;
      patterns[7728] = 29'b0_001111000110_000_0_001111000110;
      patterns[7729] = 29'b0_001111000110_001_0_000110001111;
      patterns[7730] = 29'b0_001111000110_010_0_011110001100;
      patterns[7731] = 29'b0_001111000110_011_0_111100011000;
      patterns[7732] = 29'b0_001111000110_100_0_000111100011;
      patterns[7733] = 29'b0_001111000110_101_1_000011110001;
      patterns[7734] = 29'b0_001111000110_110_0_001111000110;
      patterns[7735] = 29'b0_001111000110_111_0_001111000110;
      patterns[7736] = 29'b0_001111000111_000_0_001111000111;
      patterns[7737] = 29'b0_001111000111_001_0_000111001111;
      patterns[7738] = 29'b0_001111000111_010_0_011110001110;
      patterns[7739] = 29'b0_001111000111_011_0_111100011100;
      patterns[7740] = 29'b0_001111000111_100_1_000111100011;
      patterns[7741] = 29'b0_001111000111_101_1_100011110001;
      patterns[7742] = 29'b0_001111000111_110_0_001111000111;
      patterns[7743] = 29'b0_001111000111_111_0_001111000111;
      patterns[7744] = 29'b0_001111001000_000_0_001111001000;
      patterns[7745] = 29'b0_001111001000_001_0_001000001111;
      patterns[7746] = 29'b0_001111001000_010_0_011110010000;
      patterns[7747] = 29'b0_001111001000_011_0_111100100000;
      patterns[7748] = 29'b0_001111001000_100_0_000111100100;
      patterns[7749] = 29'b0_001111001000_101_0_000011110010;
      patterns[7750] = 29'b0_001111001000_110_0_001111001000;
      patterns[7751] = 29'b0_001111001000_111_0_001111001000;
      patterns[7752] = 29'b0_001111001001_000_0_001111001001;
      patterns[7753] = 29'b0_001111001001_001_0_001001001111;
      patterns[7754] = 29'b0_001111001001_010_0_011110010010;
      patterns[7755] = 29'b0_001111001001_011_0_111100100100;
      patterns[7756] = 29'b0_001111001001_100_1_000111100100;
      patterns[7757] = 29'b0_001111001001_101_0_100011110010;
      patterns[7758] = 29'b0_001111001001_110_0_001111001001;
      patterns[7759] = 29'b0_001111001001_111_0_001111001001;
      patterns[7760] = 29'b0_001111001010_000_0_001111001010;
      patterns[7761] = 29'b0_001111001010_001_0_001010001111;
      patterns[7762] = 29'b0_001111001010_010_0_011110010100;
      patterns[7763] = 29'b0_001111001010_011_0_111100101000;
      patterns[7764] = 29'b0_001111001010_100_0_000111100101;
      patterns[7765] = 29'b0_001111001010_101_1_000011110010;
      patterns[7766] = 29'b0_001111001010_110_0_001111001010;
      patterns[7767] = 29'b0_001111001010_111_0_001111001010;
      patterns[7768] = 29'b0_001111001011_000_0_001111001011;
      patterns[7769] = 29'b0_001111001011_001_0_001011001111;
      patterns[7770] = 29'b0_001111001011_010_0_011110010110;
      patterns[7771] = 29'b0_001111001011_011_0_111100101100;
      patterns[7772] = 29'b0_001111001011_100_1_000111100101;
      patterns[7773] = 29'b0_001111001011_101_1_100011110010;
      patterns[7774] = 29'b0_001111001011_110_0_001111001011;
      patterns[7775] = 29'b0_001111001011_111_0_001111001011;
      patterns[7776] = 29'b0_001111001100_000_0_001111001100;
      patterns[7777] = 29'b0_001111001100_001_0_001100001111;
      patterns[7778] = 29'b0_001111001100_010_0_011110011000;
      patterns[7779] = 29'b0_001111001100_011_0_111100110000;
      patterns[7780] = 29'b0_001111001100_100_0_000111100110;
      patterns[7781] = 29'b0_001111001100_101_0_000011110011;
      patterns[7782] = 29'b0_001111001100_110_0_001111001100;
      patterns[7783] = 29'b0_001111001100_111_0_001111001100;
      patterns[7784] = 29'b0_001111001101_000_0_001111001101;
      patterns[7785] = 29'b0_001111001101_001_0_001101001111;
      patterns[7786] = 29'b0_001111001101_010_0_011110011010;
      patterns[7787] = 29'b0_001111001101_011_0_111100110100;
      patterns[7788] = 29'b0_001111001101_100_1_000111100110;
      patterns[7789] = 29'b0_001111001101_101_0_100011110011;
      patterns[7790] = 29'b0_001111001101_110_0_001111001101;
      patterns[7791] = 29'b0_001111001101_111_0_001111001101;
      patterns[7792] = 29'b0_001111001110_000_0_001111001110;
      patterns[7793] = 29'b0_001111001110_001_0_001110001111;
      patterns[7794] = 29'b0_001111001110_010_0_011110011100;
      patterns[7795] = 29'b0_001111001110_011_0_111100111000;
      patterns[7796] = 29'b0_001111001110_100_0_000111100111;
      patterns[7797] = 29'b0_001111001110_101_1_000011110011;
      patterns[7798] = 29'b0_001111001110_110_0_001111001110;
      patterns[7799] = 29'b0_001111001110_111_0_001111001110;
      patterns[7800] = 29'b0_001111001111_000_0_001111001111;
      patterns[7801] = 29'b0_001111001111_001_0_001111001111;
      patterns[7802] = 29'b0_001111001111_010_0_011110011110;
      patterns[7803] = 29'b0_001111001111_011_0_111100111100;
      patterns[7804] = 29'b0_001111001111_100_1_000111100111;
      patterns[7805] = 29'b0_001111001111_101_1_100011110011;
      patterns[7806] = 29'b0_001111001111_110_0_001111001111;
      patterns[7807] = 29'b0_001111001111_111_0_001111001111;
      patterns[7808] = 29'b0_001111010000_000_0_001111010000;
      patterns[7809] = 29'b0_001111010000_001_0_010000001111;
      patterns[7810] = 29'b0_001111010000_010_0_011110100000;
      patterns[7811] = 29'b0_001111010000_011_0_111101000000;
      patterns[7812] = 29'b0_001111010000_100_0_000111101000;
      patterns[7813] = 29'b0_001111010000_101_0_000011110100;
      patterns[7814] = 29'b0_001111010000_110_0_001111010000;
      patterns[7815] = 29'b0_001111010000_111_0_001111010000;
      patterns[7816] = 29'b0_001111010001_000_0_001111010001;
      patterns[7817] = 29'b0_001111010001_001_0_010001001111;
      patterns[7818] = 29'b0_001111010001_010_0_011110100010;
      patterns[7819] = 29'b0_001111010001_011_0_111101000100;
      patterns[7820] = 29'b0_001111010001_100_1_000111101000;
      patterns[7821] = 29'b0_001111010001_101_0_100011110100;
      patterns[7822] = 29'b0_001111010001_110_0_001111010001;
      patterns[7823] = 29'b0_001111010001_111_0_001111010001;
      patterns[7824] = 29'b0_001111010010_000_0_001111010010;
      patterns[7825] = 29'b0_001111010010_001_0_010010001111;
      patterns[7826] = 29'b0_001111010010_010_0_011110100100;
      patterns[7827] = 29'b0_001111010010_011_0_111101001000;
      patterns[7828] = 29'b0_001111010010_100_0_000111101001;
      patterns[7829] = 29'b0_001111010010_101_1_000011110100;
      patterns[7830] = 29'b0_001111010010_110_0_001111010010;
      patterns[7831] = 29'b0_001111010010_111_0_001111010010;
      patterns[7832] = 29'b0_001111010011_000_0_001111010011;
      patterns[7833] = 29'b0_001111010011_001_0_010011001111;
      patterns[7834] = 29'b0_001111010011_010_0_011110100110;
      patterns[7835] = 29'b0_001111010011_011_0_111101001100;
      patterns[7836] = 29'b0_001111010011_100_1_000111101001;
      patterns[7837] = 29'b0_001111010011_101_1_100011110100;
      patterns[7838] = 29'b0_001111010011_110_0_001111010011;
      patterns[7839] = 29'b0_001111010011_111_0_001111010011;
      patterns[7840] = 29'b0_001111010100_000_0_001111010100;
      patterns[7841] = 29'b0_001111010100_001_0_010100001111;
      patterns[7842] = 29'b0_001111010100_010_0_011110101000;
      patterns[7843] = 29'b0_001111010100_011_0_111101010000;
      patterns[7844] = 29'b0_001111010100_100_0_000111101010;
      patterns[7845] = 29'b0_001111010100_101_0_000011110101;
      patterns[7846] = 29'b0_001111010100_110_0_001111010100;
      patterns[7847] = 29'b0_001111010100_111_0_001111010100;
      patterns[7848] = 29'b0_001111010101_000_0_001111010101;
      patterns[7849] = 29'b0_001111010101_001_0_010101001111;
      patterns[7850] = 29'b0_001111010101_010_0_011110101010;
      patterns[7851] = 29'b0_001111010101_011_0_111101010100;
      patterns[7852] = 29'b0_001111010101_100_1_000111101010;
      patterns[7853] = 29'b0_001111010101_101_0_100011110101;
      patterns[7854] = 29'b0_001111010101_110_0_001111010101;
      patterns[7855] = 29'b0_001111010101_111_0_001111010101;
      patterns[7856] = 29'b0_001111010110_000_0_001111010110;
      patterns[7857] = 29'b0_001111010110_001_0_010110001111;
      patterns[7858] = 29'b0_001111010110_010_0_011110101100;
      patterns[7859] = 29'b0_001111010110_011_0_111101011000;
      patterns[7860] = 29'b0_001111010110_100_0_000111101011;
      patterns[7861] = 29'b0_001111010110_101_1_000011110101;
      patterns[7862] = 29'b0_001111010110_110_0_001111010110;
      patterns[7863] = 29'b0_001111010110_111_0_001111010110;
      patterns[7864] = 29'b0_001111010111_000_0_001111010111;
      patterns[7865] = 29'b0_001111010111_001_0_010111001111;
      patterns[7866] = 29'b0_001111010111_010_0_011110101110;
      patterns[7867] = 29'b0_001111010111_011_0_111101011100;
      patterns[7868] = 29'b0_001111010111_100_1_000111101011;
      patterns[7869] = 29'b0_001111010111_101_1_100011110101;
      patterns[7870] = 29'b0_001111010111_110_0_001111010111;
      patterns[7871] = 29'b0_001111010111_111_0_001111010111;
      patterns[7872] = 29'b0_001111011000_000_0_001111011000;
      patterns[7873] = 29'b0_001111011000_001_0_011000001111;
      patterns[7874] = 29'b0_001111011000_010_0_011110110000;
      patterns[7875] = 29'b0_001111011000_011_0_111101100000;
      patterns[7876] = 29'b0_001111011000_100_0_000111101100;
      patterns[7877] = 29'b0_001111011000_101_0_000011110110;
      patterns[7878] = 29'b0_001111011000_110_0_001111011000;
      patterns[7879] = 29'b0_001111011000_111_0_001111011000;
      patterns[7880] = 29'b0_001111011001_000_0_001111011001;
      patterns[7881] = 29'b0_001111011001_001_0_011001001111;
      patterns[7882] = 29'b0_001111011001_010_0_011110110010;
      patterns[7883] = 29'b0_001111011001_011_0_111101100100;
      patterns[7884] = 29'b0_001111011001_100_1_000111101100;
      patterns[7885] = 29'b0_001111011001_101_0_100011110110;
      patterns[7886] = 29'b0_001111011001_110_0_001111011001;
      patterns[7887] = 29'b0_001111011001_111_0_001111011001;
      patterns[7888] = 29'b0_001111011010_000_0_001111011010;
      patterns[7889] = 29'b0_001111011010_001_0_011010001111;
      patterns[7890] = 29'b0_001111011010_010_0_011110110100;
      patterns[7891] = 29'b0_001111011010_011_0_111101101000;
      patterns[7892] = 29'b0_001111011010_100_0_000111101101;
      patterns[7893] = 29'b0_001111011010_101_1_000011110110;
      patterns[7894] = 29'b0_001111011010_110_0_001111011010;
      patterns[7895] = 29'b0_001111011010_111_0_001111011010;
      patterns[7896] = 29'b0_001111011011_000_0_001111011011;
      patterns[7897] = 29'b0_001111011011_001_0_011011001111;
      patterns[7898] = 29'b0_001111011011_010_0_011110110110;
      patterns[7899] = 29'b0_001111011011_011_0_111101101100;
      patterns[7900] = 29'b0_001111011011_100_1_000111101101;
      patterns[7901] = 29'b0_001111011011_101_1_100011110110;
      patterns[7902] = 29'b0_001111011011_110_0_001111011011;
      patterns[7903] = 29'b0_001111011011_111_0_001111011011;
      patterns[7904] = 29'b0_001111011100_000_0_001111011100;
      patterns[7905] = 29'b0_001111011100_001_0_011100001111;
      patterns[7906] = 29'b0_001111011100_010_0_011110111000;
      patterns[7907] = 29'b0_001111011100_011_0_111101110000;
      patterns[7908] = 29'b0_001111011100_100_0_000111101110;
      patterns[7909] = 29'b0_001111011100_101_0_000011110111;
      patterns[7910] = 29'b0_001111011100_110_0_001111011100;
      patterns[7911] = 29'b0_001111011100_111_0_001111011100;
      patterns[7912] = 29'b0_001111011101_000_0_001111011101;
      patterns[7913] = 29'b0_001111011101_001_0_011101001111;
      patterns[7914] = 29'b0_001111011101_010_0_011110111010;
      patterns[7915] = 29'b0_001111011101_011_0_111101110100;
      patterns[7916] = 29'b0_001111011101_100_1_000111101110;
      patterns[7917] = 29'b0_001111011101_101_0_100011110111;
      patterns[7918] = 29'b0_001111011101_110_0_001111011101;
      patterns[7919] = 29'b0_001111011101_111_0_001111011101;
      patterns[7920] = 29'b0_001111011110_000_0_001111011110;
      patterns[7921] = 29'b0_001111011110_001_0_011110001111;
      patterns[7922] = 29'b0_001111011110_010_0_011110111100;
      patterns[7923] = 29'b0_001111011110_011_0_111101111000;
      patterns[7924] = 29'b0_001111011110_100_0_000111101111;
      patterns[7925] = 29'b0_001111011110_101_1_000011110111;
      patterns[7926] = 29'b0_001111011110_110_0_001111011110;
      patterns[7927] = 29'b0_001111011110_111_0_001111011110;
      patterns[7928] = 29'b0_001111011111_000_0_001111011111;
      patterns[7929] = 29'b0_001111011111_001_0_011111001111;
      patterns[7930] = 29'b0_001111011111_010_0_011110111110;
      patterns[7931] = 29'b0_001111011111_011_0_111101111100;
      patterns[7932] = 29'b0_001111011111_100_1_000111101111;
      patterns[7933] = 29'b0_001111011111_101_1_100011110111;
      patterns[7934] = 29'b0_001111011111_110_0_001111011111;
      patterns[7935] = 29'b0_001111011111_111_0_001111011111;
      patterns[7936] = 29'b0_001111100000_000_0_001111100000;
      patterns[7937] = 29'b0_001111100000_001_0_100000001111;
      patterns[7938] = 29'b0_001111100000_010_0_011111000000;
      patterns[7939] = 29'b0_001111100000_011_0_111110000000;
      patterns[7940] = 29'b0_001111100000_100_0_000111110000;
      patterns[7941] = 29'b0_001111100000_101_0_000011111000;
      patterns[7942] = 29'b0_001111100000_110_0_001111100000;
      patterns[7943] = 29'b0_001111100000_111_0_001111100000;
      patterns[7944] = 29'b0_001111100001_000_0_001111100001;
      patterns[7945] = 29'b0_001111100001_001_0_100001001111;
      patterns[7946] = 29'b0_001111100001_010_0_011111000010;
      patterns[7947] = 29'b0_001111100001_011_0_111110000100;
      patterns[7948] = 29'b0_001111100001_100_1_000111110000;
      patterns[7949] = 29'b0_001111100001_101_0_100011111000;
      patterns[7950] = 29'b0_001111100001_110_0_001111100001;
      patterns[7951] = 29'b0_001111100001_111_0_001111100001;
      patterns[7952] = 29'b0_001111100010_000_0_001111100010;
      patterns[7953] = 29'b0_001111100010_001_0_100010001111;
      patterns[7954] = 29'b0_001111100010_010_0_011111000100;
      patterns[7955] = 29'b0_001111100010_011_0_111110001000;
      patterns[7956] = 29'b0_001111100010_100_0_000111110001;
      patterns[7957] = 29'b0_001111100010_101_1_000011111000;
      patterns[7958] = 29'b0_001111100010_110_0_001111100010;
      patterns[7959] = 29'b0_001111100010_111_0_001111100010;
      patterns[7960] = 29'b0_001111100011_000_0_001111100011;
      patterns[7961] = 29'b0_001111100011_001_0_100011001111;
      patterns[7962] = 29'b0_001111100011_010_0_011111000110;
      patterns[7963] = 29'b0_001111100011_011_0_111110001100;
      patterns[7964] = 29'b0_001111100011_100_1_000111110001;
      patterns[7965] = 29'b0_001111100011_101_1_100011111000;
      patterns[7966] = 29'b0_001111100011_110_0_001111100011;
      patterns[7967] = 29'b0_001111100011_111_0_001111100011;
      patterns[7968] = 29'b0_001111100100_000_0_001111100100;
      patterns[7969] = 29'b0_001111100100_001_0_100100001111;
      patterns[7970] = 29'b0_001111100100_010_0_011111001000;
      patterns[7971] = 29'b0_001111100100_011_0_111110010000;
      patterns[7972] = 29'b0_001111100100_100_0_000111110010;
      patterns[7973] = 29'b0_001111100100_101_0_000011111001;
      patterns[7974] = 29'b0_001111100100_110_0_001111100100;
      patterns[7975] = 29'b0_001111100100_111_0_001111100100;
      patterns[7976] = 29'b0_001111100101_000_0_001111100101;
      patterns[7977] = 29'b0_001111100101_001_0_100101001111;
      patterns[7978] = 29'b0_001111100101_010_0_011111001010;
      patterns[7979] = 29'b0_001111100101_011_0_111110010100;
      patterns[7980] = 29'b0_001111100101_100_1_000111110010;
      patterns[7981] = 29'b0_001111100101_101_0_100011111001;
      patterns[7982] = 29'b0_001111100101_110_0_001111100101;
      patterns[7983] = 29'b0_001111100101_111_0_001111100101;
      patterns[7984] = 29'b0_001111100110_000_0_001111100110;
      patterns[7985] = 29'b0_001111100110_001_0_100110001111;
      patterns[7986] = 29'b0_001111100110_010_0_011111001100;
      patterns[7987] = 29'b0_001111100110_011_0_111110011000;
      patterns[7988] = 29'b0_001111100110_100_0_000111110011;
      patterns[7989] = 29'b0_001111100110_101_1_000011111001;
      patterns[7990] = 29'b0_001111100110_110_0_001111100110;
      patterns[7991] = 29'b0_001111100110_111_0_001111100110;
      patterns[7992] = 29'b0_001111100111_000_0_001111100111;
      patterns[7993] = 29'b0_001111100111_001_0_100111001111;
      patterns[7994] = 29'b0_001111100111_010_0_011111001110;
      patterns[7995] = 29'b0_001111100111_011_0_111110011100;
      patterns[7996] = 29'b0_001111100111_100_1_000111110011;
      patterns[7997] = 29'b0_001111100111_101_1_100011111001;
      patterns[7998] = 29'b0_001111100111_110_0_001111100111;
      patterns[7999] = 29'b0_001111100111_111_0_001111100111;
      patterns[8000] = 29'b0_001111101000_000_0_001111101000;
      patterns[8001] = 29'b0_001111101000_001_0_101000001111;
      patterns[8002] = 29'b0_001111101000_010_0_011111010000;
      patterns[8003] = 29'b0_001111101000_011_0_111110100000;
      patterns[8004] = 29'b0_001111101000_100_0_000111110100;
      patterns[8005] = 29'b0_001111101000_101_0_000011111010;
      patterns[8006] = 29'b0_001111101000_110_0_001111101000;
      patterns[8007] = 29'b0_001111101000_111_0_001111101000;
      patterns[8008] = 29'b0_001111101001_000_0_001111101001;
      patterns[8009] = 29'b0_001111101001_001_0_101001001111;
      patterns[8010] = 29'b0_001111101001_010_0_011111010010;
      patterns[8011] = 29'b0_001111101001_011_0_111110100100;
      patterns[8012] = 29'b0_001111101001_100_1_000111110100;
      patterns[8013] = 29'b0_001111101001_101_0_100011111010;
      patterns[8014] = 29'b0_001111101001_110_0_001111101001;
      patterns[8015] = 29'b0_001111101001_111_0_001111101001;
      patterns[8016] = 29'b0_001111101010_000_0_001111101010;
      patterns[8017] = 29'b0_001111101010_001_0_101010001111;
      patterns[8018] = 29'b0_001111101010_010_0_011111010100;
      patterns[8019] = 29'b0_001111101010_011_0_111110101000;
      patterns[8020] = 29'b0_001111101010_100_0_000111110101;
      patterns[8021] = 29'b0_001111101010_101_1_000011111010;
      patterns[8022] = 29'b0_001111101010_110_0_001111101010;
      patterns[8023] = 29'b0_001111101010_111_0_001111101010;
      patterns[8024] = 29'b0_001111101011_000_0_001111101011;
      patterns[8025] = 29'b0_001111101011_001_0_101011001111;
      patterns[8026] = 29'b0_001111101011_010_0_011111010110;
      patterns[8027] = 29'b0_001111101011_011_0_111110101100;
      patterns[8028] = 29'b0_001111101011_100_1_000111110101;
      patterns[8029] = 29'b0_001111101011_101_1_100011111010;
      patterns[8030] = 29'b0_001111101011_110_0_001111101011;
      patterns[8031] = 29'b0_001111101011_111_0_001111101011;
      patterns[8032] = 29'b0_001111101100_000_0_001111101100;
      patterns[8033] = 29'b0_001111101100_001_0_101100001111;
      patterns[8034] = 29'b0_001111101100_010_0_011111011000;
      patterns[8035] = 29'b0_001111101100_011_0_111110110000;
      patterns[8036] = 29'b0_001111101100_100_0_000111110110;
      patterns[8037] = 29'b0_001111101100_101_0_000011111011;
      patterns[8038] = 29'b0_001111101100_110_0_001111101100;
      patterns[8039] = 29'b0_001111101100_111_0_001111101100;
      patterns[8040] = 29'b0_001111101101_000_0_001111101101;
      patterns[8041] = 29'b0_001111101101_001_0_101101001111;
      patterns[8042] = 29'b0_001111101101_010_0_011111011010;
      patterns[8043] = 29'b0_001111101101_011_0_111110110100;
      patterns[8044] = 29'b0_001111101101_100_1_000111110110;
      patterns[8045] = 29'b0_001111101101_101_0_100011111011;
      patterns[8046] = 29'b0_001111101101_110_0_001111101101;
      patterns[8047] = 29'b0_001111101101_111_0_001111101101;
      patterns[8048] = 29'b0_001111101110_000_0_001111101110;
      patterns[8049] = 29'b0_001111101110_001_0_101110001111;
      patterns[8050] = 29'b0_001111101110_010_0_011111011100;
      patterns[8051] = 29'b0_001111101110_011_0_111110111000;
      patterns[8052] = 29'b0_001111101110_100_0_000111110111;
      patterns[8053] = 29'b0_001111101110_101_1_000011111011;
      patterns[8054] = 29'b0_001111101110_110_0_001111101110;
      patterns[8055] = 29'b0_001111101110_111_0_001111101110;
      patterns[8056] = 29'b0_001111101111_000_0_001111101111;
      patterns[8057] = 29'b0_001111101111_001_0_101111001111;
      patterns[8058] = 29'b0_001111101111_010_0_011111011110;
      patterns[8059] = 29'b0_001111101111_011_0_111110111100;
      patterns[8060] = 29'b0_001111101111_100_1_000111110111;
      patterns[8061] = 29'b0_001111101111_101_1_100011111011;
      patterns[8062] = 29'b0_001111101111_110_0_001111101111;
      patterns[8063] = 29'b0_001111101111_111_0_001111101111;
      patterns[8064] = 29'b0_001111110000_000_0_001111110000;
      patterns[8065] = 29'b0_001111110000_001_0_110000001111;
      patterns[8066] = 29'b0_001111110000_010_0_011111100000;
      patterns[8067] = 29'b0_001111110000_011_0_111111000000;
      patterns[8068] = 29'b0_001111110000_100_0_000111111000;
      patterns[8069] = 29'b0_001111110000_101_0_000011111100;
      patterns[8070] = 29'b0_001111110000_110_0_001111110000;
      patterns[8071] = 29'b0_001111110000_111_0_001111110000;
      patterns[8072] = 29'b0_001111110001_000_0_001111110001;
      patterns[8073] = 29'b0_001111110001_001_0_110001001111;
      patterns[8074] = 29'b0_001111110001_010_0_011111100010;
      patterns[8075] = 29'b0_001111110001_011_0_111111000100;
      patterns[8076] = 29'b0_001111110001_100_1_000111111000;
      patterns[8077] = 29'b0_001111110001_101_0_100011111100;
      patterns[8078] = 29'b0_001111110001_110_0_001111110001;
      patterns[8079] = 29'b0_001111110001_111_0_001111110001;
      patterns[8080] = 29'b0_001111110010_000_0_001111110010;
      patterns[8081] = 29'b0_001111110010_001_0_110010001111;
      patterns[8082] = 29'b0_001111110010_010_0_011111100100;
      patterns[8083] = 29'b0_001111110010_011_0_111111001000;
      patterns[8084] = 29'b0_001111110010_100_0_000111111001;
      patterns[8085] = 29'b0_001111110010_101_1_000011111100;
      patterns[8086] = 29'b0_001111110010_110_0_001111110010;
      patterns[8087] = 29'b0_001111110010_111_0_001111110010;
      patterns[8088] = 29'b0_001111110011_000_0_001111110011;
      patterns[8089] = 29'b0_001111110011_001_0_110011001111;
      patterns[8090] = 29'b0_001111110011_010_0_011111100110;
      patterns[8091] = 29'b0_001111110011_011_0_111111001100;
      patterns[8092] = 29'b0_001111110011_100_1_000111111001;
      patterns[8093] = 29'b0_001111110011_101_1_100011111100;
      patterns[8094] = 29'b0_001111110011_110_0_001111110011;
      patterns[8095] = 29'b0_001111110011_111_0_001111110011;
      patterns[8096] = 29'b0_001111110100_000_0_001111110100;
      patterns[8097] = 29'b0_001111110100_001_0_110100001111;
      patterns[8098] = 29'b0_001111110100_010_0_011111101000;
      patterns[8099] = 29'b0_001111110100_011_0_111111010000;
      patterns[8100] = 29'b0_001111110100_100_0_000111111010;
      patterns[8101] = 29'b0_001111110100_101_0_000011111101;
      patterns[8102] = 29'b0_001111110100_110_0_001111110100;
      patterns[8103] = 29'b0_001111110100_111_0_001111110100;
      patterns[8104] = 29'b0_001111110101_000_0_001111110101;
      patterns[8105] = 29'b0_001111110101_001_0_110101001111;
      patterns[8106] = 29'b0_001111110101_010_0_011111101010;
      patterns[8107] = 29'b0_001111110101_011_0_111111010100;
      patterns[8108] = 29'b0_001111110101_100_1_000111111010;
      patterns[8109] = 29'b0_001111110101_101_0_100011111101;
      patterns[8110] = 29'b0_001111110101_110_0_001111110101;
      patterns[8111] = 29'b0_001111110101_111_0_001111110101;
      patterns[8112] = 29'b0_001111110110_000_0_001111110110;
      patterns[8113] = 29'b0_001111110110_001_0_110110001111;
      patterns[8114] = 29'b0_001111110110_010_0_011111101100;
      patterns[8115] = 29'b0_001111110110_011_0_111111011000;
      patterns[8116] = 29'b0_001111110110_100_0_000111111011;
      patterns[8117] = 29'b0_001111110110_101_1_000011111101;
      patterns[8118] = 29'b0_001111110110_110_0_001111110110;
      patterns[8119] = 29'b0_001111110110_111_0_001111110110;
      patterns[8120] = 29'b0_001111110111_000_0_001111110111;
      patterns[8121] = 29'b0_001111110111_001_0_110111001111;
      patterns[8122] = 29'b0_001111110111_010_0_011111101110;
      patterns[8123] = 29'b0_001111110111_011_0_111111011100;
      patterns[8124] = 29'b0_001111110111_100_1_000111111011;
      patterns[8125] = 29'b0_001111110111_101_1_100011111101;
      patterns[8126] = 29'b0_001111110111_110_0_001111110111;
      patterns[8127] = 29'b0_001111110111_111_0_001111110111;
      patterns[8128] = 29'b0_001111111000_000_0_001111111000;
      patterns[8129] = 29'b0_001111111000_001_0_111000001111;
      patterns[8130] = 29'b0_001111111000_010_0_011111110000;
      patterns[8131] = 29'b0_001111111000_011_0_111111100000;
      patterns[8132] = 29'b0_001111111000_100_0_000111111100;
      patterns[8133] = 29'b0_001111111000_101_0_000011111110;
      patterns[8134] = 29'b0_001111111000_110_0_001111111000;
      patterns[8135] = 29'b0_001111111000_111_0_001111111000;
      patterns[8136] = 29'b0_001111111001_000_0_001111111001;
      patterns[8137] = 29'b0_001111111001_001_0_111001001111;
      patterns[8138] = 29'b0_001111111001_010_0_011111110010;
      patterns[8139] = 29'b0_001111111001_011_0_111111100100;
      patterns[8140] = 29'b0_001111111001_100_1_000111111100;
      patterns[8141] = 29'b0_001111111001_101_0_100011111110;
      patterns[8142] = 29'b0_001111111001_110_0_001111111001;
      patterns[8143] = 29'b0_001111111001_111_0_001111111001;
      patterns[8144] = 29'b0_001111111010_000_0_001111111010;
      patterns[8145] = 29'b0_001111111010_001_0_111010001111;
      patterns[8146] = 29'b0_001111111010_010_0_011111110100;
      patterns[8147] = 29'b0_001111111010_011_0_111111101000;
      patterns[8148] = 29'b0_001111111010_100_0_000111111101;
      patterns[8149] = 29'b0_001111111010_101_1_000011111110;
      patterns[8150] = 29'b0_001111111010_110_0_001111111010;
      patterns[8151] = 29'b0_001111111010_111_0_001111111010;
      patterns[8152] = 29'b0_001111111011_000_0_001111111011;
      patterns[8153] = 29'b0_001111111011_001_0_111011001111;
      patterns[8154] = 29'b0_001111111011_010_0_011111110110;
      patterns[8155] = 29'b0_001111111011_011_0_111111101100;
      patterns[8156] = 29'b0_001111111011_100_1_000111111101;
      patterns[8157] = 29'b0_001111111011_101_1_100011111110;
      patterns[8158] = 29'b0_001111111011_110_0_001111111011;
      patterns[8159] = 29'b0_001111111011_111_0_001111111011;
      patterns[8160] = 29'b0_001111111100_000_0_001111111100;
      patterns[8161] = 29'b0_001111111100_001_0_111100001111;
      patterns[8162] = 29'b0_001111111100_010_0_011111111000;
      patterns[8163] = 29'b0_001111111100_011_0_111111110000;
      patterns[8164] = 29'b0_001111111100_100_0_000111111110;
      patterns[8165] = 29'b0_001111111100_101_0_000011111111;
      patterns[8166] = 29'b0_001111111100_110_0_001111111100;
      patterns[8167] = 29'b0_001111111100_111_0_001111111100;
      patterns[8168] = 29'b0_001111111101_000_0_001111111101;
      patterns[8169] = 29'b0_001111111101_001_0_111101001111;
      patterns[8170] = 29'b0_001111111101_010_0_011111111010;
      patterns[8171] = 29'b0_001111111101_011_0_111111110100;
      patterns[8172] = 29'b0_001111111101_100_1_000111111110;
      patterns[8173] = 29'b0_001111111101_101_0_100011111111;
      patterns[8174] = 29'b0_001111111101_110_0_001111111101;
      patterns[8175] = 29'b0_001111111101_111_0_001111111101;
      patterns[8176] = 29'b0_001111111110_000_0_001111111110;
      patterns[8177] = 29'b0_001111111110_001_0_111110001111;
      patterns[8178] = 29'b0_001111111110_010_0_011111111100;
      patterns[8179] = 29'b0_001111111110_011_0_111111111000;
      patterns[8180] = 29'b0_001111111110_100_0_000111111111;
      patterns[8181] = 29'b0_001111111110_101_1_000011111111;
      patterns[8182] = 29'b0_001111111110_110_0_001111111110;
      patterns[8183] = 29'b0_001111111110_111_0_001111111110;
      patterns[8184] = 29'b0_001111111111_000_0_001111111111;
      patterns[8185] = 29'b0_001111111111_001_0_111111001111;
      patterns[8186] = 29'b0_001111111111_010_0_011111111110;
      patterns[8187] = 29'b0_001111111111_011_0_111111111100;
      patterns[8188] = 29'b0_001111111111_100_1_000111111111;
      patterns[8189] = 29'b0_001111111111_101_1_100011111111;
      patterns[8190] = 29'b0_001111111111_110_0_001111111111;
      patterns[8191] = 29'b0_001111111111_111_0_001111111111;
      patterns[8192] = 29'b0_010000000000_000_0_010000000000;
      patterns[8193] = 29'b0_010000000000_001_0_000000010000;
      patterns[8194] = 29'b0_010000000000_010_0_100000000000;
      patterns[8195] = 29'b0_010000000000_011_1_000000000000;
      patterns[8196] = 29'b0_010000000000_100_0_001000000000;
      patterns[8197] = 29'b0_010000000000_101_0_000100000000;
      patterns[8198] = 29'b0_010000000000_110_0_010000000000;
      patterns[8199] = 29'b0_010000000000_111_0_010000000000;
      patterns[8200] = 29'b0_010000000001_000_0_010000000001;
      patterns[8201] = 29'b0_010000000001_001_0_000001010000;
      patterns[8202] = 29'b0_010000000001_010_0_100000000010;
      patterns[8203] = 29'b0_010000000001_011_1_000000000100;
      patterns[8204] = 29'b0_010000000001_100_1_001000000000;
      patterns[8205] = 29'b0_010000000001_101_0_100100000000;
      patterns[8206] = 29'b0_010000000001_110_0_010000000001;
      patterns[8207] = 29'b0_010000000001_111_0_010000000001;
      patterns[8208] = 29'b0_010000000010_000_0_010000000010;
      patterns[8209] = 29'b0_010000000010_001_0_000010010000;
      patterns[8210] = 29'b0_010000000010_010_0_100000000100;
      patterns[8211] = 29'b0_010000000010_011_1_000000001000;
      patterns[8212] = 29'b0_010000000010_100_0_001000000001;
      patterns[8213] = 29'b0_010000000010_101_1_000100000000;
      patterns[8214] = 29'b0_010000000010_110_0_010000000010;
      patterns[8215] = 29'b0_010000000010_111_0_010000000010;
      patterns[8216] = 29'b0_010000000011_000_0_010000000011;
      patterns[8217] = 29'b0_010000000011_001_0_000011010000;
      patterns[8218] = 29'b0_010000000011_010_0_100000000110;
      patterns[8219] = 29'b0_010000000011_011_1_000000001100;
      patterns[8220] = 29'b0_010000000011_100_1_001000000001;
      patterns[8221] = 29'b0_010000000011_101_1_100100000000;
      patterns[8222] = 29'b0_010000000011_110_0_010000000011;
      patterns[8223] = 29'b0_010000000011_111_0_010000000011;
      patterns[8224] = 29'b0_010000000100_000_0_010000000100;
      patterns[8225] = 29'b0_010000000100_001_0_000100010000;
      patterns[8226] = 29'b0_010000000100_010_0_100000001000;
      patterns[8227] = 29'b0_010000000100_011_1_000000010000;
      patterns[8228] = 29'b0_010000000100_100_0_001000000010;
      patterns[8229] = 29'b0_010000000100_101_0_000100000001;
      patterns[8230] = 29'b0_010000000100_110_0_010000000100;
      patterns[8231] = 29'b0_010000000100_111_0_010000000100;
      patterns[8232] = 29'b0_010000000101_000_0_010000000101;
      patterns[8233] = 29'b0_010000000101_001_0_000101010000;
      patterns[8234] = 29'b0_010000000101_010_0_100000001010;
      patterns[8235] = 29'b0_010000000101_011_1_000000010100;
      patterns[8236] = 29'b0_010000000101_100_1_001000000010;
      patterns[8237] = 29'b0_010000000101_101_0_100100000001;
      patterns[8238] = 29'b0_010000000101_110_0_010000000101;
      patterns[8239] = 29'b0_010000000101_111_0_010000000101;
      patterns[8240] = 29'b0_010000000110_000_0_010000000110;
      patterns[8241] = 29'b0_010000000110_001_0_000110010000;
      patterns[8242] = 29'b0_010000000110_010_0_100000001100;
      patterns[8243] = 29'b0_010000000110_011_1_000000011000;
      patterns[8244] = 29'b0_010000000110_100_0_001000000011;
      patterns[8245] = 29'b0_010000000110_101_1_000100000001;
      patterns[8246] = 29'b0_010000000110_110_0_010000000110;
      patterns[8247] = 29'b0_010000000110_111_0_010000000110;
      patterns[8248] = 29'b0_010000000111_000_0_010000000111;
      patterns[8249] = 29'b0_010000000111_001_0_000111010000;
      patterns[8250] = 29'b0_010000000111_010_0_100000001110;
      patterns[8251] = 29'b0_010000000111_011_1_000000011100;
      patterns[8252] = 29'b0_010000000111_100_1_001000000011;
      patterns[8253] = 29'b0_010000000111_101_1_100100000001;
      patterns[8254] = 29'b0_010000000111_110_0_010000000111;
      patterns[8255] = 29'b0_010000000111_111_0_010000000111;
      patterns[8256] = 29'b0_010000001000_000_0_010000001000;
      patterns[8257] = 29'b0_010000001000_001_0_001000010000;
      patterns[8258] = 29'b0_010000001000_010_0_100000010000;
      patterns[8259] = 29'b0_010000001000_011_1_000000100000;
      patterns[8260] = 29'b0_010000001000_100_0_001000000100;
      patterns[8261] = 29'b0_010000001000_101_0_000100000010;
      patterns[8262] = 29'b0_010000001000_110_0_010000001000;
      patterns[8263] = 29'b0_010000001000_111_0_010000001000;
      patterns[8264] = 29'b0_010000001001_000_0_010000001001;
      patterns[8265] = 29'b0_010000001001_001_0_001001010000;
      patterns[8266] = 29'b0_010000001001_010_0_100000010010;
      patterns[8267] = 29'b0_010000001001_011_1_000000100100;
      patterns[8268] = 29'b0_010000001001_100_1_001000000100;
      patterns[8269] = 29'b0_010000001001_101_0_100100000010;
      patterns[8270] = 29'b0_010000001001_110_0_010000001001;
      patterns[8271] = 29'b0_010000001001_111_0_010000001001;
      patterns[8272] = 29'b0_010000001010_000_0_010000001010;
      patterns[8273] = 29'b0_010000001010_001_0_001010010000;
      patterns[8274] = 29'b0_010000001010_010_0_100000010100;
      patterns[8275] = 29'b0_010000001010_011_1_000000101000;
      patterns[8276] = 29'b0_010000001010_100_0_001000000101;
      patterns[8277] = 29'b0_010000001010_101_1_000100000010;
      patterns[8278] = 29'b0_010000001010_110_0_010000001010;
      patterns[8279] = 29'b0_010000001010_111_0_010000001010;
      patterns[8280] = 29'b0_010000001011_000_0_010000001011;
      patterns[8281] = 29'b0_010000001011_001_0_001011010000;
      patterns[8282] = 29'b0_010000001011_010_0_100000010110;
      patterns[8283] = 29'b0_010000001011_011_1_000000101100;
      patterns[8284] = 29'b0_010000001011_100_1_001000000101;
      patterns[8285] = 29'b0_010000001011_101_1_100100000010;
      patterns[8286] = 29'b0_010000001011_110_0_010000001011;
      patterns[8287] = 29'b0_010000001011_111_0_010000001011;
      patterns[8288] = 29'b0_010000001100_000_0_010000001100;
      patterns[8289] = 29'b0_010000001100_001_0_001100010000;
      patterns[8290] = 29'b0_010000001100_010_0_100000011000;
      patterns[8291] = 29'b0_010000001100_011_1_000000110000;
      patterns[8292] = 29'b0_010000001100_100_0_001000000110;
      patterns[8293] = 29'b0_010000001100_101_0_000100000011;
      patterns[8294] = 29'b0_010000001100_110_0_010000001100;
      patterns[8295] = 29'b0_010000001100_111_0_010000001100;
      patterns[8296] = 29'b0_010000001101_000_0_010000001101;
      patterns[8297] = 29'b0_010000001101_001_0_001101010000;
      patterns[8298] = 29'b0_010000001101_010_0_100000011010;
      patterns[8299] = 29'b0_010000001101_011_1_000000110100;
      patterns[8300] = 29'b0_010000001101_100_1_001000000110;
      patterns[8301] = 29'b0_010000001101_101_0_100100000011;
      patterns[8302] = 29'b0_010000001101_110_0_010000001101;
      patterns[8303] = 29'b0_010000001101_111_0_010000001101;
      patterns[8304] = 29'b0_010000001110_000_0_010000001110;
      patterns[8305] = 29'b0_010000001110_001_0_001110010000;
      patterns[8306] = 29'b0_010000001110_010_0_100000011100;
      patterns[8307] = 29'b0_010000001110_011_1_000000111000;
      patterns[8308] = 29'b0_010000001110_100_0_001000000111;
      patterns[8309] = 29'b0_010000001110_101_1_000100000011;
      patterns[8310] = 29'b0_010000001110_110_0_010000001110;
      patterns[8311] = 29'b0_010000001110_111_0_010000001110;
      patterns[8312] = 29'b0_010000001111_000_0_010000001111;
      patterns[8313] = 29'b0_010000001111_001_0_001111010000;
      patterns[8314] = 29'b0_010000001111_010_0_100000011110;
      patterns[8315] = 29'b0_010000001111_011_1_000000111100;
      patterns[8316] = 29'b0_010000001111_100_1_001000000111;
      patterns[8317] = 29'b0_010000001111_101_1_100100000011;
      patterns[8318] = 29'b0_010000001111_110_0_010000001111;
      patterns[8319] = 29'b0_010000001111_111_0_010000001111;
      patterns[8320] = 29'b0_010000010000_000_0_010000010000;
      patterns[8321] = 29'b0_010000010000_001_0_010000010000;
      patterns[8322] = 29'b0_010000010000_010_0_100000100000;
      patterns[8323] = 29'b0_010000010000_011_1_000001000000;
      patterns[8324] = 29'b0_010000010000_100_0_001000001000;
      patterns[8325] = 29'b0_010000010000_101_0_000100000100;
      patterns[8326] = 29'b0_010000010000_110_0_010000010000;
      patterns[8327] = 29'b0_010000010000_111_0_010000010000;
      patterns[8328] = 29'b0_010000010001_000_0_010000010001;
      patterns[8329] = 29'b0_010000010001_001_0_010001010000;
      patterns[8330] = 29'b0_010000010001_010_0_100000100010;
      patterns[8331] = 29'b0_010000010001_011_1_000001000100;
      patterns[8332] = 29'b0_010000010001_100_1_001000001000;
      patterns[8333] = 29'b0_010000010001_101_0_100100000100;
      patterns[8334] = 29'b0_010000010001_110_0_010000010001;
      patterns[8335] = 29'b0_010000010001_111_0_010000010001;
      patterns[8336] = 29'b0_010000010010_000_0_010000010010;
      patterns[8337] = 29'b0_010000010010_001_0_010010010000;
      patterns[8338] = 29'b0_010000010010_010_0_100000100100;
      patterns[8339] = 29'b0_010000010010_011_1_000001001000;
      patterns[8340] = 29'b0_010000010010_100_0_001000001001;
      patterns[8341] = 29'b0_010000010010_101_1_000100000100;
      patterns[8342] = 29'b0_010000010010_110_0_010000010010;
      patterns[8343] = 29'b0_010000010010_111_0_010000010010;
      patterns[8344] = 29'b0_010000010011_000_0_010000010011;
      patterns[8345] = 29'b0_010000010011_001_0_010011010000;
      patterns[8346] = 29'b0_010000010011_010_0_100000100110;
      patterns[8347] = 29'b0_010000010011_011_1_000001001100;
      patterns[8348] = 29'b0_010000010011_100_1_001000001001;
      patterns[8349] = 29'b0_010000010011_101_1_100100000100;
      patterns[8350] = 29'b0_010000010011_110_0_010000010011;
      patterns[8351] = 29'b0_010000010011_111_0_010000010011;
      patterns[8352] = 29'b0_010000010100_000_0_010000010100;
      patterns[8353] = 29'b0_010000010100_001_0_010100010000;
      patterns[8354] = 29'b0_010000010100_010_0_100000101000;
      patterns[8355] = 29'b0_010000010100_011_1_000001010000;
      patterns[8356] = 29'b0_010000010100_100_0_001000001010;
      patterns[8357] = 29'b0_010000010100_101_0_000100000101;
      patterns[8358] = 29'b0_010000010100_110_0_010000010100;
      patterns[8359] = 29'b0_010000010100_111_0_010000010100;
      patterns[8360] = 29'b0_010000010101_000_0_010000010101;
      patterns[8361] = 29'b0_010000010101_001_0_010101010000;
      patterns[8362] = 29'b0_010000010101_010_0_100000101010;
      patterns[8363] = 29'b0_010000010101_011_1_000001010100;
      patterns[8364] = 29'b0_010000010101_100_1_001000001010;
      patterns[8365] = 29'b0_010000010101_101_0_100100000101;
      patterns[8366] = 29'b0_010000010101_110_0_010000010101;
      patterns[8367] = 29'b0_010000010101_111_0_010000010101;
      patterns[8368] = 29'b0_010000010110_000_0_010000010110;
      patterns[8369] = 29'b0_010000010110_001_0_010110010000;
      patterns[8370] = 29'b0_010000010110_010_0_100000101100;
      patterns[8371] = 29'b0_010000010110_011_1_000001011000;
      patterns[8372] = 29'b0_010000010110_100_0_001000001011;
      patterns[8373] = 29'b0_010000010110_101_1_000100000101;
      patterns[8374] = 29'b0_010000010110_110_0_010000010110;
      patterns[8375] = 29'b0_010000010110_111_0_010000010110;
      patterns[8376] = 29'b0_010000010111_000_0_010000010111;
      patterns[8377] = 29'b0_010000010111_001_0_010111010000;
      patterns[8378] = 29'b0_010000010111_010_0_100000101110;
      patterns[8379] = 29'b0_010000010111_011_1_000001011100;
      patterns[8380] = 29'b0_010000010111_100_1_001000001011;
      patterns[8381] = 29'b0_010000010111_101_1_100100000101;
      patterns[8382] = 29'b0_010000010111_110_0_010000010111;
      patterns[8383] = 29'b0_010000010111_111_0_010000010111;
      patterns[8384] = 29'b0_010000011000_000_0_010000011000;
      patterns[8385] = 29'b0_010000011000_001_0_011000010000;
      patterns[8386] = 29'b0_010000011000_010_0_100000110000;
      patterns[8387] = 29'b0_010000011000_011_1_000001100000;
      patterns[8388] = 29'b0_010000011000_100_0_001000001100;
      patterns[8389] = 29'b0_010000011000_101_0_000100000110;
      patterns[8390] = 29'b0_010000011000_110_0_010000011000;
      patterns[8391] = 29'b0_010000011000_111_0_010000011000;
      patterns[8392] = 29'b0_010000011001_000_0_010000011001;
      patterns[8393] = 29'b0_010000011001_001_0_011001010000;
      patterns[8394] = 29'b0_010000011001_010_0_100000110010;
      patterns[8395] = 29'b0_010000011001_011_1_000001100100;
      patterns[8396] = 29'b0_010000011001_100_1_001000001100;
      patterns[8397] = 29'b0_010000011001_101_0_100100000110;
      patterns[8398] = 29'b0_010000011001_110_0_010000011001;
      patterns[8399] = 29'b0_010000011001_111_0_010000011001;
      patterns[8400] = 29'b0_010000011010_000_0_010000011010;
      patterns[8401] = 29'b0_010000011010_001_0_011010010000;
      patterns[8402] = 29'b0_010000011010_010_0_100000110100;
      patterns[8403] = 29'b0_010000011010_011_1_000001101000;
      patterns[8404] = 29'b0_010000011010_100_0_001000001101;
      patterns[8405] = 29'b0_010000011010_101_1_000100000110;
      patterns[8406] = 29'b0_010000011010_110_0_010000011010;
      patterns[8407] = 29'b0_010000011010_111_0_010000011010;
      patterns[8408] = 29'b0_010000011011_000_0_010000011011;
      patterns[8409] = 29'b0_010000011011_001_0_011011010000;
      patterns[8410] = 29'b0_010000011011_010_0_100000110110;
      patterns[8411] = 29'b0_010000011011_011_1_000001101100;
      patterns[8412] = 29'b0_010000011011_100_1_001000001101;
      patterns[8413] = 29'b0_010000011011_101_1_100100000110;
      patterns[8414] = 29'b0_010000011011_110_0_010000011011;
      patterns[8415] = 29'b0_010000011011_111_0_010000011011;
      patterns[8416] = 29'b0_010000011100_000_0_010000011100;
      patterns[8417] = 29'b0_010000011100_001_0_011100010000;
      patterns[8418] = 29'b0_010000011100_010_0_100000111000;
      patterns[8419] = 29'b0_010000011100_011_1_000001110000;
      patterns[8420] = 29'b0_010000011100_100_0_001000001110;
      patterns[8421] = 29'b0_010000011100_101_0_000100000111;
      patterns[8422] = 29'b0_010000011100_110_0_010000011100;
      patterns[8423] = 29'b0_010000011100_111_0_010000011100;
      patterns[8424] = 29'b0_010000011101_000_0_010000011101;
      patterns[8425] = 29'b0_010000011101_001_0_011101010000;
      patterns[8426] = 29'b0_010000011101_010_0_100000111010;
      patterns[8427] = 29'b0_010000011101_011_1_000001110100;
      patterns[8428] = 29'b0_010000011101_100_1_001000001110;
      patterns[8429] = 29'b0_010000011101_101_0_100100000111;
      patterns[8430] = 29'b0_010000011101_110_0_010000011101;
      patterns[8431] = 29'b0_010000011101_111_0_010000011101;
      patterns[8432] = 29'b0_010000011110_000_0_010000011110;
      patterns[8433] = 29'b0_010000011110_001_0_011110010000;
      patterns[8434] = 29'b0_010000011110_010_0_100000111100;
      patterns[8435] = 29'b0_010000011110_011_1_000001111000;
      patterns[8436] = 29'b0_010000011110_100_0_001000001111;
      patterns[8437] = 29'b0_010000011110_101_1_000100000111;
      patterns[8438] = 29'b0_010000011110_110_0_010000011110;
      patterns[8439] = 29'b0_010000011110_111_0_010000011110;
      patterns[8440] = 29'b0_010000011111_000_0_010000011111;
      patterns[8441] = 29'b0_010000011111_001_0_011111010000;
      patterns[8442] = 29'b0_010000011111_010_0_100000111110;
      patterns[8443] = 29'b0_010000011111_011_1_000001111100;
      patterns[8444] = 29'b0_010000011111_100_1_001000001111;
      patterns[8445] = 29'b0_010000011111_101_1_100100000111;
      patterns[8446] = 29'b0_010000011111_110_0_010000011111;
      patterns[8447] = 29'b0_010000011111_111_0_010000011111;
      patterns[8448] = 29'b0_010000100000_000_0_010000100000;
      patterns[8449] = 29'b0_010000100000_001_0_100000010000;
      patterns[8450] = 29'b0_010000100000_010_0_100001000000;
      patterns[8451] = 29'b0_010000100000_011_1_000010000000;
      patterns[8452] = 29'b0_010000100000_100_0_001000010000;
      patterns[8453] = 29'b0_010000100000_101_0_000100001000;
      patterns[8454] = 29'b0_010000100000_110_0_010000100000;
      patterns[8455] = 29'b0_010000100000_111_0_010000100000;
      patterns[8456] = 29'b0_010000100001_000_0_010000100001;
      patterns[8457] = 29'b0_010000100001_001_0_100001010000;
      patterns[8458] = 29'b0_010000100001_010_0_100001000010;
      patterns[8459] = 29'b0_010000100001_011_1_000010000100;
      patterns[8460] = 29'b0_010000100001_100_1_001000010000;
      patterns[8461] = 29'b0_010000100001_101_0_100100001000;
      patterns[8462] = 29'b0_010000100001_110_0_010000100001;
      patterns[8463] = 29'b0_010000100001_111_0_010000100001;
      patterns[8464] = 29'b0_010000100010_000_0_010000100010;
      patterns[8465] = 29'b0_010000100010_001_0_100010010000;
      patterns[8466] = 29'b0_010000100010_010_0_100001000100;
      patterns[8467] = 29'b0_010000100010_011_1_000010001000;
      patterns[8468] = 29'b0_010000100010_100_0_001000010001;
      patterns[8469] = 29'b0_010000100010_101_1_000100001000;
      patterns[8470] = 29'b0_010000100010_110_0_010000100010;
      patterns[8471] = 29'b0_010000100010_111_0_010000100010;
      patterns[8472] = 29'b0_010000100011_000_0_010000100011;
      patterns[8473] = 29'b0_010000100011_001_0_100011010000;
      patterns[8474] = 29'b0_010000100011_010_0_100001000110;
      patterns[8475] = 29'b0_010000100011_011_1_000010001100;
      patterns[8476] = 29'b0_010000100011_100_1_001000010001;
      patterns[8477] = 29'b0_010000100011_101_1_100100001000;
      patterns[8478] = 29'b0_010000100011_110_0_010000100011;
      patterns[8479] = 29'b0_010000100011_111_0_010000100011;
      patterns[8480] = 29'b0_010000100100_000_0_010000100100;
      patterns[8481] = 29'b0_010000100100_001_0_100100010000;
      patterns[8482] = 29'b0_010000100100_010_0_100001001000;
      patterns[8483] = 29'b0_010000100100_011_1_000010010000;
      patterns[8484] = 29'b0_010000100100_100_0_001000010010;
      patterns[8485] = 29'b0_010000100100_101_0_000100001001;
      patterns[8486] = 29'b0_010000100100_110_0_010000100100;
      patterns[8487] = 29'b0_010000100100_111_0_010000100100;
      patterns[8488] = 29'b0_010000100101_000_0_010000100101;
      patterns[8489] = 29'b0_010000100101_001_0_100101010000;
      patterns[8490] = 29'b0_010000100101_010_0_100001001010;
      patterns[8491] = 29'b0_010000100101_011_1_000010010100;
      patterns[8492] = 29'b0_010000100101_100_1_001000010010;
      patterns[8493] = 29'b0_010000100101_101_0_100100001001;
      patterns[8494] = 29'b0_010000100101_110_0_010000100101;
      patterns[8495] = 29'b0_010000100101_111_0_010000100101;
      patterns[8496] = 29'b0_010000100110_000_0_010000100110;
      patterns[8497] = 29'b0_010000100110_001_0_100110010000;
      patterns[8498] = 29'b0_010000100110_010_0_100001001100;
      patterns[8499] = 29'b0_010000100110_011_1_000010011000;
      patterns[8500] = 29'b0_010000100110_100_0_001000010011;
      patterns[8501] = 29'b0_010000100110_101_1_000100001001;
      patterns[8502] = 29'b0_010000100110_110_0_010000100110;
      patterns[8503] = 29'b0_010000100110_111_0_010000100110;
      patterns[8504] = 29'b0_010000100111_000_0_010000100111;
      patterns[8505] = 29'b0_010000100111_001_0_100111010000;
      patterns[8506] = 29'b0_010000100111_010_0_100001001110;
      patterns[8507] = 29'b0_010000100111_011_1_000010011100;
      patterns[8508] = 29'b0_010000100111_100_1_001000010011;
      patterns[8509] = 29'b0_010000100111_101_1_100100001001;
      patterns[8510] = 29'b0_010000100111_110_0_010000100111;
      patterns[8511] = 29'b0_010000100111_111_0_010000100111;
      patterns[8512] = 29'b0_010000101000_000_0_010000101000;
      patterns[8513] = 29'b0_010000101000_001_0_101000010000;
      patterns[8514] = 29'b0_010000101000_010_0_100001010000;
      patterns[8515] = 29'b0_010000101000_011_1_000010100000;
      patterns[8516] = 29'b0_010000101000_100_0_001000010100;
      patterns[8517] = 29'b0_010000101000_101_0_000100001010;
      patterns[8518] = 29'b0_010000101000_110_0_010000101000;
      patterns[8519] = 29'b0_010000101000_111_0_010000101000;
      patterns[8520] = 29'b0_010000101001_000_0_010000101001;
      patterns[8521] = 29'b0_010000101001_001_0_101001010000;
      patterns[8522] = 29'b0_010000101001_010_0_100001010010;
      patterns[8523] = 29'b0_010000101001_011_1_000010100100;
      patterns[8524] = 29'b0_010000101001_100_1_001000010100;
      patterns[8525] = 29'b0_010000101001_101_0_100100001010;
      patterns[8526] = 29'b0_010000101001_110_0_010000101001;
      patterns[8527] = 29'b0_010000101001_111_0_010000101001;
      patterns[8528] = 29'b0_010000101010_000_0_010000101010;
      patterns[8529] = 29'b0_010000101010_001_0_101010010000;
      patterns[8530] = 29'b0_010000101010_010_0_100001010100;
      patterns[8531] = 29'b0_010000101010_011_1_000010101000;
      patterns[8532] = 29'b0_010000101010_100_0_001000010101;
      patterns[8533] = 29'b0_010000101010_101_1_000100001010;
      patterns[8534] = 29'b0_010000101010_110_0_010000101010;
      patterns[8535] = 29'b0_010000101010_111_0_010000101010;
      patterns[8536] = 29'b0_010000101011_000_0_010000101011;
      patterns[8537] = 29'b0_010000101011_001_0_101011010000;
      patterns[8538] = 29'b0_010000101011_010_0_100001010110;
      patterns[8539] = 29'b0_010000101011_011_1_000010101100;
      patterns[8540] = 29'b0_010000101011_100_1_001000010101;
      patterns[8541] = 29'b0_010000101011_101_1_100100001010;
      patterns[8542] = 29'b0_010000101011_110_0_010000101011;
      patterns[8543] = 29'b0_010000101011_111_0_010000101011;
      patterns[8544] = 29'b0_010000101100_000_0_010000101100;
      patterns[8545] = 29'b0_010000101100_001_0_101100010000;
      patterns[8546] = 29'b0_010000101100_010_0_100001011000;
      patterns[8547] = 29'b0_010000101100_011_1_000010110000;
      patterns[8548] = 29'b0_010000101100_100_0_001000010110;
      patterns[8549] = 29'b0_010000101100_101_0_000100001011;
      patterns[8550] = 29'b0_010000101100_110_0_010000101100;
      patterns[8551] = 29'b0_010000101100_111_0_010000101100;
      patterns[8552] = 29'b0_010000101101_000_0_010000101101;
      patterns[8553] = 29'b0_010000101101_001_0_101101010000;
      patterns[8554] = 29'b0_010000101101_010_0_100001011010;
      patterns[8555] = 29'b0_010000101101_011_1_000010110100;
      patterns[8556] = 29'b0_010000101101_100_1_001000010110;
      patterns[8557] = 29'b0_010000101101_101_0_100100001011;
      patterns[8558] = 29'b0_010000101101_110_0_010000101101;
      patterns[8559] = 29'b0_010000101101_111_0_010000101101;
      patterns[8560] = 29'b0_010000101110_000_0_010000101110;
      patterns[8561] = 29'b0_010000101110_001_0_101110010000;
      patterns[8562] = 29'b0_010000101110_010_0_100001011100;
      patterns[8563] = 29'b0_010000101110_011_1_000010111000;
      patterns[8564] = 29'b0_010000101110_100_0_001000010111;
      patterns[8565] = 29'b0_010000101110_101_1_000100001011;
      patterns[8566] = 29'b0_010000101110_110_0_010000101110;
      patterns[8567] = 29'b0_010000101110_111_0_010000101110;
      patterns[8568] = 29'b0_010000101111_000_0_010000101111;
      patterns[8569] = 29'b0_010000101111_001_0_101111010000;
      patterns[8570] = 29'b0_010000101111_010_0_100001011110;
      patterns[8571] = 29'b0_010000101111_011_1_000010111100;
      patterns[8572] = 29'b0_010000101111_100_1_001000010111;
      patterns[8573] = 29'b0_010000101111_101_1_100100001011;
      patterns[8574] = 29'b0_010000101111_110_0_010000101111;
      patterns[8575] = 29'b0_010000101111_111_0_010000101111;
      patterns[8576] = 29'b0_010000110000_000_0_010000110000;
      patterns[8577] = 29'b0_010000110000_001_0_110000010000;
      patterns[8578] = 29'b0_010000110000_010_0_100001100000;
      patterns[8579] = 29'b0_010000110000_011_1_000011000000;
      patterns[8580] = 29'b0_010000110000_100_0_001000011000;
      patterns[8581] = 29'b0_010000110000_101_0_000100001100;
      patterns[8582] = 29'b0_010000110000_110_0_010000110000;
      patterns[8583] = 29'b0_010000110000_111_0_010000110000;
      patterns[8584] = 29'b0_010000110001_000_0_010000110001;
      patterns[8585] = 29'b0_010000110001_001_0_110001010000;
      patterns[8586] = 29'b0_010000110001_010_0_100001100010;
      patterns[8587] = 29'b0_010000110001_011_1_000011000100;
      patterns[8588] = 29'b0_010000110001_100_1_001000011000;
      patterns[8589] = 29'b0_010000110001_101_0_100100001100;
      patterns[8590] = 29'b0_010000110001_110_0_010000110001;
      patterns[8591] = 29'b0_010000110001_111_0_010000110001;
      patterns[8592] = 29'b0_010000110010_000_0_010000110010;
      patterns[8593] = 29'b0_010000110010_001_0_110010010000;
      patterns[8594] = 29'b0_010000110010_010_0_100001100100;
      patterns[8595] = 29'b0_010000110010_011_1_000011001000;
      patterns[8596] = 29'b0_010000110010_100_0_001000011001;
      patterns[8597] = 29'b0_010000110010_101_1_000100001100;
      patterns[8598] = 29'b0_010000110010_110_0_010000110010;
      patterns[8599] = 29'b0_010000110010_111_0_010000110010;
      patterns[8600] = 29'b0_010000110011_000_0_010000110011;
      patterns[8601] = 29'b0_010000110011_001_0_110011010000;
      patterns[8602] = 29'b0_010000110011_010_0_100001100110;
      patterns[8603] = 29'b0_010000110011_011_1_000011001100;
      patterns[8604] = 29'b0_010000110011_100_1_001000011001;
      patterns[8605] = 29'b0_010000110011_101_1_100100001100;
      patterns[8606] = 29'b0_010000110011_110_0_010000110011;
      patterns[8607] = 29'b0_010000110011_111_0_010000110011;
      patterns[8608] = 29'b0_010000110100_000_0_010000110100;
      patterns[8609] = 29'b0_010000110100_001_0_110100010000;
      patterns[8610] = 29'b0_010000110100_010_0_100001101000;
      patterns[8611] = 29'b0_010000110100_011_1_000011010000;
      patterns[8612] = 29'b0_010000110100_100_0_001000011010;
      patterns[8613] = 29'b0_010000110100_101_0_000100001101;
      patterns[8614] = 29'b0_010000110100_110_0_010000110100;
      patterns[8615] = 29'b0_010000110100_111_0_010000110100;
      patterns[8616] = 29'b0_010000110101_000_0_010000110101;
      patterns[8617] = 29'b0_010000110101_001_0_110101010000;
      patterns[8618] = 29'b0_010000110101_010_0_100001101010;
      patterns[8619] = 29'b0_010000110101_011_1_000011010100;
      patterns[8620] = 29'b0_010000110101_100_1_001000011010;
      patterns[8621] = 29'b0_010000110101_101_0_100100001101;
      patterns[8622] = 29'b0_010000110101_110_0_010000110101;
      patterns[8623] = 29'b0_010000110101_111_0_010000110101;
      patterns[8624] = 29'b0_010000110110_000_0_010000110110;
      patterns[8625] = 29'b0_010000110110_001_0_110110010000;
      patterns[8626] = 29'b0_010000110110_010_0_100001101100;
      patterns[8627] = 29'b0_010000110110_011_1_000011011000;
      patterns[8628] = 29'b0_010000110110_100_0_001000011011;
      patterns[8629] = 29'b0_010000110110_101_1_000100001101;
      patterns[8630] = 29'b0_010000110110_110_0_010000110110;
      patterns[8631] = 29'b0_010000110110_111_0_010000110110;
      patterns[8632] = 29'b0_010000110111_000_0_010000110111;
      patterns[8633] = 29'b0_010000110111_001_0_110111010000;
      patterns[8634] = 29'b0_010000110111_010_0_100001101110;
      patterns[8635] = 29'b0_010000110111_011_1_000011011100;
      patterns[8636] = 29'b0_010000110111_100_1_001000011011;
      patterns[8637] = 29'b0_010000110111_101_1_100100001101;
      patterns[8638] = 29'b0_010000110111_110_0_010000110111;
      patterns[8639] = 29'b0_010000110111_111_0_010000110111;
      patterns[8640] = 29'b0_010000111000_000_0_010000111000;
      patterns[8641] = 29'b0_010000111000_001_0_111000010000;
      patterns[8642] = 29'b0_010000111000_010_0_100001110000;
      patterns[8643] = 29'b0_010000111000_011_1_000011100000;
      patterns[8644] = 29'b0_010000111000_100_0_001000011100;
      patterns[8645] = 29'b0_010000111000_101_0_000100001110;
      patterns[8646] = 29'b0_010000111000_110_0_010000111000;
      patterns[8647] = 29'b0_010000111000_111_0_010000111000;
      patterns[8648] = 29'b0_010000111001_000_0_010000111001;
      patterns[8649] = 29'b0_010000111001_001_0_111001010000;
      patterns[8650] = 29'b0_010000111001_010_0_100001110010;
      patterns[8651] = 29'b0_010000111001_011_1_000011100100;
      patterns[8652] = 29'b0_010000111001_100_1_001000011100;
      patterns[8653] = 29'b0_010000111001_101_0_100100001110;
      patterns[8654] = 29'b0_010000111001_110_0_010000111001;
      patterns[8655] = 29'b0_010000111001_111_0_010000111001;
      patterns[8656] = 29'b0_010000111010_000_0_010000111010;
      patterns[8657] = 29'b0_010000111010_001_0_111010010000;
      patterns[8658] = 29'b0_010000111010_010_0_100001110100;
      patterns[8659] = 29'b0_010000111010_011_1_000011101000;
      patterns[8660] = 29'b0_010000111010_100_0_001000011101;
      patterns[8661] = 29'b0_010000111010_101_1_000100001110;
      patterns[8662] = 29'b0_010000111010_110_0_010000111010;
      patterns[8663] = 29'b0_010000111010_111_0_010000111010;
      patterns[8664] = 29'b0_010000111011_000_0_010000111011;
      patterns[8665] = 29'b0_010000111011_001_0_111011010000;
      patterns[8666] = 29'b0_010000111011_010_0_100001110110;
      patterns[8667] = 29'b0_010000111011_011_1_000011101100;
      patterns[8668] = 29'b0_010000111011_100_1_001000011101;
      patterns[8669] = 29'b0_010000111011_101_1_100100001110;
      patterns[8670] = 29'b0_010000111011_110_0_010000111011;
      patterns[8671] = 29'b0_010000111011_111_0_010000111011;
      patterns[8672] = 29'b0_010000111100_000_0_010000111100;
      patterns[8673] = 29'b0_010000111100_001_0_111100010000;
      patterns[8674] = 29'b0_010000111100_010_0_100001111000;
      patterns[8675] = 29'b0_010000111100_011_1_000011110000;
      patterns[8676] = 29'b0_010000111100_100_0_001000011110;
      patterns[8677] = 29'b0_010000111100_101_0_000100001111;
      patterns[8678] = 29'b0_010000111100_110_0_010000111100;
      patterns[8679] = 29'b0_010000111100_111_0_010000111100;
      patterns[8680] = 29'b0_010000111101_000_0_010000111101;
      patterns[8681] = 29'b0_010000111101_001_0_111101010000;
      patterns[8682] = 29'b0_010000111101_010_0_100001111010;
      patterns[8683] = 29'b0_010000111101_011_1_000011110100;
      patterns[8684] = 29'b0_010000111101_100_1_001000011110;
      patterns[8685] = 29'b0_010000111101_101_0_100100001111;
      patterns[8686] = 29'b0_010000111101_110_0_010000111101;
      patterns[8687] = 29'b0_010000111101_111_0_010000111101;
      patterns[8688] = 29'b0_010000111110_000_0_010000111110;
      patterns[8689] = 29'b0_010000111110_001_0_111110010000;
      patterns[8690] = 29'b0_010000111110_010_0_100001111100;
      patterns[8691] = 29'b0_010000111110_011_1_000011111000;
      patterns[8692] = 29'b0_010000111110_100_0_001000011111;
      patterns[8693] = 29'b0_010000111110_101_1_000100001111;
      patterns[8694] = 29'b0_010000111110_110_0_010000111110;
      patterns[8695] = 29'b0_010000111110_111_0_010000111110;
      patterns[8696] = 29'b0_010000111111_000_0_010000111111;
      patterns[8697] = 29'b0_010000111111_001_0_111111010000;
      patterns[8698] = 29'b0_010000111111_010_0_100001111110;
      patterns[8699] = 29'b0_010000111111_011_1_000011111100;
      patterns[8700] = 29'b0_010000111111_100_1_001000011111;
      patterns[8701] = 29'b0_010000111111_101_1_100100001111;
      patterns[8702] = 29'b0_010000111111_110_0_010000111111;
      patterns[8703] = 29'b0_010000111111_111_0_010000111111;
      patterns[8704] = 29'b0_010001000000_000_0_010001000000;
      patterns[8705] = 29'b0_010001000000_001_0_000000010001;
      patterns[8706] = 29'b0_010001000000_010_0_100010000000;
      patterns[8707] = 29'b0_010001000000_011_1_000100000000;
      patterns[8708] = 29'b0_010001000000_100_0_001000100000;
      patterns[8709] = 29'b0_010001000000_101_0_000100010000;
      patterns[8710] = 29'b0_010001000000_110_0_010001000000;
      patterns[8711] = 29'b0_010001000000_111_0_010001000000;
      patterns[8712] = 29'b0_010001000001_000_0_010001000001;
      patterns[8713] = 29'b0_010001000001_001_0_000001010001;
      patterns[8714] = 29'b0_010001000001_010_0_100010000010;
      patterns[8715] = 29'b0_010001000001_011_1_000100000100;
      patterns[8716] = 29'b0_010001000001_100_1_001000100000;
      patterns[8717] = 29'b0_010001000001_101_0_100100010000;
      patterns[8718] = 29'b0_010001000001_110_0_010001000001;
      patterns[8719] = 29'b0_010001000001_111_0_010001000001;
      patterns[8720] = 29'b0_010001000010_000_0_010001000010;
      patterns[8721] = 29'b0_010001000010_001_0_000010010001;
      patterns[8722] = 29'b0_010001000010_010_0_100010000100;
      patterns[8723] = 29'b0_010001000010_011_1_000100001000;
      patterns[8724] = 29'b0_010001000010_100_0_001000100001;
      patterns[8725] = 29'b0_010001000010_101_1_000100010000;
      patterns[8726] = 29'b0_010001000010_110_0_010001000010;
      patterns[8727] = 29'b0_010001000010_111_0_010001000010;
      patterns[8728] = 29'b0_010001000011_000_0_010001000011;
      patterns[8729] = 29'b0_010001000011_001_0_000011010001;
      patterns[8730] = 29'b0_010001000011_010_0_100010000110;
      patterns[8731] = 29'b0_010001000011_011_1_000100001100;
      patterns[8732] = 29'b0_010001000011_100_1_001000100001;
      patterns[8733] = 29'b0_010001000011_101_1_100100010000;
      patterns[8734] = 29'b0_010001000011_110_0_010001000011;
      patterns[8735] = 29'b0_010001000011_111_0_010001000011;
      patterns[8736] = 29'b0_010001000100_000_0_010001000100;
      patterns[8737] = 29'b0_010001000100_001_0_000100010001;
      patterns[8738] = 29'b0_010001000100_010_0_100010001000;
      patterns[8739] = 29'b0_010001000100_011_1_000100010000;
      patterns[8740] = 29'b0_010001000100_100_0_001000100010;
      patterns[8741] = 29'b0_010001000100_101_0_000100010001;
      patterns[8742] = 29'b0_010001000100_110_0_010001000100;
      patterns[8743] = 29'b0_010001000100_111_0_010001000100;
      patterns[8744] = 29'b0_010001000101_000_0_010001000101;
      patterns[8745] = 29'b0_010001000101_001_0_000101010001;
      patterns[8746] = 29'b0_010001000101_010_0_100010001010;
      patterns[8747] = 29'b0_010001000101_011_1_000100010100;
      patterns[8748] = 29'b0_010001000101_100_1_001000100010;
      patterns[8749] = 29'b0_010001000101_101_0_100100010001;
      patterns[8750] = 29'b0_010001000101_110_0_010001000101;
      patterns[8751] = 29'b0_010001000101_111_0_010001000101;
      patterns[8752] = 29'b0_010001000110_000_0_010001000110;
      patterns[8753] = 29'b0_010001000110_001_0_000110010001;
      patterns[8754] = 29'b0_010001000110_010_0_100010001100;
      patterns[8755] = 29'b0_010001000110_011_1_000100011000;
      patterns[8756] = 29'b0_010001000110_100_0_001000100011;
      patterns[8757] = 29'b0_010001000110_101_1_000100010001;
      patterns[8758] = 29'b0_010001000110_110_0_010001000110;
      patterns[8759] = 29'b0_010001000110_111_0_010001000110;
      patterns[8760] = 29'b0_010001000111_000_0_010001000111;
      patterns[8761] = 29'b0_010001000111_001_0_000111010001;
      patterns[8762] = 29'b0_010001000111_010_0_100010001110;
      patterns[8763] = 29'b0_010001000111_011_1_000100011100;
      patterns[8764] = 29'b0_010001000111_100_1_001000100011;
      patterns[8765] = 29'b0_010001000111_101_1_100100010001;
      patterns[8766] = 29'b0_010001000111_110_0_010001000111;
      patterns[8767] = 29'b0_010001000111_111_0_010001000111;
      patterns[8768] = 29'b0_010001001000_000_0_010001001000;
      patterns[8769] = 29'b0_010001001000_001_0_001000010001;
      patterns[8770] = 29'b0_010001001000_010_0_100010010000;
      patterns[8771] = 29'b0_010001001000_011_1_000100100000;
      patterns[8772] = 29'b0_010001001000_100_0_001000100100;
      patterns[8773] = 29'b0_010001001000_101_0_000100010010;
      patterns[8774] = 29'b0_010001001000_110_0_010001001000;
      patterns[8775] = 29'b0_010001001000_111_0_010001001000;
      patterns[8776] = 29'b0_010001001001_000_0_010001001001;
      patterns[8777] = 29'b0_010001001001_001_0_001001010001;
      patterns[8778] = 29'b0_010001001001_010_0_100010010010;
      patterns[8779] = 29'b0_010001001001_011_1_000100100100;
      patterns[8780] = 29'b0_010001001001_100_1_001000100100;
      patterns[8781] = 29'b0_010001001001_101_0_100100010010;
      patterns[8782] = 29'b0_010001001001_110_0_010001001001;
      patterns[8783] = 29'b0_010001001001_111_0_010001001001;
      patterns[8784] = 29'b0_010001001010_000_0_010001001010;
      patterns[8785] = 29'b0_010001001010_001_0_001010010001;
      patterns[8786] = 29'b0_010001001010_010_0_100010010100;
      patterns[8787] = 29'b0_010001001010_011_1_000100101000;
      patterns[8788] = 29'b0_010001001010_100_0_001000100101;
      patterns[8789] = 29'b0_010001001010_101_1_000100010010;
      patterns[8790] = 29'b0_010001001010_110_0_010001001010;
      patterns[8791] = 29'b0_010001001010_111_0_010001001010;
      patterns[8792] = 29'b0_010001001011_000_0_010001001011;
      patterns[8793] = 29'b0_010001001011_001_0_001011010001;
      patterns[8794] = 29'b0_010001001011_010_0_100010010110;
      patterns[8795] = 29'b0_010001001011_011_1_000100101100;
      patterns[8796] = 29'b0_010001001011_100_1_001000100101;
      patterns[8797] = 29'b0_010001001011_101_1_100100010010;
      patterns[8798] = 29'b0_010001001011_110_0_010001001011;
      patterns[8799] = 29'b0_010001001011_111_0_010001001011;
      patterns[8800] = 29'b0_010001001100_000_0_010001001100;
      patterns[8801] = 29'b0_010001001100_001_0_001100010001;
      patterns[8802] = 29'b0_010001001100_010_0_100010011000;
      patterns[8803] = 29'b0_010001001100_011_1_000100110000;
      patterns[8804] = 29'b0_010001001100_100_0_001000100110;
      patterns[8805] = 29'b0_010001001100_101_0_000100010011;
      patterns[8806] = 29'b0_010001001100_110_0_010001001100;
      patterns[8807] = 29'b0_010001001100_111_0_010001001100;
      patterns[8808] = 29'b0_010001001101_000_0_010001001101;
      patterns[8809] = 29'b0_010001001101_001_0_001101010001;
      patterns[8810] = 29'b0_010001001101_010_0_100010011010;
      patterns[8811] = 29'b0_010001001101_011_1_000100110100;
      patterns[8812] = 29'b0_010001001101_100_1_001000100110;
      patterns[8813] = 29'b0_010001001101_101_0_100100010011;
      patterns[8814] = 29'b0_010001001101_110_0_010001001101;
      patterns[8815] = 29'b0_010001001101_111_0_010001001101;
      patterns[8816] = 29'b0_010001001110_000_0_010001001110;
      patterns[8817] = 29'b0_010001001110_001_0_001110010001;
      patterns[8818] = 29'b0_010001001110_010_0_100010011100;
      patterns[8819] = 29'b0_010001001110_011_1_000100111000;
      patterns[8820] = 29'b0_010001001110_100_0_001000100111;
      patterns[8821] = 29'b0_010001001110_101_1_000100010011;
      patterns[8822] = 29'b0_010001001110_110_0_010001001110;
      patterns[8823] = 29'b0_010001001110_111_0_010001001110;
      patterns[8824] = 29'b0_010001001111_000_0_010001001111;
      patterns[8825] = 29'b0_010001001111_001_0_001111010001;
      patterns[8826] = 29'b0_010001001111_010_0_100010011110;
      patterns[8827] = 29'b0_010001001111_011_1_000100111100;
      patterns[8828] = 29'b0_010001001111_100_1_001000100111;
      patterns[8829] = 29'b0_010001001111_101_1_100100010011;
      patterns[8830] = 29'b0_010001001111_110_0_010001001111;
      patterns[8831] = 29'b0_010001001111_111_0_010001001111;
      patterns[8832] = 29'b0_010001010000_000_0_010001010000;
      patterns[8833] = 29'b0_010001010000_001_0_010000010001;
      patterns[8834] = 29'b0_010001010000_010_0_100010100000;
      patterns[8835] = 29'b0_010001010000_011_1_000101000000;
      patterns[8836] = 29'b0_010001010000_100_0_001000101000;
      patterns[8837] = 29'b0_010001010000_101_0_000100010100;
      patterns[8838] = 29'b0_010001010000_110_0_010001010000;
      patterns[8839] = 29'b0_010001010000_111_0_010001010000;
      patterns[8840] = 29'b0_010001010001_000_0_010001010001;
      patterns[8841] = 29'b0_010001010001_001_0_010001010001;
      patterns[8842] = 29'b0_010001010001_010_0_100010100010;
      patterns[8843] = 29'b0_010001010001_011_1_000101000100;
      patterns[8844] = 29'b0_010001010001_100_1_001000101000;
      patterns[8845] = 29'b0_010001010001_101_0_100100010100;
      patterns[8846] = 29'b0_010001010001_110_0_010001010001;
      patterns[8847] = 29'b0_010001010001_111_0_010001010001;
      patterns[8848] = 29'b0_010001010010_000_0_010001010010;
      patterns[8849] = 29'b0_010001010010_001_0_010010010001;
      patterns[8850] = 29'b0_010001010010_010_0_100010100100;
      patterns[8851] = 29'b0_010001010010_011_1_000101001000;
      patterns[8852] = 29'b0_010001010010_100_0_001000101001;
      patterns[8853] = 29'b0_010001010010_101_1_000100010100;
      patterns[8854] = 29'b0_010001010010_110_0_010001010010;
      patterns[8855] = 29'b0_010001010010_111_0_010001010010;
      patterns[8856] = 29'b0_010001010011_000_0_010001010011;
      patterns[8857] = 29'b0_010001010011_001_0_010011010001;
      patterns[8858] = 29'b0_010001010011_010_0_100010100110;
      patterns[8859] = 29'b0_010001010011_011_1_000101001100;
      patterns[8860] = 29'b0_010001010011_100_1_001000101001;
      patterns[8861] = 29'b0_010001010011_101_1_100100010100;
      patterns[8862] = 29'b0_010001010011_110_0_010001010011;
      patterns[8863] = 29'b0_010001010011_111_0_010001010011;
      patterns[8864] = 29'b0_010001010100_000_0_010001010100;
      patterns[8865] = 29'b0_010001010100_001_0_010100010001;
      patterns[8866] = 29'b0_010001010100_010_0_100010101000;
      patterns[8867] = 29'b0_010001010100_011_1_000101010000;
      patterns[8868] = 29'b0_010001010100_100_0_001000101010;
      patterns[8869] = 29'b0_010001010100_101_0_000100010101;
      patterns[8870] = 29'b0_010001010100_110_0_010001010100;
      patterns[8871] = 29'b0_010001010100_111_0_010001010100;
      patterns[8872] = 29'b0_010001010101_000_0_010001010101;
      patterns[8873] = 29'b0_010001010101_001_0_010101010001;
      patterns[8874] = 29'b0_010001010101_010_0_100010101010;
      patterns[8875] = 29'b0_010001010101_011_1_000101010100;
      patterns[8876] = 29'b0_010001010101_100_1_001000101010;
      patterns[8877] = 29'b0_010001010101_101_0_100100010101;
      patterns[8878] = 29'b0_010001010101_110_0_010001010101;
      patterns[8879] = 29'b0_010001010101_111_0_010001010101;
      patterns[8880] = 29'b0_010001010110_000_0_010001010110;
      patterns[8881] = 29'b0_010001010110_001_0_010110010001;
      patterns[8882] = 29'b0_010001010110_010_0_100010101100;
      patterns[8883] = 29'b0_010001010110_011_1_000101011000;
      patterns[8884] = 29'b0_010001010110_100_0_001000101011;
      patterns[8885] = 29'b0_010001010110_101_1_000100010101;
      patterns[8886] = 29'b0_010001010110_110_0_010001010110;
      patterns[8887] = 29'b0_010001010110_111_0_010001010110;
      patterns[8888] = 29'b0_010001010111_000_0_010001010111;
      patterns[8889] = 29'b0_010001010111_001_0_010111010001;
      patterns[8890] = 29'b0_010001010111_010_0_100010101110;
      patterns[8891] = 29'b0_010001010111_011_1_000101011100;
      patterns[8892] = 29'b0_010001010111_100_1_001000101011;
      patterns[8893] = 29'b0_010001010111_101_1_100100010101;
      patterns[8894] = 29'b0_010001010111_110_0_010001010111;
      patterns[8895] = 29'b0_010001010111_111_0_010001010111;
      patterns[8896] = 29'b0_010001011000_000_0_010001011000;
      patterns[8897] = 29'b0_010001011000_001_0_011000010001;
      patterns[8898] = 29'b0_010001011000_010_0_100010110000;
      patterns[8899] = 29'b0_010001011000_011_1_000101100000;
      patterns[8900] = 29'b0_010001011000_100_0_001000101100;
      patterns[8901] = 29'b0_010001011000_101_0_000100010110;
      patterns[8902] = 29'b0_010001011000_110_0_010001011000;
      patterns[8903] = 29'b0_010001011000_111_0_010001011000;
      patterns[8904] = 29'b0_010001011001_000_0_010001011001;
      patterns[8905] = 29'b0_010001011001_001_0_011001010001;
      patterns[8906] = 29'b0_010001011001_010_0_100010110010;
      patterns[8907] = 29'b0_010001011001_011_1_000101100100;
      patterns[8908] = 29'b0_010001011001_100_1_001000101100;
      patterns[8909] = 29'b0_010001011001_101_0_100100010110;
      patterns[8910] = 29'b0_010001011001_110_0_010001011001;
      patterns[8911] = 29'b0_010001011001_111_0_010001011001;
      patterns[8912] = 29'b0_010001011010_000_0_010001011010;
      patterns[8913] = 29'b0_010001011010_001_0_011010010001;
      patterns[8914] = 29'b0_010001011010_010_0_100010110100;
      patterns[8915] = 29'b0_010001011010_011_1_000101101000;
      patterns[8916] = 29'b0_010001011010_100_0_001000101101;
      patterns[8917] = 29'b0_010001011010_101_1_000100010110;
      patterns[8918] = 29'b0_010001011010_110_0_010001011010;
      patterns[8919] = 29'b0_010001011010_111_0_010001011010;
      patterns[8920] = 29'b0_010001011011_000_0_010001011011;
      patterns[8921] = 29'b0_010001011011_001_0_011011010001;
      patterns[8922] = 29'b0_010001011011_010_0_100010110110;
      patterns[8923] = 29'b0_010001011011_011_1_000101101100;
      patterns[8924] = 29'b0_010001011011_100_1_001000101101;
      patterns[8925] = 29'b0_010001011011_101_1_100100010110;
      patterns[8926] = 29'b0_010001011011_110_0_010001011011;
      patterns[8927] = 29'b0_010001011011_111_0_010001011011;
      patterns[8928] = 29'b0_010001011100_000_0_010001011100;
      patterns[8929] = 29'b0_010001011100_001_0_011100010001;
      patterns[8930] = 29'b0_010001011100_010_0_100010111000;
      patterns[8931] = 29'b0_010001011100_011_1_000101110000;
      patterns[8932] = 29'b0_010001011100_100_0_001000101110;
      patterns[8933] = 29'b0_010001011100_101_0_000100010111;
      patterns[8934] = 29'b0_010001011100_110_0_010001011100;
      patterns[8935] = 29'b0_010001011100_111_0_010001011100;
      patterns[8936] = 29'b0_010001011101_000_0_010001011101;
      patterns[8937] = 29'b0_010001011101_001_0_011101010001;
      patterns[8938] = 29'b0_010001011101_010_0_100010111010;
      patterns[8939] = 29'b0_010001011101_011_1_000101110100;
      patterns[8940] = 29'b0_010001011101_100_1_001000101110;
      patterns[8941] = 29'b0_010001011101_101_0_100100010111;
      patterns[8942] = 29'b0_010001011101_110_0_010001011101;
      patterns[8943] = 29'b0_010001011101_111_0_010001011101;
      patterns[8944] = 29'b0_010001011110_000_0_010001011110;
      patterns[8945] = 29'b0_010001011110_001_0_011110010001;
      patterns[8946] = 29'b0_010001011110_010_0_100010111100;
      patterns[8947] = 29'b0_010001011110_011_1_000101111000;
      patterns[8948] = 29'b0_010001011110_100_0_001000101111;
      patterns[8949] = 29'b0_010001011110_101_1_000100010111;
      patterns[8950] = 29'b0_010001011110_110_0_010001011110;
      patterns[8951] = 29'b0_010001011110_111_0_010001011110;
      patterns[8952] = 29'b0_010001011111_000_0_010001011111;
      patterns[8953] = 29'b0_010001011111_001_0_011111010001;
      patterns[8954] = 29'b0_010001011111_010_0_100010111110;
      patterns[8955] = 29'b0_010001011111_011_1_000101111100;
      patterns[8956] = 29'b0_010001011111_100_1_001000101111;
      patterns[8957] = 29'b0_010001011111_101_1_100100010111;
      patterns[8958] = 29'b0_010001011111_110_0_010001011111;
      patterns[8959] = 29'b0_010001011111_111_0_010001011111;
      patterns[8960] = 29'b0_010001100000_000_0_010001100000;
      patterns[8961] = 29'b0_010001100000_001_0_100000010001;
      patterns[8962] = 29'b0_010001100000_010_0_100011000000;
      patterns[8963] = 29'b0_010001100000_011_1_000110000000;
      patterns[8964] = 29'b0_010001100000_100_0_001000110000;
      patterns[8965] = 29'b0_010001100000_101_0_000100011000;
      patterns[8966] = 29'b0_010001100000_110_0_010001100000;
      patterns[8967] = 29'b0_010001100000_111_0_010001100000;
      patterns[8968] = 29'b0_010001100001_000_0_010001100001;
      patterns[8969] = 29'b0_010001100001_001_0_100001010001;
      patterns[8970] = 29'b0_010001100001_010_0_100011000010;
      patterns[8971] = 29'b0_010001100001_011_1_000110000100;
      patterns[8972] = 29'b0_010001100001_100_1_001000110000;
      patterns[8973] = 29'b0_010001100001_101_0_100100011000;
      patterns[8974] = 29'b0_010001100001_110_0_010001100001;
      patterns[8975] = 29'b0_010001100001_111_0_010001100001;
      patterns[8976] = 29'b0_010001100010_000_0_010001100010;
      patterns[8977] = 29'b0_010001100010_001_0_100010010001;
      patterns[8978] = 29'b0_010001100010_010_0_100011000100;
      patterns[8979] = 29'b0_010001100010_011_1_000110001000;
      patterns[8980] = 29'b0_010001100010_100_0_001000110001;
      patterns[8981] = 29'b0_010001100010_101_1_000100011000;
      patterns[8982] = 29'b0_010001100010_110_0_010001100010;
      patterns[8983] = 29'b0_010001100010_111_0_010001100010;
      patterns[8984] = 29'b0_010001100011_000_0_010001100011;
      patterns[8985] = 29'b0_010001100011_001_0_100011010001;
      patterns[8986] = 29'b0_010001100011_010_0_100011000110;
      patterns[8987] = 29'b0_010001100011_011_1_000110001100;
      patterns[8988] = 29'b0_010001100011_100_1_001000110001;
      patterns[8989] = 29'b0_010001100011_101_1_100100011000;
      patterns[8990] = 29'b0_010001100011_110_0_010001100011;
      patterns[8991] = 29'b0_010001100011_111_0_010001100011;
      patterns[8992] = 29'b0_010001100100_000_0_010001100100;
      patterns[8993] = 29'b0_010001100100_001_0_100100010001;
      patterns[8994] = 29'b0_010001100100_010_0_100011001000;
      patterns[8995] = 29'b0_010001100100_011_1_000110010000;
      patterns[8996] = 29'b0_010001100100_100_0_001000110010;
      patterns[8997] = 29'b0_010001100100_101_0_000100011001;
      patterns[8998] = 29'b0_010001100100_110_0_010001100100;
      patterns[8999] = 29'b0_010001100100_111_0_010001100100;
      patterns[9000] = 29'b0_010001100101_000_0_010001100101;
      patterns[9001] = 29'b0_010001100101_001_0_100101010001;
      patterns[9002] = 29'b0_010001100101_010_0_100011001010;
      patterns[9003] = 29'b0_010001100101_011_1_000110010100;
      patterns[9004] = 29'b0_010001100101_100_1_001000110010;
      patterns[9005] = 29'b0_010001100101_101_0_100100011001;
      patterns[9006] = 29'b0_010001100101_110_0_010001100101;
      patterns[9007] = 29'b0_010001100101_111_0_010001100101;
      patterns[9008] = 29'b0_010001100110_000_0_010001100110;
      patterns[9009] = 29'b0_010001100110_001_0_100110010001;
      patterns[9010] = 29'b0_010001100110_010_0_100011001100;
      patterns[9011] = 29'b0_010001100110_011_1_000110011000;
      patterns[9012] = 29'b0_010001100110_100_0_001000110011;
      patterns[9013] = 29'b0_010001100110_101_1_000100011001;
      patterns[9014] = 29'b0_010001100110_110_0_010001100110;
      patterns[9015] = 29'b0_010001100110_111_0_010001100110;
      patterns[9016] = 29'b0_010001100111_000_0_010001100111;
      patterns[9017] = 29'b0_010001100111_001_0_100111010001;
      patterns[9018] = 29'b0_010001100111_010_0_100011001110;
      patterns[9019] = 29'b0_010001100111_011_1_000110011100;
      patterns[9020] = 29'b0_010001100111_100_1_001000110011;
      patterns[9021] = 29'b0_010001100111_101_1_100100011001;
      patterns[9022] = 29'b0_010001100111_110_0_010001100111;
      patterns[9023] = 29'b0_010001100111_111_0_010001100111;
      patterns[9024] = 29'b0_010001101000_000_0_010001101000;
      patterns[9025] = 29'b0_010001101000_001_0_101000010001;
      patterns[9026] = 29'b0_010001101000_010_0_100011010000;
      patterns[9027] = 29'b0_010001101000_011_1_000110100000;
      patterns[9028] = 29'b0_010001101000_100_0_001000110100;
      patterns[9029] = 29'b0_010001101000_101_0_000100011010;
      patterns[9030] = 29'b0_010001101000_110_0_010001101000;
      patterns[9031] = 29'b0_010001101000_111_0_010001101000;
      patterns[9032] = 29'b0_010001101001_000_0_010001101001;
      patterns[9033] = 29'b0_010001101001_001_0_101001010001;
      patterns[9034] = 29'b0_010001101001_010_0_100011010010;
      patterns[9035] = 29'b0_010001101001_011_1_000110100100;
      patterns[9036] = 29'b0_010001101001_100_1_001000110100;
      patterns[9037] = 29'b0_010001101001_101_0_100100011010;
      patterns[9038] = 29'b0_010001101001_110_0_010001101001;
      patterns[9039] = 29'b0_010001101001_111_0_010001101001;
      patterns[9040] = 29'b0_010001101010_000_0_010001101010;
      patterns[9041] = 29'b0_010001101010_001_0_101010010001;
      patterns[9042] = 29'b0_010001101010_010_0_100011010100;
      patterns[9043] = 29'b0_010001101010_011_1_000110101000;
      patterns[9044] = 29'b0_010001101010_100_0_001000110101;
      patterns[9045] = 29'b0_010001101010_101_1_000100011010;
      patterns[9046] = 29'b0_010001101010_110_0_010001101010;
      patterns[9047] = 29'b0_010001101010_111_0_010001101010;
      patterns[9048] = 29'b0_010001101011_000_0_010001101011;
      patterns[9049] = 29'b0_010001101011_001_0_101011010001;
      patterns[9050] = 29'b0_010001101011_010_0_100011010110;
      patterns[9051] = 29'b0_010001101011_011_1_000110101100;
      patterns[9052] = 29'b0_010001101011_100_1_001000110101;
      patterns[9053] = 29'b0_010001101011_101_1_100100011010;
      patterns[9054] = 29'b0_010001101011_110_0_010001101011;
      patterns[9055] = 29'b0_010001101011_111_0_010001101011;
      patterns[9056] = 29'b0_010001101100_000_0_010001101100;
      patterns[9057] = 29'b0_010001101100_001_0_101100010001;
      patterns[9058] = 29'b0_010001101100_010_0_100011011000;
      patterns[9059] = 29'b0_010001101100_011_1_000110110000;
      patterns[9060] = 29'b0_010001101100_100_0_001000110110;
      patterns[9061] = 29'b0_010001101100_101_0_000100011011;
      patterns[9062] = 29'b0_010001101100_110_0_010001101100;
      patterns[9063] = 29'b0_010001101100_111_0_010001101100;
      patterns[9064] = 29'b0_010001101101_000_0_010001101101;
      patterns[9065] = 29'b0_010001101101_001_0_101101010001;
      patterns[9066] = 29'b0_010001101101_010_0_100011011010;
      patterns[9067] = 29'b0_010001101101_011_1_000110110100;
      patterns[9068] = 29'b0_010001101101_100_1_001000110110;
      patterns[9069] = 29'b0_010001101101_101_0_100100011011;
      patterns[9070] = 29'b0_010001101101_110_0_010001101101;
      patterns[9071] = 29'b0_010001101101_111_0_010001101101;
      patterns[9072] = 29'b0_010001101110_000_0_010001101110;
      patterns[9073] = 29'b0_010001101110_001_0_101110010001;
      patterns[9074] = 29'b0_010001101110_010_0_100011011100;
      patterns[9075] = 29'b0_010001101110_011_1_000110111000;
      patterns[9076] = 29'b0_010001101110_100_0_001000110111;
      patterns[9077] = 29'b0_010001101110_101_1_000100011011;
      patterns[9078] = 29'b0_010001101110_110_0_010001101110;
      patterns[9079] = 29'b0_010001101110_111_0_010001101110;
      patterns[9080] = 29'b0_010001101111_000_0_010001101111;
      patterns[9081] = 29'b0_010001101111_001_0_101111010001;
      patterns[9082] = 29'b0_010001101111_010_0_100011011110;
      patterns[9083] = 29'b0_010001101111_011_1_000110111100;
      patterns[9084] = 29'b0_010001101111_100_1_001000110111;
      patterns[9085] = 29'b0_010001101111_101_1_100100011011;
      patterns[9086] = 29'b0_010001101111_110_0_010001101111;
      patterns[9087] = 29'b0_010001101111_111_0_010001101111;
      patterns[9088] = 29'b0_010001110000_000_0_010001110000;
      patterns[9089] = 29'b0_010001110000_001_0_110000010001;
      patterns[9090] = 29'b0_010001110000_010_0_100011100000;
      patterns[9091] = 29'b0_010001110000_011_1_000111000000;
      patterns[9092] = 29'b0_010001110000_100_0_001000111000;
      patterns[9093] = 29'b0_010001110000_101_0_000100011100;
      patterns[9094] = 29'b0_010001110000_110_0_010001110000;
      patterns[9095] = 29'b0_010001110000_111_0_010001110000;
      patterns[9096] = 29'b0_010001110001_000_0_010001110001;
      patterns[9097] = 29'b0_010001110001_001_0_110001010001;
      patterns[9098] = 29'b0_010001110001_010_0_100011100010;
      patterns[9099] = 29'b0_010001110001_011_1_000111000100;
      patterns[9100] = 29'b0_010001110001_100_1_001000111000;
      patterns[9101] = 29'b0_010001110001_101_0_100100011100;
      patterns[9102] = 29'b0_010001110001_110_0_010001110001;
      patterns[9103] = 29'b0_010001110001_111_0_010001110001;
      patterns[9104] = 29'b0_010001110010_000_0_010001110010;
      patterns[9105] = 29'b0_010001110010_001_0_110010010001;
      patterns[9106] = 29'b0_010001110010_010_0_100011100100;
      patterns[9107] = 29'b0_010001110010_011_1_000111001000;
      patterns[9108] = 29'b0_010001110010_100_0_001000111001;
      patterns[9109] = 29'b0_010001110010_101_1_000100011100;
      patterns[9110] = 29'b0_010001110010_110_0_010001110010;
      patterns[9111] = 29'b0_010001110010_111_0_010001110010;
      patterns[9112] = 29'b0_010001110011_000_0_010001110011;
      patterns[9113] = 29'b0_010001110011_001_0_110011010001;
      patterns[9114] = 29'b0_010001110011_010_0_100011100110;
      patterns[9115] = 29'b0_010001110011_011_1_000111001100;
      patterns[9116] = 29'b0_010001110011_100_1_001000111001;
      patterns[9117] = 29'b0_010001110011_101_1_100100011100;
      patterns[9118] = 29'b0_010001110011_110_0_010001110011;
      patterns[9119] = 29'b0_010001110011_111_0_010001110011;
      patterns[9120] = 29'b0_010001110100_000_0_010001110100;
      patterns[9121] = 29'b0_010001110100_001_0_110100010001;
      patterns[9122] = 29'b0_010001110100_010_0_100011101000;
      patterns[9123] = 29'b0_010001110100_011_1_000111010000;
      patterns[9124] = 29'b0_010001110100_100_0_001000111010;
      patterns[9125] = 29'b0_010001110100_101_0_000100011101;
      patterns[9126] = 29'b0_010001110100_110_0_010001110100;
      patterns[9127] = 29'b0_010001110100_111_0_010001110100;
      patterns[9128] = 29'b0_010001110101_000_0_010001110101;
      patterns[9129] = 29'b0_010001110101_001_0_110101010001;
      patterns[9130] = 29'b0_010001110101_010_0_100011101010;
      patterns[9131] = 29'b0_010001110101_011_1_000111010100;
      patterns[9132] = 29'b0_010001110101_100_1_001000111010;
      patterns[9133] = 29'b0_010001110101_101_0_100100011101;
      patterns[9134] = 29'b0_010001110101_110_0_010001110101;
      patterns[9135] = 29'b0_010001110101_111_0_010001110101;
      patterns[9136] = 29'b0_010001110110_000_0_010001110110;
      patterns[9137] = 29'b0_010001110110_001_0_110110010001;
      patterns[9138] = 29'b0_010001110110_010_0_100011101100;
      patterns[9139] = 29'b0_010001110110_011_1_000111011000;
      patterns[9140] = 29'b0_010001110110_100_0_001000111011;
      patterns[9141] = 29'b0_010001110110_101_1_000100011101;
      patterns[9142] = 29'b0_010001110110_110_0_010001110110;
      patterns[9143] = 29'b0_010001110110_111_0_010001110110;
      patterns[9144] = 29'b0_010001110111_000_0_010001110111;
      patterns[9145] = 29'b0_010001110111_001_0_110111010001;
      patterns[9146] = 29'b0_010001110111_010_0_100011101110;
      patterns[9147] = 29'b0_010001110111_011_1_000111011100;
      patterns[9148] = 29'b0_010001110111_100_1_001000111011;
      patterns[9149] = 29'b0_010001110111_101_1_100100011101;
      patterns[9150] = 29'b0_010001110111_110_0_010001110111;
      patterns[9151] = 29'b0_010001110111_111_0_010001110111;
      patterns[9152] = 29'b0_010001111000_000_0_010001111000;
      patterns[9153] = 29'b0_010001111000_001_0_111000010001;
      patterns[9154] = 29'b0_010001111000_010_0_100011110000;
      patterns[9155] = 29'b0_010001111000_011_1_000111100000;
      patterns[9156] = 29'b0_010001111000_100_0_001000111100;
      patterns[9157] = 29'b0_010001111000_101_0_000100011110;
      patterns[9158] = 29'b0_010001111000_110_0_010001111000;
      patterns[9159] = 29'b0_010001111000_111_0_010001111000;
      patterns[9160] = 29'b0_010001111001_000_0_010001111001;
      patterns[9161] = 29'b0_010001111001_001_0_111001010001;
      patterns[9162] = 29'b0_010001111001_010_0_100011110010;
      patterns[9163] = 29'b0_010001111001_011_1_000111100100;
      patterns[9164] = 29'b0_010001111001_100_1_001000111100;
      patterns[9165] = 29'b0_010001111001_101_0_100100011110;
      patterns[9166] = 29'b0_010001111001_110_0_010001111001;
      patterns[9167] = 29'b0_010001111001_111_0_010001111001;
      patterns[9168] = 29'b0_010001111010_000_0_010001111010;
      patterns[9169] = 29'b0_010001111010_001_0_111010010001;
      patterns[9170] = 29'b0_010001111010_010_0_100011110100;
      patterns[9171] = 29'b0_010001111010_011_1_000111101000;
      patterns[9172] = 29'b0_010001111010_100_0_001000111101;
      patterns[9173] = 29'b0_010001111010_101_1_000100011110;
      patterns[9174] = 29'b0_010001111010_110_0_010001111010;
      patterns[9175] = 29'b0_010001111010_111_0_010001111010;
      patterns[9176] = 29'b0_010001111011_000_0_010001111011;
      patterns[9177] = 29'b0_010001111011_001_0_111011010001;
      patterns[9178] = 29'b0_010001111011_010_0_100011110110;
      patterns[9179] = 29'b0_010001111011_011_1_000111101100;
      patterns[9180] = 29'b0_010001111011_100_1_001000111101;
      patterns[9181] = 29'b0_010001111011_101_1_100100011110;
      patterns[9182] = 29'b0_010001111011_110_0_010001111011;
      patterns[9183] = 29'b0_010001111011_111_0_010001111011;
      patterns[9184] = 29'b0_010001111100_000_0_010001111100;
      patterns[9185] = 29'b0_010001111100_001_0_111100010001;
      patterns[9186] = 29'b0_010001111100_010_0_100011111000;
      patterns[9187] = 29'b0_010001111100_011_1_000111110000;
      patterns[9188] = 29'b0_010001111100_100_0_001000111110;
      patterns[9189] = 29'b0_010001111100_101_0_000100011111;
      patterns[9190] = 29'b0_010001111100_110_0_010001111100;
      patterns[9191] = 29'b0_010001111100_111_0_010001111100;
      patterns[9192] = 29'b0_010001111101_000_0_010001111101;
      patterns[9193] = 29'b0_010001111101_001_0_111101010001;
      patterns[9194] = 29'b0_010001111101_010_0_100011111010;
      patterns[9195] = 29'b0_010001111101_011_1_000111110100;
      patterns[9196] = 29'b0_010001111101_100_1_001000111110;
      patterns[9197] = 29'b0_010001111101_101_0_100100011111;
      patterns[9198] = 29'b0_010001111101_110_0_010001111101;
      patterns[9199] = 29'b0_010001111101_111_0_010001111101;
      patterns[9200] = 29'b0_010001111110_000_0_010001111110;
      patterns[9201] = 29'b0_010001111110_001_0_111110010001;
      patterns[9202] = 29'b0_010001111110_010_0_100011111100;
      patterns[9203] = 29'b0_010001111110_011_1_000111111000;
      patterns[9204] = 29'b0_010001111110_100_0_001000111111;
      patterns[9205] = 29'b0_010001111110_101_1_000100011111;
      patterns[9206] = 29'b0_010001111110_110_0_010001111110;
      patterns[9207] = 29'b0_010001111110_111_0_010001111110;
      patterns[9208] = 29'b0_010001111111_000_0_010001111111;
      patterns[9209] = 29'b0_010001111111_001_0_111111010001;
      patterns[9210] = 29'b0_010001111111_010_0_100011111110;
      patterns[9211] = 29'b0_010001111111_011_1_000111111100;
      patterns[9212] = 29'b0_010001111111_100_1_001000111111;
      patterns[9213] = 29'b0_010001111111_101_1_100100011111;
      patterns[9214] = 29'b0_010001111111_110_0_010001111111;
      patterns[9215] = 29'b0_010001111111_111_0_010001111111;
      patterns[9216] = 29'b0_010010000000_000_0_010010000000;
      patterns[9217] = 29'b0_010010000000_001_0_000000010010;
      patterns[9218] = 29'b0_010010000000_010_0_100100000000;
      patterns[9219] = 29'b0_010010000000_011_1_001000000000;
      patterns[9220] = 29'b0_010010000000_100_0_001001000000;
      patterns[9221] = 29'b0_010010000000_101_0_000100100000;
      patterns[9222] = 29'b0_010010000000_110_0_010010000000;
      patterns[9223] = 29'b0_010010000000_111_0_010010000000;
      patterns[9224] = 29'b0_010010000001_000_0_010010000001;
      patterns[9225] = 29'b0_010010000001_001_0_000001010010;
      patterns[9226] = 29'b0_010010000001_010_0_100100000010;
      patterns[9227] = 29'b0_010010000001_011_1_001000000100;
      patterns[9228] = 29'b0_010010000001_100_1_001001000000;
      patterns[9229] = 29'b0_010010000001_101_0_100100100000;
      patterns[9230] = 29'b0_010010000001_110_0_010010000001;
      patterns[9231] = 29'b0_010010000001_111_0_010010000001;
      patterns[9232] = 29'b0_010010000010_000_0_010010000010;
      patterns[9233] = 29'b0_010010000010_001_0_000010010010;
      patterns[9234] = 29'b0_010010000010_010_0_100100000100;
      patterns[9235] = 29'b0_010010000010_011_1_001000001000;
      patterns[9236] = 29'b0_010010000010_100_0_001001000001;
      patterns[9237] = 29'b0_010010000010_101_1_000100100000;
      patterns[9238] = 29'b0_010010000010_110_0_010010000010;
      patterns[9239] = 29'b0_010010000010_111_0_010010000010;
      patterns[9240] = 29'b0_010010000011_000_0_010010000011;
      patterns[9241] = 29'b0_010010000011_001_0_000011010010;
      patterns[9242] = 29'b0_010010000011_010_0_100100000110;
      patterns[9243] = 29'b0_010010000011_011_1_001000001100;
      patterns[9244] = 29'b0_010010000011_100_1_001001000001;
      patterns[9245] = 29'b0_010010000011_101_1_100100100000;
      patterns[9246] = 29'b0_010010000011_110_0_010010000011;
      patterns[9247] = 29'b0_010010000011_111_0_010010000011;
      patterns[9248] = 29'b0_010010000100_000_0_010010000100;
      patterns[9249] = 29'b0_010010000100_001_0_000100010010;
      patterns[9250] = 29'b0_010010000100_010_0_100100001000;
      patterns[9251] = 29'b0_010010000100_011_1_001000010000;
      patterns[9252] = 29'b0_010010000100_100_0_001001000010;
      patterns[9253] = 29'b0_010010000100_101_0_000100100001;
      patterns[9254] = 29'b0_010010000100_110_0_010010000100;
      patterns[9255] = 29'b0_010010000100_111_0_010010000100;
      patterns[9256] = 29'b0_010010000101_000_0_010010000101;
      patterns[9257] = 29'b0_010010000101_001_0_000101010010;
      patterns[9258] = 29'b0_010010000101_010_0_100100001010;
      patterns[9259] = 29'b0_010010000101_011_1_001000010100;
      patterns[9260] = 29'b0_010010000101_100_1_001001000010;
      patterns[9261] = 29'b0_010010000101_101_0_100100100001;
      patterns[9262] = 29'b0_010010000101_110_0_010010000101;
      patterns[9263] = 29'b0_010010000101_111_0_010010000101;
      patterns[9264] = 29'b0_010010000110_000_0_010010000110;
      patterns[9265] = 29'b0_010010000110_001_0_000110010010;
      patterns[9266] = 29'b0_010010000110_010_0_100100001100;
      patterns[9267] = 29'b0_010010000110_011_1_001000011000;
      patterns[9268] = 29'b0_010010000110_100_0_001001000011;
      patterns[9269] = 29'b0_010010000110_101_1_000100100001;
      patterns[9270] = 29'b0_010010000110_110_0_010010000110;
      patterns[9271] = 29'b0_010010000110_111_0_010010000110;
      patterns[9272] = 29'b0_010010000111_000_0_010010000111;
      patterns[9273] = 29'b0_010010000111_001_0_000111010010;
      patterns[9274] = 29'b0_010010000111_010_0_100100001110;
      patterns[9275] = 29'b0_010010000111_011_1_001000011100;
      patterns[9276] = 29'b0_010010000111_100_1_001001000011;
      patterns[9277] = 29'b0_010010000111_101_1_100100100001;
      patterns[9278] = 29'b0_010010000111_110_0_010010000111;
      patterns[9279] = 29'b0_010010000111_111_0_010010000111;
      patterns[9280] = 29'b0_010010001000_000_0_010010001000;
      patterns[9281] = 29'b0_010010001000_001_0_001000010010;
      patterns[9282] = 29'b0_010010001000_010_0_100100010000;
      patterns[9283] = 29'b0_010010001000_011_1_001000100000;
      patterns[9284] = 29'b0_010010001000_100_0_001001000100;
      patterns[9285] = 29'b0_010010001000_101_0_000100100010;
      patterns[9286] = 29'b0_010010001000_110_0_010010001000;
      patterns[9287] = 29'b0_010010001000_111_0_010010001000;
      patterns[9288] = 29'b0_010010001001_000_0_010010001001;
      patterns[9289] = 29'b0_010010001001_001_0_001001010010;
      patterns[9290] = 29'b0_010010001001_010_0_100100010010;
      patterns[9291] = 29'b0_010010001001_011_1_001000100100;
      patterns[9292] = 29'b0_010010001001_100_1_001001000100;
      patterns[9293] = 29'b0_010010001001_101_0_100100100010;
      patterns[9294] = 29'b0_010010001001_110_0_010010001001;
      patterns[9295] = 29'b0_010010001001_111_0_010010001001;
      patterns[9296] = 29'b0_010010001010_000_0_010010001010;
      patterns[9297] = 29'b0_010010001010_001_0_001010010010;
      patterns[9298] = 29'b0_010010001010_010_0_100100010100;
      patterns[9299] = 29'b0_010010001010_011_1_001000101000;
      patterns[9300] = 29'b0_010010001010_100_0_001001000101;
      patterns[9301] = 29'b0_010010001010_101_1_000100100010;
      patterns[9302] = 29'b0_010010001010_110_0_010010001010;
      patterns[9303] = 29'b0_010010001010_111_0_010010001010;
      patterns[9304] = 29'b0_010010001011_000_0_010010001011;
      patterns[9305] = 29'b0_010010001011_001_0_001011010010;
      patterns[9306] = 29'b0_010010001011_010_0_100100010110;
      patterns[9307] = 29'b0_010010001011_011_1_001000101100;
      patterns[9308] = 29'b0_010010001011_100_1_001001000101;
      patterns[9309] = 29'b0_010010001011_101_1_100100100010;
      patterns[9310] = 29'b0_010010001011_110_0_010010001011;
      patterns[9311] = 29'b0_010010001011_111_0_010010001011;
      patterns[9312] = 29'b0_010010001100_000_0_010010001100;
      patterns[9313] = 29'b0_010010001100_001_0_001100010010;
      patterns[9314] = 29'b0_010010001100_010_0_100100011000;
      patterns[9315] = 29'b0_010010001100_011_1_001000110000;
      patterns[9316] = 29'b0_010010001100_100_0_001001000110;
      patterns[9317] = 29'b0_010010001100_101_0_000100100011;
      patterns[9318] = 29'b0_010010001100_110_0_010010001100;
      patterns[9319] = 29'b0_010010001100_111_0_010010001100;
      patterns[9320] = 29'b0_010010001101_000_0_010010001101;
      patterns[9321] = 29'b0_010010001101_001_0_001101010010;
      patterns[9322] = 29'b0_010010001101_010_0_100100011010;
      patterns[9323] = 29'b0_010010001101_011_1_001000110100;
      patterns[9324] = 29'b0_010010001101_100_1_001001000110;
      patterns[9325] = 29'b0_010010001101_101_0_100100100011;
      patterns[9326] = 29'b0_010010001101_110_0_010010001101;
      patterns[9327] = 29'b0_010010001101_111_0_010010001101;
      patterns[9328] = 29'b0_010010001110_000_0_010010001110;
      patterns[9329] = 29'b0_010010001110_001_0_001110010010;
      patterns[9330] = 29'b0_010010001110_010_0_100100011100;
      patterns[9331] = 29'b0_010010001110_011_1_001000111000;
      patterns[9332] = 29'b0_010010001110_100_0_001001000111;
      patterns[9333] = 29'b0_010010001110_101_1_000100100011;
      patterns[9334] = 29'b0_010010001110_110_0_010010001110;
      patterns[9335] = 29'b0_010010001110_111_0_010010001110;
      patterns[9336] = 29'b0_010010001111_000_0_010010001111;
      patterns[9337] = 29'b0_010010001111_001_0_001111010010;
      patterns[9338] = 29'b0_010010001111_010_0_100100011110;
      patterns[9339] = 29'b0_010010001111_011_1_001000111100;
      patterns[9340] = 29'b0_010010001111_100_1_001001000111;
      patterns[9341] = 29'b0_010010001111_101_1_100100100011;
      patterns[9342] = 29'b0_010010001111_110_0_010010001111;
      patterns[9343] = 29'b0_010010001111_111_0_010010001111;
      patterns[9344] = 29'b0_010010010000_000_0_010010010000;
      patterns[9345] = 29'b0_010010010000_001_0_010000010010;
      patterns[9346] = 29'b0_010010010000_010_0_100100100000;
      patterns[9347] = 29'b0_010010010000_011_1_001001000000;
      patterns[9348] = 29'b0_010010010000_100_0_001001001000;
      patterns[9349] = 29'b0_010010010000_101_0_000100100100;
      patterns[9350] = 29'b0_010010010000_110_0_010010010000;
      patterns[9351] = 29'b0_010010010000_111_0_010010010000;
      patterns[9352] = 29'b0_010010010001_000_0_010010010001;
      patterns[9353] = 29'b0_010010010001_001_0_010001010010;
      patterns[9354] = 29'b0_010010010001_010_0_100100100010;
      patterns[9355] = 29'b0_010010010001_011_1_001001000100;
      patterns[9356] = 29'b0_010010010001_100_1_001001001000;
      patterns[9357] = 29'b0_010010010001_101_0_100100100100;
      patterns[9358] = 29'b0_010010010001_110_0_010010010001;
      patterns[9359] = 29'b0_010010010001_111_0_010010010001;
      patterns[9360] = 29'b0_010010010010_000_0_010010010010;
      patterns[9361] = 29'b0_010010010010_001_0_010010010010;
      patterns[9362] = 29'b0_010010010010_010_0_100100100100;
      patterns[9363] = 29'b0_010010010010_011_1_001001001000;
      patterns[9364] = 29'b0_010010010010_100_0_001001001001;
      patterns[9365] = 29'b0_010010010010_101_1_000100100100;
      patterns[9366] = 29'b0_010010010010_110_0_010010010010;
      patterns[9367] = 29'b0_010010010010_111_0_010010010010;
      patterns[9368] = 29'b0_010010010011_000_0_010010010011;
      patterns[9369] = 29'b0_010010010011_001_0_010011010010;
      patterns[9370] = 29'b0_010010010011_010_0_100100100110;
      patterns[9371] = 29'b0_010010010011_011_1_001001001100;
      patterns[9372] = 29'b0_010010010011_100_1_001001001001;
      patterns[9373] = 29'b0_010010010011_101_1_100100100100;
      patterns[9374] = 29'b0_010010010011_110_0_010010010011;
      patterns[9375] = 29'b0_010010010011_111_0_010010010011;
      patterns[9376] = 29'b0_010010010100_000_0_010010010100;
      patterns[9377] = 29'b0_010010010100_001_0_010100010010;
      patterns[9378] = 29'b0_010010010100_010_0_100100101000;
      patterns[9379] = 29'b0_010010010100_011_1_001001010000;
      patterns[9380] = 29'b0_010010010100_100_0_001001001010;
      patterns[9381] = 29'b0_010010010100_101_0_000100100101;
      patterns[9382] = 29'b0_010010010100_110_0_010010010100;
      patterns[9383] = 29'b0_010010010100_111_0_010010010100;
      patterns[9384] = 29'b0_010010010101_000_0_010010010101;
      patterns[9385] = 29'b0_010010010101_001_0_010101010010;
      patterns[9386] = 29'b0_010010010101_010_0_100100101010;
      patterns[9387] = 29'b0_010010010101_011_1_001001010100;
      patterns[9388] = 29'b0_010010010101_100_1_001001001010;
      patterns[9389] = 29'b0_010010010101_101_0_100100100101;
      patterns[9390] = 29'b0_010010010101_110_0_010010010101;
      patterns[9391] = 29'b0_010010010101_111_0_010010010101;
      patterns[9392] = 29'b0_010010010110_000_0_010010010110;
      patterns[9393] = 29'b0_010010010110_001_0_010110010010;
      patterns[9394] = 29'b0_010010010110_010_0_100100101100;
      patterns[9395] = 29'b0_010010010110_011_1_001001011000;
      patterns[9396] = 29'b0_010010010110_100_0_001001001011;
      patterns[9397] = 29'b0_010010010110_101_1_000100100101;
      patterns[9398] = 29'b0_010010010110_110_0_010010010110;
      patterns[9399] = 29'b0_010010010110_111_0_010010010110;
      patterns[9400] = 29'b0_010010010111_000_0_010010010111;
      patterns[9401] = 29'b0_010010010111_001_0_010111010010;
      patterns[9402] = 29'b0_010010010111_010_0_100100101110;
      patterns[9403] = 29'b0_010010010111_011_1_001001011100;
      patterns[9404] = 29'b0_010010010111_100_1_001001001011;
      patterns[9405] = 29'b0_010010010111_101_1_100100100101;
      patterns[9406] = 29'b0_010010010111_110_0_010010010111;
      patterns[9407] = 29'b0_010010010111_111_0_010010010111;
      patterns[9408] = 29'b0_010010011000_000_0_010010011000;
      patterns[9409] = 29'b0_010010011000_001_0_011000010010;
      patterns[9410] = 29'b0_010010011000_010_0_100100110000;
      patterns[9411] = 29'b0_010010011000_011_1_001001100000;
      patterns[9412] = 29'b0_010010011000_100_0_001001001100;
      patterns[9413] = 29'b0_010010011000_101_0_000100100110;
      patterns[9414] = 29'b0_010010011000_110_0_010010011000;
      patterns[9415] = 29'b0_010010011000_111_0_010010011000;
      patterns[9416] = 29'b0_010010011001_000_0_010010011001;
      patterns[9417] = 29'b0_010010011001_001_0_011001010010;
      patterns[9418] = 29'b0_010010011001_010_0_100100110010;
      patterns[9419] = 29'b0_010010011001_011_1_001001100100;
      patterns[9420] = 29'b0_010010011001_100_1_001001001100;
      patterns[9421] = 29'b0_010010011001_101_0_100100100110;
      patterns[9422] = 29'b0_010010011001_110_0_010010011001;
      patterns[9423] = 29'b0_010010011001_111_0_010010011001;
      patterns[9424] = 29'b0_010010011010_000_0_010010011010;
      patterns[9425] = 29'b0_010010011010_001_0_011010010010;
      patterns[9426] = 29'b0_010010011010_010_0_100100110100;
      patterns[9427] = 29'b0_010010011010_011_1_001001101000;
      patterns[9428] = 29'b0_010010011010_100_0_001001001101;
      patterns[9429] = 29'b0_010010011010_101_1_000100100110;
      patterns[9430] = 29'b0_010010011010_110_0_010010011010;
      patterns[9431] = 29'b0_010010011010_111_0_010010011010;
      patterns[9432] = 29'b0_010010011011_000_0_010010011011;
      patterns[9433] = 29'b0_010010011011_001_0_011011010010;
      patterns[9434] = 29'b0_010010011011_010_0_100100110110;
      patterns[9435] = 29'b0_010010011011_011_1_001001101100;
      patterns[9436] = 29'b0_010010011011_100_1_001001001101;
      patterns[9437] = 29'b0_010010011011_101_1_100100100110;
      patterns[9438] = 29'b0_010010011011_110_0_010010011011;
      patterns[9439] = 29'b0_010010011011_111_0_010010011011;
      patterns[9440] = 29'b0_010010011100_000_0_010010011100;
      patterns[9441] = 29'b0_010010011100_001_0_011100010010;
      patterns[9442] = 29'b0_010010011100_010_0_100100111000;
      patterns[9443] = 29'b0_010010011100_011_1_001001110000;
      patterns[9444] = 29'b0_010010011100_100_0_001001001110;
      patterns[9445] = 29'b0_010010011100_101_0_000100100111;
      patterns[9446] = 29'b0_010010011100_110_0_010010011100;
      patterns[9447] = 29'b0_010010011100_111_0_010010011100;
      patterns[9448] = 29'b0_010010011101_000_0_010010011101;
      patterns[9449] = 29'b0_010010011101_001_0_011101010010;
      patterns[9450] = 29'b0_010010011101_010_0_100100111010;
      patterns[9451] = 29'b0_010010011101_011_1_001001110100;
      patterns[9452] = 29'b0_010010011101_100_1_001001001110;
      patterns[9453] = 29'b0_010010011101_101_0_100100100111;
      patterns[9454] = 29'b0_010010011101_110_0_010010011101;
      patterns[9455] = 29'b0_010010011101_111_0_010010011101;
      patterns[9456] = 29'b0_010010011110_000_0_010010011110;
      patterns[9457] = 29'b0_010010011110_001_0_011110010010;
      patterns[9458] = 29'b0_010010011110_010_0_100100111100;
      patterns[9459] = 29'b0_010010011110_011_1_001001111000;
      patterns[9460] = 29'b0_010010011110_100_0_001001001111;
      patterns[9461] = 29'b0_010010011110_101_1_000100100111;
      patterns[9462] = 29'b0_010010011110_110_0_010010011110;
      patterns[9463] = 29'b0_010010011110_111_0_010010011110;
      patterns[9464] = 29'b0_010010011111_000_0_010010011111;
      patterns[9465] = 29'b0_010010011111_001_0_011111010010;
      patterns[9466] = 29'b0_010010011111_010_0_100100111110;
      patterns[9467] = 29'b0_010010011111_011_1_001001111100;
      patterns[9468] = 29'b0_010010011111_100_1_001001001111;
      patterns[9469] = 29'b0_010010011111_101_1_100100100111;
      patterns[9470] = 29'b0_010010011111_110_0_010010011111;
      patterns[9471] = 29'b0_010010011111_111_0_010010011111;
      patterns[9472] = 29'b0_010010100000_000_0_010010100000;
      patterns[9473] = 29'b0_010010100000_001_0_100000010010;
      patterns[9474] = 29'b0_010010100000_010_0_100101000000;
      patterns[9475] = 29'b0_010010100000_011_1_001010000000;
      patterns[9476] = 29'b0_010010100000_100_0_001001010000;
      patterns[9477] = 29'b0_010010100000_101_0_000100101000;
      patterns[9478] = 29'b0_010010100000_110_0_010010100000;
      patterns[9479] = 29'b0_010010100000_111_0_010010100000;
      patterns[9480] = 29'b0_010010100001_000_0_010010100001;
      patterns[9481] = 29'b0_010010100001_001_0_100001010010;
      patterns[9482] = 29'b0_010010100001_010_0_100101000010;
      patterns[9483] = 29'b0_010010100001_011_1_001010000100;
      patterns[9484] = 29'b0_010010100001_100_1_001001010000;
      patterns[9485] = 29'b0_010010100001_101_0_100100101000;
      patterns[9486] = 29'b0_010010100001_110_0_010010100001;
      patterns[9487] = 29'b0_010010100001_111_0_010010100001;
      patterns[9488] = 29'b0_010010100010_000_0_010010100010;
      patterns[9489] = 29'b0_010010100010_001_0_100010010010;
      patterns[9490] = 29'b0_010010100010_010_0_100101000100;
      patterns[9491] = 29'b0_010010100010_011_1_001010001000;
      patterns[9492] = 29'b0_010010100010_100_0_001001010001;
      patterns[9493] = 29'b0_010010100010_101_1_000100101000;
      patterns[9494] = 29'b0_010010100010_110_0_010010100010;
      patterns[9495] = 29'b0_010010100010_111_0_010010100010;
      patterns[9496] = 29'b0_010010100011_000_0_010010100011;
      patterns[9497] = 29'b0_010010100011_001_0_100011010010;
      patterns[9498] = 29'b0_010010100011_010_0_100101000110;
      patterns[9499] = 29'b0_010010100011_011_1_001010001100;
      patterns[9500] = 29'b0_010010100011_100_1_001001010001;
      patterns[9501] = 29'b0_010010100011_101_1_100100101000;
      patterns[9502] = 29'b0_010010100011_110_0_010010100011;
      patterns[9503] = 29'b0_010010100011_111_0_010010100011;
      patterns[9504] = 29'b0_010010100100_000_0_010010100100;
      patterns[9505] = 29'b0_010010100100_001_0_100100010010;
      patterns[9506] = 29'b0_010010100100_010_0_100101001000;
      patterns[9507] = 29'b0_010010100100_011_1_001010010000;
      patterns[9508] = 29'b0_010010100100_100_0_001001010010;
      patterns[9509] = 29'b0_010010100100_101_0_000100101001;
      patterns[9510] = 29'b0_010010100100_110_0_010010100100;
      patterns[9511] = 29'b0_010010100100_111_0_010010100100;
      patterns[9512] = 29'b0_010010100101_000_0_010010100101;
      patterns[9513] = 29'b0_010010100101_001_0_100101010010;
      patterns[9514] = 29'b0_010010100101_010_0_100101001010;
      patterns[9515] = 29'b0_010010100101_011_1_001010010100;
      patterns[9516] = 29'b0_010010100101_100_1_001001010010;
      patterns[9517] = 29'b0_010010100101_101_0_100100101001;
      patterns[9518] = 29'b0_010010100101_110_0_010010100101;
      patterns[9519] = 29'b0_010010100101_111_0_010010100101;
      patterns[9520] = 29'b0_010010100110_000_0_010010100110;
      patterns[9521] = 29'b0_010010100110_001_0_100110010010;
      patterns[9522] = 29'b0_010010100110_010_0_100101001100;
      patterns[9523] = 29'b0_010010100110_011_1_001010011000;
      patterns[9524] = 29'b0_010010100110_100_0_001001010011;
      patterns[9525] = 29'b0_010010100110_101_1_000100101001;
      patterns[9526] = 29'b0_010010100110_110_0_010010100110;
      patterns[9527] = 29'b0_010010100110_111_0_010010100110;
      patterns[9528] = 29'b0_010010100111_000_0_010010100111;
      patterns[9529] = 29'b0_010010100111_001_0_100111010010;
      patterns[9530] = 29'b0_010010100111_010_0_100101001110;
      patterns[9531] = 29'b0_010010100111_011_1_001010011100;
      patterns[9532] = 29'b0_010010100111_100_1_001001010011;
      patterns[9533] = 29'b0_010010100111_101_1_100100101001;
      patterns[9534] = 29'b0_010010100111_110_0_010010100111;
      patterns[9535] = 29'b0_010010100111_111_0_010010100111;
      patterns[9536] = 29'b0_010010101000_000_0_010010101000;
      patterns[9537] = 29'b0_010010101000_001_0_101000010010;
      patterns[9538] = 29'b0_010010101000_010_0_100101010000;
      patterns[9539] = 29'b0_010010101000_011_1_001010100000;
      patterns[9540] = 29'b0_010010101000_100_0_001001010100;
      patterns[9541] = 29'b0_010010101000_101_0_000100101010;
      patterns[9542] = 29'b0_010010101000_110_0_010010101000;
      patterns[9543] = 29'b0_010010101000_111_0_010010101000;
      patterns[9544] = 29'b0_010010101001_000_0_010010101001;
      patterns[9545] = 29'b0_010010101001_001_0_101001010010;
      patterns[9546] = 29'b0_010010101001_010_0_100101010010;
      patterns[9547] = 29'b0_010010101001_011_1_001010100100;
      patterns[9548] = 29'b0_010010101001_100_1_001001010100;
      patterns[9549] = 29'b0_010010101001_101_0_100100101010;
      patterns[9550] = 29'b0_010010101001_110_0_010010101001;
      patterns[9551] = 29'b0_010010101001_111_0_010010101001;
      patterns[9552] = 29'b0_010010101010_000_0_010010101010;
      patterns[9553] = 29'b0_010010101010_001_0_101010010010;
      patterns[9554] = 29'b0_010010101010_010_0_100101010100;
      patterns[9555] = 29'b0_010010101010_011_1_001010101000;
      patterns[9556] = 29'b0_010010101010_100_0_001001010101;
      patterns[9557] = 29'b0_010010101010_101_1_000100101010;
      patterns[9558] = 29'b0_010010101010_110_0_010010101010;
      patterns[9559] = 29'b0_010010101010_111_0_010010101010;
      patterns[9560] = 29'b0_010010101011_000_0_010010101011;
      patterns[9561] = 29'b0_010010101011_001_0_101011010010;
      patterns[9562] = 29'b0_010010101011_010_0_100101010110;
      patterns[9563] = 29'b0_010010101011_011_1_001010101100;
      patterns[9564] = 29'b0_010010101011_100_1_001001010101;
      patterns[9565] = 29'b0_010010101011_101_1_100100101010;
      patterns[9566] = 29'b0_010010101011_110_0_010010101011;
      patterns[9567] = 29'b0_010010101011_111_0_010010101011;
      patterns[9568] = 29'b0_010010101100_000_0_010010101100;
      patterns[9569] = 29'b0_010010101100_001_0_101100010010;
      patterns[9570] = 29'b0_010010101100_010_0_100101011000;
      patterns[9571] = 29'b0_010010101100_011_1_001010110000;
      patterns[9572] = 29'b0_010010101100_100_0_001001010110;
      patterns[9573] = 29'b0_010010101100_101_0_000100101011;
      patterns[9574] = 29'b0_010010101100_110_0_010010101100;
      patterns[9575] = 29'b0_010010101100_111_0_010010101100;
      patterns[9576] = 29'b0_010010101101_000_0_010010101101;
      patterns[9577] = 29'b0_010010101101_001_0_101101010010;
      patterns[9578] = 29'b0_010010101101_010_0_100101011010;
      patterns[9579] = 29'b0_010010101101_011_1_001010110100;
      patterns[9580] = 29'b0_010010101101_100_1_001001010110;
      patterns[9581] = 29'b0_010010101101_101_0_100100101011;
      patterns[9582] = 29'b0_010010101101_110_0_010010101101;
      patterns[9583] = 29'b0_010010101101_111_0_010010101101;
      patterns[9584] = 29'b0_010010101110_000_0_010010101110;
      patterns[9585] = 29'b0_010010101110_001_0_101110010010;
      patterns[9586] = 29'b0_010010101110_010_0_100101011100;
      patterns[9587] = 29'b0_010010101110_011_1_001010111000;
      patterns[9588] = 29'b0_010010101110_100_0_001001010111;
      patterns[9589] = 29'b0_010010101110_101_1_000100101011;
      patterns[9590] = 29'b0_010010101110_110_0_010010101110;
      patterns[9591] = 29'b0_010010101110_111_0_010010101110;
      patterns[9592] = 29'b0_010010101111_000_0_010010101111;
      patterns[9593] = 29'b0_010010101111_001_0_101111010010;
      patterns[9594] = 29'b0_010010101111_010_0_100101011110;
      patterns[9595] = 29'b0_010010101111_011_1_001010111100;
      patterns[9596] = 29'b0_010010101111_100_1_001001010111;
      patterns[9597] = 29'b0_010010101111_101_1_100100101011;
      patterns[9598] = 29'b0_010010101111_110_0_010010101111;
      patterns[9599] = 29'b0_010010101111_111_0_010010101111;
      patterns[9600] = 29'b0_010010110000_000_0_010010110000;
      patterns[9601] = 29'b0_010010110000_001_0_110000010010;
      patterns[9602] = 29'b0_010010110000_010_0_100101100000;
      patterns[9603] = 29'b0_010010110000_011_1_001011000000;
      patterns[9604] = 29'b0_010010110000_100_0_001001011000;
      patterns[9605] = 29'b0_010010110000_101_0_000100101100;
      patterns[9606] = 29'b0_010010110000_110_0_010010110000;
      patterns[9607] = 29'b0_010010110000_111_0_010010110000;
      patterns[9608] = 29'b0_010010110001_000_0_010010110001;
      patterns[9609] = 29'b0_010010110001_001_0_110001010010;
      patterns[9610] = 29'b0_010010110001_010_0_100101100010;
      patterns[9611] = 29'b0_010010110001_011_1_001011000100;
      patterns[9612] = 29'b0_010010110001_100_1_001001011000;
      patterns[9613] = 29'b0_010010110001_101_0_100100101100;
      patterns[9614] = 29'b0_010010110001_110_0_010010110001;
      patterns[9615] = 29'b0_010010110001_111_0_010010110001;
      patterns[9616] = 29'b0_010010110010_000_0_010010110010;
      patterns[9617] = 29'b0_010010110010_001_0_110010010010;
      patterns[9618] = 29'b0_010010110010_010_0_100101100100;
      patterns[9619] = 29'b0_010010110010_011_1_001011001000;
      patterns[9620] = 29'b0_010010110010_100_0_001001011001;
      patterns[9621] = 29'b0_010010110010_101_1_000100101100;
      patterns[9622] = 29'b0_010010110010_110_0_010010110010;
      patterns[9623] = 29'b0_010010110010_111_0_010010110010;
      patterns[9624] = 29'b0_010010110011_000_0_010010110011;
      patterns[9625] = 29'b0_010010110011_001_0_110011010010;
      patterns[9626] = 29'b0_010010110011_010_0_100101100110;
      patterns[9627] = 29'b0_010010110011_011_1_001011001100;
      patterns[9628] = 29'b0_010010110011_100_1_001001011001;
      patterns[9629] = 29'b0_010010110011_101_1_100100101100;
      patterns[9630] = 29'b0_010010110011_110_0_010010110011;
      patterns[9631] = 29'b0_010010110011_111_0_010010110011;
      patterns[9632] = 29'b0_010010110100_000_0_010010110100;
      patterns[9633] = 29'b0_010010110100_001_0_110100010010;
      patterns[9634] = 29'b0_010010110100_010_0_100101101000;
      patterns[9635] = 29'b0_010010110100_011_1_001011010000;
      patterns[9636] = 29'b0_010010110100_100_0_001001011010;
      patterns[9637] = 29'b0_010010110100_101_0_000100101101;
      patterns[9638] = 29'b0_010010110100_110_0_010010110100;
      patterns[9639] = 29'b0_010010110100_111_0_010010110100;
      patterns[9640] = 29'b0_010010110101_000_0_010010110101;
      patterns[9641] = 29'b0_010010110101_001_0_110101010010;
      patterns[9642] = 29'b0_010010110101_010_0_100101101010;
      patterns[9643] = 29'b0_010010110101_011_1_001011010100;
      patterns[9644] = 29'b0_010010110101_100_1_001001011010;
      patterns[9645] = 29'b0_010010110101_101_0_100100101101;
      patterns[9646] = 29'b0_010010110101_110_0_010010110101;
      patterns[9647] = 29'b0_010010110101_111_0_010010110101;
      patterns[9648] = 29'b0_010010110110_000_0_010010110110;
      patterns[9649] = 29'b0_010010110110_001_0_110110010010;
      patterns[9650] = 29'b0_010010110110_010_0_100101101100;
      patterns[9651] = 29'b0_010010110110_011_1_001011011000;
      patterns[9652] = 29'b0_010010110110_100_0_001001011011;
      patterns[9653] = 29'b0_010010110110_101_1_000100101101;
      patterns[9654] = 29'b0_010010110110_110_0_010010110110;
      patterns[9655] = 29'b0_010010110110_111_0_010010110110;
      patterns[9656] = 29'b0_010010110111_000_0_010010110111;
      patterns[9657] = 29'b0_010010110111_001_0_110111010010;
      patterns[9658] = 29'b0_010010110111_010_0_100101101110;
      patterns[9659] = 29'b0_010010110111_011_1_001011011100;
      patterns[9660] = 29'b0_010010110111_100_1_001001011011;
      patterns[9661] = 29'b0_010010110111_101_1_100100101101;
      patterns[9662] = 29'b0_010010110111_110_0_010010110111;
      patterns[9663] = 29'b0_010010110111_111_0_010010110111;
      patterns[9664] = 29'b0_010010111000_000_0_010010111000;
      patterns[9665] = 29'b0_010010111000_001_0_111000010010;
      patterns[9666] = 29'b0_010010111000_010_0_100101110000;
      patterns[9667] = 29'b0_010010111000_011_1_001011100000;
      patterns[9668] = 29'b0_010010111000_100_0_001001011100;
      patterns[9669] = 29'b0_010010111000_101_0_000100101110;
      patterns[9670] = 29'b0_010010111000_110_0_010010111000;
      patterns[9671] = 29'b0_010010111000_111_0_010010111000;
      patterns[9672] = 29'b0_010010111001_000_0_010010111001;
      patterns[9673] = 29'b0_010010111001_001_0_111001010010;
      patterns[9674] = 29'b0_010010111001_010_0_100101110010;
      patterns[9675] = 29'b0_010010111001_011_1_001011100100;
      patterns[9676] = 29'b0_010010111001_100_1_001001011100;
      patterns[9677] = 29'b0_010010111001_101_0_100100101110;
      patterns[9678] = 29'b0_010010111001_110_0_010010111001;
      patterns[9679] = 29'b0_010010111001_111_0_010010111001;
      patterns[9680] = 29'b0_010010111010_000_0_010010111010;
      patterns[9681] = 29'b0_010010111010_001_0_111010010010;
      patterns[9682] = 29'b0_010010111010_010_0_100101110100;
      patterns[9683] = 29'b0_010010111010_011_1_001011101000;
      patterns[9684] = 29'b0_010010111010_100_0_001001011101;
      patterns[9685] = 29'b0_010010111010_101_1_000100101110;
      patterns[9686] = 29'b0_010010111010_110_0_010010111010;
      patterns[9687] = 29'b0_010010111010_111_0_010010111010;
      patterns[9688] = 29'b0_010010111011_000_0_010010111011;
      patterns[9689] = 29'b0_010010111011_001_0_111011010010;
      patterns[9690] = 29'b0_010010111011_010_0_100101110110;
      patterns[9691] = 29'b0_010010111011_011_1_001011101100;
      patterns[9692] = 29'b0_010010111011_100_1_001001011101;
      patterns[9693] = 29'b0_010010111011_101_1_100100101110;
      patterns[9694] = 29'b0_010010111011_110_0_010010111011;
      patterns[9695] = 29'b0_010010111011_111_0_010010111011;
      patterns[9696] = 29'b0_010010111100_000_0_010010111100;
      patterns[9697] = 29'b0_010010111100_001_0_111100010010;
      patterns[9698] = 29'b0_010010111100_010_0_100101111000;
      patterns[9699] = 29'b0_010010111100_011_1_001011110000;
      patterns[9700] = 29'b0_010010111100_100_0_001001011110;
      patterns[9701] = 29'b0_010010111100_101_0_000100101111;
      patterns[9702] = 29'b0_010010111100_110_0_010010111100;
      patterns[9703] = 29'b0_010010111100_111_0_010010111100;
      patterns[9704] = 29'b0_010010111101_000_0_010010111101;
      patterns[9705] = 29'b0_010010111101_001_0_111101010010;
      patterns[9706] = 29'b0_010010111101_010_0_100101111010;
      patterns[9707] = 29'b0_010010111101_011_1_001011110100;
      patterns[9708] = 29'b0_010010111101_100_1_001001011110;
      patterns[9709] = 29'b0_010010111101_101_0_100100101111;
      patterns[9710] = 29'b0_010010111101_110_0_010010111101;
      patterns[9711] = 29'b0_010010111101_111_0_010010111101;
      patterns[9712] = 29'b0_010010111110_000_0_010010111110;
      patterns[9713] = 29'b0_010010111110_001_0_111110010010;
      patterns[9714] = 29'b0_010010111110_010_0_100101111100;
      patterns[9715] = 29'b0_010010111110_011_1_001011111000;
      patterns[9716] = 29'b0_010010111110_100_0_001001011111;
      patterns[9717] = 29'b0_010010111110_101_1_000100101111;
      patterns[9718] = 29'b0_010010111110_110_0_010010111110;
      patterns[9719] = 29'b0_010010111110_111_0_010010111110;
      patterns[9720] = 29'b0_010010111111_000_0_010010111111;
      patterns[9721] = 29'b0_010010111111_001_0_111111010010;
      patterns[9722] = 29'b0_010010111111_010_0_100101111110;
      patterns[9723] = 29'b0_010010111111_011_1_001011111100;
      patterns[9724] = 29'b0_010010111111_100_1_001001011111;
      patterns[9725] = 29'b0_010010111111_101_1_100100101111;
      patterns[9726] = 29'b0_010010111111_110_0_010010111111;
      patterns[9727] = 29'b0_010010111111_111_0_010010111111;
      patterns[9728] = 29'b0_010011000000_000_0_010011000000;
      patterns[9729] = 29'b0_010011000000_001_0_000000010011;
      patterns[9730] = 29'b0_010011000000_010_0_100110000000;
      patterns[9731] = 29'b0_010011000000_011_1_001100000000;
      patterns[9732] = 29'b0_010011000000_100_0_001001100000;
      patterns[9733] = 29'b0_010011000000_101_0_000100110000;
      patterns[9734] = 29'b0_010011000000_110_0_010011000000;
      patterns[9735] = 29'b0_010011000000_111_0_010011000000;
      patterns[9736] = 29'b0_010011000001_000_0_010011000001;
      patterns[9737] = 29'b0_010011000001_001_0_000001010011;
      patterns[9738] = 29'b0_010011000001_010_0_100110000010;
      patterns[9739] = 29'b0_010011000001_011_1_001100000100;
      patterns[9740] = 29'b0_010011000001_100_1_001001100000;
      patterns[9741] = 29'b0_010011000001_101_0_100100110000;
      patterns[9742] = 29'b0_010011000001_110_0_010011000001;
      patterns[9743] = 29'b0_010011000001_111_0_010011000001;
      patterns[9744] = 29'b0_010011000010_000_0_010011000010;
      patterns[9745] = 29'b0_010011000010_001_0_000010010011;
      patterns[9746] = 29'b0_010011000010_010_0_100110000100;
      patterns[9747] = 29'b0_010011000010_011_1_001100001000;
      patterns[9748] = 29'b0_010011000010_100_0_001001100001;
      patterns[9749] = 29'b0_010011000010_101_1_000100110000;
      patterns[9750] = 29'b0_010011000010_110_0_010011000010;
      patterns[9751] = 29'b0_010011000010_111_0_010011000010;
      patterns[9752] = 29'b0_010011000011_000_0_010011000011;
      patterns[9753] = 29'b0_010011000011_001_0_000011010011;
      patterns[9754] = 29'b0_010011000011_010_0_100110000110;
      patterns[9755] = 29'b0_010011000011_011_1_001100001100;
      patterns[9756] = 29'b0_010011000011_100_1_001001100001;
      patterns[9757] = 29'b0_010011000011_101_1_100100110000;
      patterns[9758] = 29'b0_010011000011_110_0_010011000011;
      patterns[9759] = 29'b0_010011000011_111_0_010011000011;
      patterns[9760] = 29'b0_010011000100_000_0_010011000100;
      patterns[9761] = 29'b0_010011000100_001_0_000100010011;
      patterns[9762] = 29'b0_010011000100_010_0_100110001000;
      patterns[9763] = 29'b0_010011000100_011_1_001100010000;
      patterns[9764] = 29'b0_010011000100_100_0_001001100010;
      patterns[9765] = 29'b0_010011000100_101_0_000100110001;
      patterns[9766] = 29'b0_010011000100_110_0_010011000100;
      patterns[9767] = 29'b0_010011000100_111_0_010011000100;
      patterns[9768] = 29'b0_010011000101_000_0_010011000101;
      patterns[9769] = 29'b0_010011000101_001_0_000101010011;
      patterns[9770] = 29'b0_010011000101_010_0_100110001010;
      patterns[9771] = 29'b0_010011000101_011_1_001100010100;
      patterns[9772] = 29'b0_010011000101_100_1_001001100010;
      patterns[9773] = 29'b0_010011000101_101_0_100100110001;
      patterns[9774] = 29'b0_010011000101_110_0_010011000101;
      patterns[9775] = 29'b0_010011000101_111_0_010011000101;
      patterns[9776] = 29'b0_010011000110_000_0_010011000110;
      patterns[9777] = 29'b0_010011000110_001_0_000110010011;
      patterns[9778] = 29'b0_010011000110_010_0_100110001100;
      patterns[9779] = 29'b0_010011000110_011_1_001100011000;
      patterns[9780] = 29'b0_010011000110_100_0_001001100011;
      patterns[9781] = 29'b0_010011000110_101_1_000100110001;
      patterns[9782] = 29'b0_010011000110_110_0_010011000110;
      patterns[9783] = 29'b0_010011000110_111_0_010011000110;
      patterns[9784] = 29'b0_010011000111_000_0_010011000111;
      patterns[9785] = 29'b0_010011000111_001_0_000111010011;
      patterns[9786] = 29'b0_010011000111_010_0_100110001110;
      patterns[9787] = 29'b0_010011000111_011_1_001100011100;
      patterns[9788] = 29'b0_010011000111_100_1_001001100011;
      patterns[9789] = 29'b0_010011000111_101_1_100100110001;
      patterns[9790] = 29'b0_010011000111_110_0_010011000111;
      patterns[9791] = 29'b0_010011000111_111_0_010011000111;
      patterns[9792] = 29'b0_010011001000_000_0_010011001000;
      patterns[9793] = 29'b0_010011001000_001_0_001000010011;
      patterns[9794] = 29'b0_010011001000_010_0_100110010000;
      patterns[9795] = 29'b0_010011001000_011_1_001100100000;
      patterns[9796] = 29'b0_010011001000_100_0_001001100100;
      patterns[9797] = 29'b0_010011001000_101_0_000100110010;
      patterns[9798] = 29'b0_010011001000_110_0_010011001000;
      patterns[9799] = 29'b0_010011001000_111_0_010011001000;
      patterns[9800] = 29'b0_010011001001_000_0_010011001001;
      patterns[9801] = 29'b0_010011001001_001_0_001001010011;
      patterns[9802] = 29'b0_010011001001_010_0_100110010010;
      patterns[9803] = 29'b0_010011001001_011_1_001100100100;
      patterns[9804] = 29'b0_010011001001_100_1_001001100100;
      patterns[9805] = 29'b0_010011001001_101_0_100100110010;
      patterns[9806] = 29'b0_010011001001_110_0_010011001001;
      patterns[9807] = 29'b0_010011001001_111_0_010011001001;
      patterns[9808] = 29'b0_010011001010_000_0_010011001010;
      patterns[9809] = 29'b0_010011001010_001_0_001010010011;
      patterns[9810] = 29'b0_010011001010_010_0_100110010100;
      patterns[9811] = 29'b0_010011001010_011_1_001100101000;
      patterns[9812] = 29'b0_010011001010_100_0_001001100101;
      patterns[9813] = 29'b0_010011001010_101_1_000100110010;
      patterns[9814] = 29'b0_010011001010_110_0_010011001010;
      patterns[9815] = 29'b0_010011001010_111_0_010011001010;
      patterns[9816] = 29'b0_010011001011_000_0_010011001011;
      patterns[9817] = 29'b0_010011001011_001_0_001011010011;
      patterns[9818] = 29'b0_010011001011_010_0_100110010110;
      patterns[9819] = 29'b0_010011001011_011_1_001100101100;
      patterns[9820] = 29'b0_010011001011_100_1_001001100101;
      patterns[9821] = 29'b0_010011001011_101_1_100100110010;
      patterns[9822] = 29'b0_010011001011_110_0_010011001011;
      patterns[9823] = 29'b0_010011001011_111_0_010011001011;
      patterns[9824] = 29'b0_010011001100_000_0_010011001100;
      patterns[9825] = 29'b0_010011001100_001_0_001100010011;
      patterns[9826] = 29'b0_010011001100_010_0_100110011000;
      patterns[9827] = 29'b0_010011001100_011_1_001100110000;
      patterns[9828] = 29'b0_010011001100_100_0_001001100110;
      patterns[9829] = 29'b0_010011001100_101_0_000100110011;
      patterns[9830] = 29'b0_010011001100_110_0_010011001100;
      patterns[9831] = 29'b0_010011001100_111_0_010011001100;
      patterns[9832] = 29'b0_010011001101_000_0_010011001101;
      patterns[9833] = 29'b0_010011001101_001_0_001101010011;
      patterns[9834] = 29'b0_010011001101_010_0_100110011010;
      patterns[9835] = 29'b0_010011001101_011_1_001100110100;
      patterns[9836] = 29'b0_010011001101_100_1_001001100110;
      patterns[9837] = 29'b0_010011001101_101_0_100100110011;
      patterns[9838] = 29'b0_010011001101_110_0_010011001101;
      patterns[9839] = 29'b0_010011001101_111_0_010011001101;
      patterns[9840] = 29'b0_010011001110_000_0_010011001110;
      patterns[9841] = 29'b0_010011001110_001_0_001110010011;
      patterns[9842] = 29'b0_010011001110_010_0_100110011100;
      patterns[9843] = 29'b0_010011001110_011_1_001100111000;
      patterns[9844] = 29'b0_010011001110_100_0_001001100111;
      patterns[9845] = 29'b0_010011001110_101_1_000100110011;
      patterns[9846] = 29'b0_010011001110_110_0_010011001110;
      patterns[9847] = 29'b0_010011001110_111_0_010011001110;
      patterns[9848] = 29'b0_010011001111_000_0_010011001111;
      patterns[9849] = 29'b0_010011001111_001_0_001111010011;
      patterns[9850] = 29'b0_010011001111_010_0_100110011110;
      patterns[9851] = 29'b0_010011001111_011_1_001100111100;
      patterns[9852] = 29'b0_010011001111_100_1_001001100111;
      patterns[9853] = 29'b0_010011001111_101_1_100100110011;
      patterns[9854] = 29'b0_010011001111_110_0_010011001111;
      patterns[9855] = 29'b0_010011001111_111_0_010011001111;
      patterns[9856] = 29'b0_010011010000_000_0_010011010000;
      patterns[9857] = 29'b0_010011010000_001_0_010000010011;
      patterns[9858] = 29'b0_010011010000_010_0_100110100000;
      patterns[9859] = 29'b0_010011010000_011_1_001101000000;
      patterns[9860] = 29'b0_010011010000_100_0_001001101000;
      patterns[9861] = 29'b0_010011010000_101_0_000100110100;
      patterns[9862] = 29'b0_010011010000_110_0_010011010000;
      patterns[9863] = 29'b0_010011010000_111_0_010011010000;
      patterns[9864] = 29'b0_010011010001_000_0_010011010001;
      patterns[9865] = 29'b0_010011010001_001_0_010001010011;
      patterns[9866] = 29'b0_010011010001_010_0_100110100010;
      patterns[9867] = 29'b0_010011010001_011_1_001101000100;
      patterns[9868] = 29'b0_010011010001_100_1_001001101000;
      patterns[9869] = 29'b0_010011010001_101_0_100100110100;
      patterns[9870] = 29'b0_010011010001_110_0_010011010001;
      patterns[9871] = 29'b0_010011010001_111_0_010011010001;
      patterns[9872] = 29'b0_010011010010_000_0_010011010010;
      patterns[9873] = 29'b0_010011010010_001_0_010010010011;
      patterns[9874] = 29'b0_010011010010_010_0_100110100100;
      patterns[9875] = 29'b0_010011010010_011_1_001101001000;
      patterns[9876] = 29'b0_010011010010_100_0_001001101001;
      patterns[9877] = 29'b0_010011010010_101_1_000100110100;
      patterns[9878] = 29'b0_010011010010_110_0_010011010010;
      patterns[9879] = 29'b0_010011010010_111_0_010011010010;
      patterns[9880] = 29'b0_010011010011_000_0_010011010011;
      patterns[9881] = 29'b0_010011010011_001_0_010011010011;
      patterns[9882] = 29'b0_010011010011_010_0_100110100110;
      patterns[9883] = 29'b0_010011010011_011_1_001101001100;
      patterns[9884] = 29'b0_010011010011_100_1_001001101001;
      patterns[9885] = 29'b0_010011010011_101_1_100100110100;
      patterns[9886] = 29'b0_010011010011_110_0_010011010011;
      patterns[9887] = 29'b0_010011010011_111_0_010011010011;
      patterns[9888] = 29'b0_010011010100_000_0_010011010100;
      patterns[9889] = 29'b0_010011010100_001_0_010100010011;
      patterns[9890] = 29'b0_010011010100_010_0_100110101000;
      patterns[9891] = 29'b0_010011010100_011_1_001101010000;
      patterns[9892] = 29'b0_010011010100_100_0_001001101010;
      patterns[9893] = 29'b0_010011010100_101_0_000100110101;
      patterns[9894] = 29'b0_010011010100_110_0_010011010100;
      patterns[9895] = 29'b0_010011010100_111_0_010011010100;
      patterns[9896] = 29'b0_010011010101_000_0_010011010101;
      patterns[9897] = 29'b0_010011010101_001_0_010101010011;
      patterns[9898] = 29'b0_010011010101_010_0_100110101010;
      patterns[9899] = 29'b0_010011010101_011_1_001101010100;
      patterns[9900] = 29'b0_010011010101_100_1_001001101010;
      patterns[9901] = 29'b0_010011010101_101_0_100100110101;
      patterns[9902] = 29'b0_010011010101_110_0_010011010101;
      patterns[9903] = 29'b0_010011010101_111_0_010011010101;
      patterns[9904] = 29'b0_010011010110_000_0_010011010110;
      patterns[9905] = 29'b0_010011010110_001_0_010110010011;
      patterns[9906] = 29'b0_010011010110_010_0_100110101100;
      patterns[9907] = 29'b0_010011010110_011_1_001101011000;
      patterns[9908] = 29'b0_010011010110_100_0_001001101011;
      patterns[9909] = 29'b0_010011010110_101_1_000100110101;
      patterns[9910] = 29'b0_010011010110_110_0_010011010110;
      patterns[9911] = 29'b0_010011010110_111_0_010011010110;
      patterns[9912] = 29'b0_010011010111_000_0_010011010111;
      patterns[9913] = 29'b0_010011010111_001_0_010111010011;
      patterns[9914] = 29'b0_010011010111_010_0_100110101110;
      patterns[9915] = 29'b0_010011010111_011_1_001101011100;
      patterns[9916] = 29'b0_010011010111_100_1_001001101011;
      patterns[9917] = 29'b0_010011010111_101_1_100100110101;
      patterns[9918] = 29'b0_010011010111_110_0_010011010111;
      patterns[9919] = 29'b0_010011010111_111_0_010011010111;
      patterns[9920] = 29'b0_010011011000_000_0_010011011000;
      patterns[9921] = 29'b0_010011011000_001_0_011000010011;
      patterns[9922] = 29'b0_010011011000_010_0_100110110000;
      patterns[9923] = 29'b0_010011011000_011_1_001101100000;
      patterns[9924] = 29'b0_010011011000_100_0_001001101100;
      patterns[9925] = 29'b0_010011011000_101_0_000100110110;
      patterns[9926] = 29'b0_010011011000_110_0_010011011000;
      patterns[9927] = 29'b0_010011011000_111_0_010011011000;
      patterns[9928] = 29'b0_010011011001_000_0_010011011001;
      patterns[9929] = 29'b0_010011011001_001_0_011001010011;
      patterns[9930] = 29'b0_010011011001_010_0_100110110010;
      patterns[9931] = 29'b0_010011011001_011_1_001101100100;
      patterns[9932] = 29'b0_010011011001_100_1_001001101100;
      patterns[9933] = 29'b0_010011011001_101_0_100100110110;
      patterns[9934] = 29'b0_010011011001_110_0_010011011001;
      patterns[9935] = 29'b0_010011011001_111_0_010011011001;
      patterns[9936] = 29'b0_010011011010_000_0_010011011010;
      patterns[9937] = 29'b0_010011011010_001_0_011010010011;
      patterns[9938] = 29'b0_010011011010_010_0_100110110100;
      patterns[9939] = 29'b0_010011011010_011_1_001101101000;
      patterns[9940] = 29'b0_010011011010_100_0_001001101101;
      patterns[9941] = 29'b0_010011011010_101_1_000100110110;
      patterns[9942] = 29'b0_010011011010_110_0_010011011010;
      patterns[9943] = 29'b0_010011011010_111_0_010011011010;
      patterns[9944] = 29'b0_010011011011_000_0_010011011011;
      patterns[9945] = 29'b0_010011011011_001_0_011011010011;
      patterns[9946] = 29'b0_010011011011_010_0_100110110110;
      patterns[9947] = 29'b0_010011011011_011_1_001101101100;
      patterns[9948] = 29'b0_010011011011_100_1_001001101101;
      patterns[9949] = 29'b0_010011011011_101_1_100100110110;
      patterns[9950] = 29'b0_010011011011_110_0_010011011011;
      patterns[9951] = 29'b0_010011011011_111_0_010011011011;
      patterns[9952] = 29'b0_010011011100_000_0_010011011100;
      patterns[9953] = 29'b0_010011011100_001_0_011100010011;
      patterns[9954] = 29'b0_010011011100_010_0_100110111000;
      patterns[9955] = 29'b0_010011011100_011_1_001101110000;
      patterns[9956] = 29'b0_010011011100_100_0_001001101110;
      patterns[9957] = 29'b0_010011011100_101_0_000100110111;
      patterns[9958] = 29'b0_010011011100_110_0_010011011100;
      patterns[9959] = 29'b0_010011011100_111_0_010011011100;
      patterns[9960] = 29'b0_010011011101_000_0_010011011101;
      patterns[9961] = 29'b0_010011011101_001_0_011101010011;
      patterns[9962] = 29'b0_010011011101_010_0_100110111010;
      patterns[9963] = 29'b0_010011011101_011_1_001101110100;
      patterns[9964] = 29'b0_010011011101_100_1_001001101110;
      patterns[9965] = 29'b0_010011011101_101_0_100100110111;
      patterns[9966] = 29'b0_010011011101_110_0_010011011101;
      patterns[9967] = 29'b0_010011011101_111_0_010011011101;
      patterns[9968] = 29'b0_010011011110_000_0_010011011110;
      patterns[9969] = 29'b0_010011011110_001_0_011110010011;
      patterns[9970] = 29'b0_010011011110_010_0_100110111100;
      patterns[9971] = 29'b0_010011011110_011_1_001101111000;
      patterns[9972] = 29'b0_010011011110_100_0_001001101111;
      patterns[9973] = 29'b0_010011011110_101_1_000100110111;
      patterns[9974] = 29'b0_010011011110_110_0_010011011110;
      patterns[9975] = 29'b0_010011011110_111_0_010011011110;
      patterns[9976] = 29'b0_010011011111_000_0_010011011111;
      patterns[9977] = 29'b0_010011011111_001_0_011111010011;
      patterns[9978] = 29'b0_010011011111_010_0_100110111110;
      patterns[9979] = 29'b0_010011011111_011_1_001101111100;
      patterns[9980] = 29'b0_010011011111_100_1_001001101111;
      patterns[9981] = 29'b0_010011011111_101_1_100100110111;
      patterns[9982] = 29'b0_010011011111_110_0_010011011111;
      patterns[9983] = 29'b0_010011011111_111_0_010011011111;
      patterns[9984] = 29'b0_010011100000_000_0_010011100000;
      patterns[9985] = 29'b0_010011100000_001_0_100000010011;
      patterns[9986] = 29'b0_010011100000_010_0_100111000000;
      patterns[9987] = 29'b0_010011100000_011_1_001110000000;
      patterns[9988] = 29'b0_010011100000_100_0_001001110000;
      patterns[9989] = 29'b0_010011100000_101_0_000100111000;
      patterns[9990] = 29'b0_010011100000_110_0_010011100000;
      patterns[9991] = 29'b0_010011100000_111_0_010011100000;
      patterns[9992] = 29'b0_010011100001_000_0_010011100001;
      patterns[9993] = 29'b0_010011100001_001_0_100001010011;
      patterns[9994] = 29'b0_010011100001_010_0_100111000010;
      patterns[9995] = 29'b0_010011100001_011_1_001110000100;
      patterns[9996] = 29'b0_010011100001_100_1_001001110000;
      patterns[9997] = 29'b0_010011100001_101_0_100100111000;
      patterns[9998] = 29'b0_010011100001_110_0_010011100001;
      patterns[9999] = 29'b0_010011100001_111_0_010011100001;
      patterns[10000] = 29'b0_010011100010_000_0_010011100010;
      patterns[10001] = 29'b0_010011100010_001_0_100010010011;
      patterns[10002] = 29'b0_010011100010_010_0_100111000100;
      patterns[10003] = 29'b0_010011100010_011_1_001110001000;
      patterns[10004] = 29'b0_010011100010_100_0_001001110001;
      patterns[10005] = 29'b0_010011100010_101_1_000100111000;
      patterns[10006] = 29'b0_010011100010_110_0_010011100010;
      patterns[10007] = 29'b0_010011100010_111_0_010011100010;
      patterns[10008] = 29'b0_010011100011_000_0_010011100011;
      patterns[10009] = 29'b0_010011100011_001_0_100011010011;
      patterns[10010] = 29'b0_010011100011_010_0_100111000110;
      patterns[10011] = 29'b0_010011100011_011_1_001110001100;
      patterns[10012] = 29'b0_010011100011_100_1_001001110001;
      patterns[10013] = 29'b0_010011100011_101_1_100100111000;
      patterns[10014] = 29'b0_010011100011_110_0_010011100011;
      patterns[10015] = 29'b0_010011100011_111_0_010011100011;
      patterns[10016] = 29'b0_010011100100_000_0_010011100100;
      patterns[10017] = 29'b0_010011100100_001_0_100100010011;
      patterns[10018] = 29'b0_010011100100_010_0_100111001000;
      patterns[10019] = 29'b0_010011100100_011_1_001110010000;
      patterns[10020] = 29'b0_010011100100_100_0_001001110010;
      patterns[10021] = 29'b0_010011100100_101_0_000100111001;
      patterns[10022] = 29'b0_010011100100_110_0_010011100100;
      patterns[10023] = 29'b0_010011100100_111_0_010011100100;
      patterns[10024] = 29'b0_010011100101_000_0_010011100101;
      patterns[10025] = 29'b0_010011100101_001_0_100101010011;
      patterns[10026] = 29'b0_010011100101_010_0_100111001010;
      patterns[10027] = 29'b0_010011100101_011_1_001110010100;
      patterns[10028] = 29'b0_010011100101_100_1_001001110010;
      patterns[10029] = 29'b0_010011100101_101_0_100100111001;
      patterns[10030] = 29'b0_010011100101_110_0_010011100101;
      patterns[10031] = 29'b0_010011100101_111_0_010011100101;
      patterns[10032] = 29'b0_010011100110_000_0_010011100110;
      patterns[10033] = 29'b0_010011100110_001_0_100110010011;
      patterns[10034] = 29'b0_010011100110_010_0_100111001100;
      patterns[10035] = 29'b0_010011100110_011_1_001110011000;
      patterns[10036] = 29'b0_010011100110_100_0_001001110011;
      patterns[10037] = 29'b0_010011100110_101_1_000100111001;
      patterns[10038] = 29'b0_010011100110_110_0_010011100110;
      patterns[10039] = 29'b0_010011100110_111_0_010011100110;
      patterns[10040] = 29'b0_010011100111_000_0_010011100111;
      patterns[10041] = 29'b0_010011100111_001_0_100111010011;
      patterns[10042] = 29'b0_010011100111_010_0_100111001110;
      patterns[10043] = 29'b0_010011100111_011_1_001110011100;
      patterns[10044] = 29'b0_010011100111_100_1_001001110011;
      patterns[10045] = 29'b0_010011100111_101_1_100100111001;
      patterns[10046] = 29'b0_010011100111_110_0_010011100111;
      patterns[10047] = 29'b0_010011100111_111_0_010011100111;
      patterns[10048] = 29'b0_010011101000_000_0_010011101000;
      patterns[10049] = 29'b0_010011101000_001_0_101000010011;
      patterns[10050] = 29'b0_010011101000_010_0_100111010000;
      patterns[10051] = 29'b0_010011101000_011_1_001110100000;
      patterns[10052] = 29'b0_010011101000_100_0_001001110100;
      patterns[10053] = 29'b0_010011101000_101_0_000100111010;
      patterns[10054] = 29'b0_010011101000_110_0_010011101000;
      patterns[10055] = 29'b0_010011101000_111_0_010011101000;
      patterns[10056] = 29'b0_010011101001_000_0_010011101001;
      patterns[10057] = 29'b0_010011101001_001_0_101001010011;
      patterns[10058] = 29'b0_010011101001_010_0_100111010010;
      patterns[10059] = 29'b0_010011101001_011_1_001110100100;
      patterns[10060] = 29'b0_010011101001_100_1_001001110100;
      patterns[10061] = 29'b0_010011101001_101_0_100100111010;
      patterns[10062] = 29'b0_010011101001_110_0_010011101001;
      patterns[10063] = 29'b0_010011101001_111_0_010011101001;
      patterns[10064] = 29'b0_010011101010_000_0_010011101010;
      patterns[10065] = 29'b0_010011101010_001_0_101010010011;
      patterns[10066] = 29'b0_010011101010_010_0_100111010100;
      patterns[10067] = 29'b0_010011101010_011_1_001110101000;
      patterns[10068] = 29'b0_010011101010_100_0_001001110101;
      patterns[10069] = 29'b0_010011101010_101_1_000100111010;
      patterns[10070] = 29'b0_010011101010_110_0_010011101010;
      patterns[10071] = 29'b0_010011101010_111_0_010011101010;
      patterns[10072] = 29'b0_010011101011_000_0_010011101011;
      patterns[10073] = 29'b0_010011101011_001_0_101011010011;
      patterns[10074] = 29'b0_010011101011_010_0_100111010110;
      patterns[10075] = 29'b0_010011101011_011_1_001110101100;
      patterns[10076] = 29'b0_010011101011_100_1_001001110101;
      patterns[10077] = 29'b0_010011101011_101_1_100100111010;
      patterns[10078] = 29'b0_010011101011_110_0_010011101011;
      patterns[10079] = 29'b0_010011101011_111_0_010011101011;
      patterns[10080] = 29'b0_010011101100_000_0_010011101100;
      patterns[10081] = 29'b0_010011101100_001_0_101100010011;
      patterns[10082] = 29'b0_010011101100_010_0_100111011000;
      patterns[10083] = 29'b0_010011101100_011_1_001110110000;
      patterns[10084] = 29'b0_010011101100_100_0_001001110110;
      patterns[10085] = 29'b0_010011101100_101_0_000100111011;
      patterns[10086] = 29'b0_010011101100_110_0_010011101100;
      patterns[10087] = 29'b0_010011101100_111_0_010011101100;
      patterns[10088] = 29'b0_010011101101_000_0_010011101101;
      patterns[10089] = 29'b0_010011101101_001_0_101101010011;
      patterns[10090] = 29'b0_010011101101_010_0_100111011010;
      patterns[10091] = 29'b0_010011101101_011_1_001110110100;
      patterns[10092] = 29'b0_010011101101_100_1_001001110110;
      patterns[10093] = 29'b0_010011101101_101_0_100100111011;
      patterns[10094] = 29'b0_010011101101_110_0_010011101101;
      patterns[10095] = 29'b0_010011101101_111_0_010011101101;
      patterns[10096] = 29'b0_010011101110_000_0_010011101110;
      patterns[10097] = 29'b0_010011101110_001_0_101110010011;
      patterns[10098] = 29'b0_010011101110_010_0_100111011100;
      patterns[10099] = 29'b0_010011101110_011_1_001110111000;
      patterns[10100] = 29'b0_010011101110_100_0_001001110111;
      patterns[10101] = 29'b0_010011101110_101_1_000100111011;
      patterns[10102] = 29'b0_010011101110_110_0_010011101110;
      patterns[10103] = 29'b0_010011101110_111_0_010011101110;
      patterns[10104] = 29'b0_010011101111_000_0_010011101111;
      patterns[10105] = 29'b0_010011101111_001_0_101111010011;
      patterns[10106] = 29'b0_010011101111_010_0_100111011110;
      patterns[10107] = 29'b0_010011101111_011_1_001110111100;
      patterns[10108] = 29'b0_010011101111_100_1_001001110111;
      patterns[10109] = 29'b0_010011101111_101_1_100100111011;
      patterns[10110] = 29'b0_010011101111_110_0_010011101111;
      patterns[10111] = 29'b0_010011101111_111_0_010011101111;
      patterns[10112] = 29'b0_010011110000_000_0_010011110000;
      patterns[10113] = 29'b0_010011110000_001_0_110000010011;
      patterns[10114] = 29'b0_010011110000_010_0_100111100000;
      patterns[10115] = 29'b0_010011110000_011_1_001111000000;
      patterns[10116] = 29'b0_010011110000_100_0_001001111000;
      patterns[10117] = 29'b0_010011110000_101_0_000100111100;
      patterns[10118] = 29'b0_010011110000_110_0_010011110000;
      patterns[10119] = 29'b0_010011110000_111_0_010011110000;
      patterns[10120] = 29'b0_010011110001_000_0_010011110001;
      patterns[10121] = 29'b0_010011110001_001_0_110001010011;
      patterns[10122] = 29'b0_010011110001_010_0_100111100010;
      patterns[10123] = 29'b0_010011110001_011_1_001111000100;
      patterns[10124] = 29'b0_010011110001_100_1_001001111000;
      patterns[10125] = 29'b0_010011110001_101_0_100100111100;
      patterns[10126] = 29'b0_010011110001_110_0_010011110001;
      patterns[10127] = 29'b0_010011110001_111_0_010011110001;
      patterns[10128] = 29'b0_010011110010_000_0_010011110010;
      patterns[10129] = 29'b0_010011110010_001_0_110010010011;
      patterns[10130] = 29'b0_010011110010_010_0_100111100100;
      patterns[10131] = 29'b0_010011110010_011_1_001111001000;
      patterns[10132] = 29'b0_010011110010_100_0_001001111001;
      patterns[10133] = 29'b0_010011110010_101_1_000100111100;
      patterns[10134] = 29'b0_010011110010_110_0_010011110010;
      patterns[10135] = 29'b0_010011110010_111_0_010011110010;
      patterns[10136] = 29'b0_010011110011_000_0_010011110011;
      patterns[10137] = 29'b0_010011110011_001_0_110011010011;
      patterns[10138] = 29'b0_010011110011_010_0_100111100110;
      patterns[10139] = 29'b0_010011110011_011_1_001111001100;
      patterns[10140] = 29'b0_010011110011_100_1_001001111001;
      patterns[10141] = 29'b0_010011110011_101_1_100100111100;
      patterns[10142] = 29'b0_010011110011_110_0_010011110011;
      patterns[10143] = 29'b0_010011110011_111_0_010011110011;
      patterns[10144] = 29'b0_010011110100_000_0_010011110100;
      patterns[10145] = 29'b0_010011110100_001_0_110100010011;
      patterns[10146] = 29'b0_010011110100_010_0_100111101000;
      patterns[10147] = 29'b0_010011110100_011_1_001111010000;
      patterns[10148] = 29'b0_010011110100_100_0_001001111010;
      patterns[10149] = 29'b0_010011110100_101_0_000100111101;
      patterns[10150] = 29'b0_010011110100_110_0_010011110100;
      patterns[10151] = 29'b0_010011110100_111_0_010011110100;
      patterns[10152] = 29'b0_010011110101_000_0_010011110101;
      patterns[10153] = 29'b0_010011110101_001_0_110101010011;
      patterns[10154] = 29'b0_010011110101_010_0_100111101010;
      patterns[10155] = 29'b0_010011110101_011_1_001111010100;
      patterns[10156] = 29'b0_010011110101_100_1_001001111010;
      patterns[10157] = 29'b0_010011110101_101_0_100100111101;
      patterns[10158] = 29'b0_010011110101_110_0_010011110101;
      patterns[10159] = 29'b0_010011110101_111_0_010011110101;
      patterns[10160] = 29'b0_010011110110_000_0_010011110110;
      patterns[10161] = 29'b0_010011110110_001_0_110110010011;
      patterns[10162] = 29'b0_010011110110_010_0_100111101100;
      patterns[10163] = 29'b0_010011110110_011_1_001111011000;
      patterns[10164] = 29'b0_010011110110_100_0_001001111011;
      patterns[10165] = 29'b0_010011110110_101_1_000100111101;
      patterns[10166] = 29'b0_010011110110_110_0_010011110110;
      patterns[10167] = 29'b0_010011110110_111_0_010011110110;
      patterns[10168] = 29'b0_010011110111_000_0_010011110111;
      patterns[10169] = 29'b0_010011110111_001_0_110111010011;
      patterns[10170] = 29'b0_010011110111_010_0_100111101110;
      patterns[10171] = 29'b0_010011110111_011_1_001111011100;
      patterns[10172] = 29'b0_010011110111_100_1_001001111011;
      patterns[10173] = 29'b0_010011110111_101_1_100100111101;
      patterns[10174] = 29'b0_010011110111_110_0_010011110111;
      patterns[10175] = 29'b0_010011110111_111_0_010011110111;
      patterns[10176] = 29'b0_010011111000_000_0_010011111000;
      patterns[10177] = 29'b0_010011111000_001_0_111000010011;
      patterns[10178] = 29'b0_010011111000_010_0_100111110000;
      patterns[10179] = 29'b0_010011111000_011_1_001111100000;
      patterns[10180] = 29'b0_010011111000_100_0_001001111100;
      patterns[10181] = 29'b0_010011111000_101_0_000100111110;
      patterns[10182] = 29'b0_010011111000_110_0_010011111000;
      patterns[10183] = 29'b0_010011111000_111_0_010011111000;
      patterns[10184] = 29'b0_010011111001_000_0_010011111001;
      patterns[10185] = 29'b0_010011111001_001_0_111001010011;
      patterns[10186] = 29'b0_010011111001_010_0_100111110010;
      patterns[10187] = 29'b0_010011111001_011_1_001111100100;
      patterns[10188] = 29'b0_010011111001_100_1_001001111100;
      patterns[10189] = 29'b0_010011111001_101_0_100100111110;
      patterns[10190] = 29'b0_010011111001_110_0_010011111001;
      patterns[10191] = 29'b0_010011111001_111_0_010011111001;
      patterns[10192] = 29'b0_010011111010_000_0_010011111010;
      patterns[10193] = 29'b0_010011111010_001_0_111010010011;
      patterns[10194] = 29'b0_010011111010_010_0_100111110100;
      patterns[10195] = 29'b0_010011111010_011_1_001111101000;
      patterns[10196] = 29'b0_010011111010_100_0_001001111101;
      patterns[10197] = 29'b0_010011111010_101_1_000100111110;
      patterns[10198] = 29'b0_010011111010_110_0_010011111010;
      patterns[10199] = 29'b0_010011111010_111_0_010011111010;
      patterns[10200] = 29'b0_010011111011_000_0_010011111011;
      patterns[10201] = 29'b0_010011111011_001_0_111011010011;
      patterns[10202] = 29'b0_010011111011_010_0_100111110110;
      patterns[10203] = 29'b0_010011111011_011_1_001111101100;
      patterns[10204] = 29'b0_010011111011_100_1_001001111101;
      patterns[10205] = 29'b0_010011111011_101_1_100100111110;
      patterns[10206] = 29'b0_010011111011_110_0_010011111011;
      patterns[10207] = 29'b0_010011111011_111_0_010011111011;
      patterns[10208] = 29'b0_010011111100_000_0_010011111100;
      patterns[10209] = 29'b0_010011111100_001_0_111100010011;
      patterns[10210] = 29'b0_010011111100_010_0_100111111000;
      patterns[10211] = 29'b0_010011111100_011_1_001111110000;
      patterns[10212] = 29'b0_010011111100_100_0_001001111110;
      patterns[10213] = 29'b0_010011111100_101_0_000100111111;
      patterns[10214] = 29'b0_010011111100_110_0_010011111100;
      patterns[10215] = 29'b0_010011111100_111_0_010011111100;
      patterns[10216] = 29'b0_010011111101_000_0_010011111101;
      patterns[10217] = 29'b0_010011111101_001_0_111101010011;
      patterns[10218] = 29'b0_010011111101_010_0_100111111010;
      patterns[10219] = 29'b0_010011111101_011_1_001111110100;
      patterns[10220] = 29'b0_010011111101_100_1_001001111110;
      patterns[10221] = 29'b0_010011111101_101_0_100100111111;
      patterns[10222] = 29'b0_010011111101_110_0_010011111101;
      patterns[10223] = 29'b0_010011111101_111_0_010011111101;
      patterns[10224] = 29'b0_010011111110_000_0_010011111110;
      patterns[10225] = 29'b0_010011111110_001_0_111110010011;
      patterns[10226] = 29'b0_010011111110_010_0_100111111100;
      patterns[10227] = 29'b0_010011111110_011_1_001111111000;
      patterns[10228] = 29'b0_010011111110_100_0_001001111111;
      patterns[10229] = 29'b0_010011111110_101_1_000100111111;
      patterns[10230] = 29'b0_010011111110_110_0_010011111110;
      patterns[10231] = 29'b0_010011111110_111_0_010011111110;
      patterns[10232] = 29'b0_010011111111_000_0_010011111111;
      patterns[10233] = 29'b0_010011111111_001_0_111111010011;
      patterns[10234] = 29'b0_010011111111_010_0_100111111110;
      patterns[10235] = 29'b0_010011111111_011_1_001111111100;
      patterns[10236] = 29'b0_010011111111_100_1_001001111111;
      patterns[10237] = 29'b0_010011111111_101_1_100100111111;
      patterns[10238] = 29'b0_010011111111_110_0_010011111111;
      patterns[10239] = 29'b0_010011111111_111_0_010011111111;
      patterns[10240] = 29'b0_010100000000_000_0_010100000000;
      patterns[10241] = 29'b0_010100000000_001_0_000000010100;
      patterns[10242] = 29'b0_010100000000_010_0_101000000000;
      patterns[10243] = 29'b0_010100000000_011_1_010000000000;
      patterns[10244] = 29'b0_010100000000_100_0_001010000000;
      patterns[10245] = 29'b0_010100000000_101_0_000101000000;
      patterns[10246] = 29'b0_010100000000_110_0_010100000000;
      patterns[10247] = 29'b0_010100000000_111_0_010100000000;
      patterns[10248] = 29'b0_010100000001_000_0_010100000001;
      patterns[10249] = 29'b0_010100000001_001_0_000001010100;
      patterns[10250] = 29'b0_010100000001_010_0_101000000010;
      patterns[10251] = 29'b0_010100000001_011_1_010000000100;
      patterns[10252] = 29'b0_010100000001_100_1_001010000000;
      patterns[10253] = 29'b0_010100000001_101_0_100101000000;
      patterns[10254] = 29'b0_010100000001_110_0_010100000001;
      patterns[10255] = 29'b0_010100000001_111_0_010100000001;
      patterns[10256] = 29'b0_010100000010_000_0_010100000010;
      patterns[10257] = 29'b0_010100000010_001_0_000010010100;
      patterns[10258] = 29'b0_010100000010_010_0_101000000100;
      patterns[10259] = 29'b0_010100000010_011_1_010000001000;
      patterns[10260] = 29'b0_010100000010_100_0_001010000001;
      patterns[10261] = 29'b0_010100000010_101_1_000101000000;
      patterns[10262] = 29'b0_010100000010_110_0_010100000010;
      patterns[10263] = 29'b0_010100000010_111_0_010100000010;
      patterns[10264] = 29'b0_010100000011_000_0_010100000011;
      patterns[10265] = 29'b0_010100000011_001_0_000011010100;
      patterns[10266] = 29'b0_010100000011_010_0_101000000110;
      patterns[10267] = 29'b0_010100000011_011_1_010000001100;
      patterns[10268] = 29'b0_010100000011_100_1_001010000001;
      patterns[10269] = 29'b0_010100000011_101_1_100101000000;
      patterns[10270] = 29'b0_010100000011_110_0_010100000011;
      patterns[10271] = 29'b0_010100000011_111_0_010100000011;
      patterns[10272] = 29'b0_010100000100_000_0_010100000100;
      patterns[10273] = 29'b0_010100000100_001_0_000100010100;
      patterns[10274] = 29'b0_010100000100_010_0_101000001000;
      patterns[10275] = 29'b0_010100000100_011_1_010000010000;
      patterns[10276] = 29'b0_010100000100_100_0_001010000010;
      patterns[10277] = 29'b0_010100000100_101_0_000101000001;
      patterns[10278] = 29'b0_010100000100_110_0_010100000100;
      patterns[10279] = 29'b0_010100000100_111_0_010100000100;
      patterns[10280] = 29'b0_010100000101_000_0_010100000101;
      patterns[10281] = 29'b0_010100000101_001_0_000101010100;
      patterns[10282] = 29'b0_010100000101_010_0_101000001010;
      patterns[10283] = 29'b0_010100000101_011_1_010000010100;
      patterns[10284] = 29'b0_010100000101_100_1_001010000010;
      patterns[10285] = 29'b0_010100000101_101_0_100101000001;
      patterns[10286] = 29'b0_010100000101_110_0_010100000101;
      patterns[10287] = 29'b0_010100000101_111_0_010100000101;
      patterns[10288] = 29'b0_010100000110_000_0_010100000110;
      patterns[10289] = 29'b0_010100000110_001_0_000110010100;
      patterns[10290] = 29'b0_010100000110_010_0_101000001100;
      patterns[10291] = 29'b0_010100000110_011_1_010000011000;
      patterns[10292] = 29'b0_010100000110_100_0_001010000011;
      patterns[10293] = 29'b0_010100000110_101_1_000101000001;
      patterns[10294] = 29'b0_010100000110_110_0_010100000110;
      patterns[10295] = 29'b0_010100000110_111_0_010100000110;
      patterns[10296] = 29'b0_010100000111_000_0_010100000111;
      patterns[10297] = 29'b0_010100000111_001_0_000111010100;
      patterns[10298] = 29'b0_010100000111_010_0_101000001110;
      patterns[10299] = 29'b0_010100000111_011_1_010000011100;
      patterns[10300] = 29'b0_010100000111_100_1_001010000011;
      patterns[10301] = 29'b0_010100000111_101_1_100101000001;
      patterns[10302] = 29'b0_010100000111_110_0_010100000111;
      patterns[10303] = 29'b0_010100000111_111_0_010100000111;
      patterns[10304] = 29'b0_010100001000_000_0_010100001000;
      patterns[10305] = 29'b0_010100001000_001_0_001000010100;
      patterns[10306] = 29'b0_010100001000_010_0_101000010000;
      patterns[10307] = 29'b0_010100001000_011_1_010000100000;
      patterns[10308] = 29'b0_010100001000_100_0_001010000100;
      patterns[10309] = 29'b0_010100001000_101_0_000101000010;
      patterns[10310] = 29'b0_010100001000_110_0_010100001000;
      patterns[10311] = 29'b0_010100001000_111_0_010100001000;
      patterns[10312] = 29'b0_010100001001_000_0_010100001001;
      patterns[10313] = 29'b0_010100001001_001_0_001001010100;
      patterns[10314] = 29'b0_010100001001_010_0_101000010010;
      patterns[10315] = 29'b0_010100001001_011_1_010000100100;
      patterns[10316] = 29'b0_010100001001_100_1_001010000100;
      patterns[10317] = 29'b0_010100001001_101_0_100101000010;
      patterns[10318] = 29'b0_010100001001_110_0_010100001001;
      patterns[10319] = 29'b0_010100001001_111_0_010100001001;
      patterns[10320] = 29'b0_010100001010_000_0_010100001010;
      patterns[10321] = 29'b0_010100001010_001_0_001010010100;
      patterns[10322] = 29'b0_010100001010_010_0_101000010100;
      patterns[10323] = 29'b0_010100001010_011_1_010000101000;
      patterns[10324] = 29'b0_010100001010_100_0_001010000101;
      patterns[10325] = 29'b0_010100001010_101_1_000101000010;
      patterns[10326] = 29'b0_010100001010_110_0_010100001010;
      patterns[10327] = 29'b0_010100001010_111_0_010100001010;
      patterns[10328] = 29'b0_010100001011_000_0_010100001011;
      patterns[10329] = 29'b0_010100001011_001_0_001011010100;
      patterns[10330] = 29'b0_010100001011_010_0_101000010110;
      patterns[10331] = 29'b0_010100001011_011_1_010000101100;
      patterns[10332] = 29'b0_010100001011_100_1_001010000101;
      patterns[10333] = 29'b0_010100001011_101_1_100101000010;
      patterns[10334] = 29'b0_010100001011_110_0_010100001011;
      patterns[10335] = 29'b0_010100001011_111_0_010100001011;
      patterns[10336] = 29'b0_010100001100_000_0_010100001100;
      patterns[10337] = 29'b0_010100001100_001_0_001100010100;
      patterns[10338] = 29'b0_010100001100_010_0_101000011000;
      patterns[10339] = 29'b0_010100001100_011_1_010000110000;
      patterns[10340] = 29'b0_010100001100_100_0_001010000110;
      patterns[10341] = 29'b0_010100001100_101_0_000101000011;
      patterns[10342] = 29'b0_010100001100_110_0_010100001100;
      patterns[10343] = 29'b0_010100001100_111_0_010100001100;
      patterns[10344] = 29'b0_010100001101_000_0_010100001101;
      patterns[10345] = 29'b0_010100001101_001_0_001101010100;
      patterns[10346] = 29'b0_010100001101_010_0_101000011010;
      patterns[10347] = 29'b0_010100001101_011_1_010000110100;
      patterns[10348] = 29'b0_010100001101_100_1_001010000110;
      patterns[10349] = 29'b0_010100001101_101_0_100101000011;
      patterns[10350] = 29'b0_010100001101_110_0_010100001101;
      patterns[10351] = 29'b0_010100001101_111_0_010100001101;
      patterns[10352] = 29'b0_010100001110_000_0_010100001110;
      patterns[10353] = 29'b0_010100001110_001_0_001110010100;
      patterns[10354] = 29'b0_010100001110_010_0_101000011100;
      patterns[10355] = 29'b0_010100001110_011_1_010000111000;
      patterns[10356] = 29'b0_010100001110_100_0_001010000111;
      patterns[10357] = 29'b0_010100001110_101_1_000101000011;
      patterns[10358] = 29'b0_010100001110_110_0_010100001110;
      patterns[10359] = 29'b0_010100001110_111_0_010100001110;
      patterns[10360] = 29'b0_010100001111_000_0_010100001111;
      patterns[10361] = 29'b0_010100001111_001_0_001111010100;
      patterns[10362] = 29'b0_010100001111_010_0_101000011110;
      patterns[10363] = 29'b0_010100001111_011_1_010000111100;
      patterns[10364] = 29'b0_010100001111_100_1_001010000111;
      patterns[10365] = 29'b0_010100001111_101_1_100101000011;
      patterns[10366] = 29'b0_010100001111_110_0_010100001111;
      patterns[10367] = 29'b0_010100001111_111_0_010100001111;
      patterns[10368] = 29'b0_010100010000_000_0_010100010000;
      patterns[10369] = 29'b0_010100010000_001_0_010000010100;
      patterns[10370] = 29'b0_010100010000_010_0_101000100000;
      patterns[10371] = 29'b0_010100010000_011_1_010001000000;
      patterns[10372] = 29'b0_010100010000_100_0_001010001000;
      patterns[10373] = 29'b0_010100010000_101_0_000101000100;
      patterns[10374] = 29'b0_010100010000_110_0_010100010000;
      patterns[10375] = 29'b0_010100010000_111_0_010100010000;
      patterns[10376] = 29'b0_010100010001_000_0_010100010001;
      patterns[10377] = 29'b0_010100010001_001_0_010001010100;
      patterns[10378] = 29'b0_010100010001_010_0_101000100010;
      patterns[10379] = 29'b0_010100010001_011_1_010001000100;
      patterns[10380] = 29'b0_010100010001_100_1_001010001000;
      patterns[10381] = 29'b0_010100010001_101_0_100101000100;
      patterns[10382] = 29'b0_010100010001_110_0_010100010001;
      patterns[10383] = 29'b0_010100010001_111_0_010100010001;
      patterns[10384] = 29'b0_010100010010_000_0_010100010010;
      patterns[10385] = 29'b0_010100010010_001_0_010010010100;
      patterns[10386] = 29'b0_010100010010_010_0_101000100100;
      patterns[10387] = 29'b0_010100010010_011_1_010001001000;
      patterns[10388] = 29'b0_010100010010_100_0_001010001001;
      patterns[10389] = 29'b0_010100010010_101_1_000101000100;
      patterns[10390] = 29'b0_010100010010_110_0_010100010010;
      patterns[10391] = 29'b0_010100010010_111_0_010100010010;
      patterns[10392] = 29'b0_010100010011_000_0_010100010011;
      patterns[10393] = 29'b0_010100010011_001_0_010011010100;
      patterns[10394] = 29'b0_010100010011_010_0_101000100110;
      patterns[10395] = 29'b0_010100010011_011_1_010001001100;
      patterns[10396] = 29'b0_010100010011_100_1_001010001001;
      patterns[10397] = 29'b0_010100010011_101_1_100101000100;
      patterns[10398] = 29'b0_010100010011_110_0_010100010011;
      patterns[10399] = 29'b0_010100010011_111_0_010100010011;
      patterns[10400] = 29'b0_010100010100_000_0_010100010100;
      patterns[10401] = 29'b0_010100010100_001_0_010100010100;
      patterns[10402] = 29'b0_010100010100_010_0_101000101000;
      patterns[10403] = 29'b0_010100010100_011_1_010001010000;
      patterns[10404] = 29'b0_010100010100_100_0_001010001010;
      patterns[10405] = 29'b0_010100010100_101_0_000101000101;
      patterns[10406] = 29'b0_010100010100_110_0_010100010100;
      patterns[10407] = 29'b0_010100010100_111_0_010100010100;
      patterns[10408] = 29'b0_010100010101_000_0_010100010101;
      patterns[10409] = 29'b0_010100010101_001_0_010101010100;
      patterns[10410] = 29'b0_010100010101_010_0_101000101010;
      patterns[10411] = 29'b0_010100010101_011_1_010001010100;
      patterns[10412] = 29'b0_010100010101_100_1_001010001010;
      patterns[10413] = 29'b0_010100010101_101_0_100101000101;
      patterns[10414] = 29'b0_010100010101_110_0_010100010101;
      patterns[10415] = 29'b0_010100010101_111_0_010100010101;
      patterns[10416] = 29'b0_010100010110_000_0_010100010110;
      patterns[10417] = 29'b0_010100010110_001_0_010110010100;
      patterns[10418] = 29'b0_010100010110_010_0_101000101100;
      patterns[10419] = 29'b0_010100010110_011_1_010001011000;
      patterns[10420] = 29'b0_010100010110_100_0_001010001011;
      patterns[10421] = 29'b0_010100010110_101_1_000101000101;
      patterns[10422] = 29'b0_010100010110_110_0_010100010110;
      patterns[10423] = 29'b0_010100010110_111_0_010100010110;
      patterns[10424] = 29'b0_010100010111_000_0_010100010111;
      patterns[10425] = 29'b0_010100010111_001_0_010111010100;
      patterns[10426] = 29'b0_010100010111_010_0_101000101110;
      patterns[10427] = 29'b0_010100010111_011_1_010001011100;
      patterns[10428] = 29'b0_010100010111_100_1_001010001011;
      patterns[10429] = 29'b0_010100010111_101_1_100101000101;
      patterns[10430] = 29'b0_010100010111_110_0_010100010111;
      patterns[10431] = 29'b0_010100010111_111_0_010100010111;
      patterns[10432] = 29'b0_010100011000_000_0_010100011000;
      patterns[10433] = 29'b0_010100011000_001_0_011000010100;
      patterns[10434] = 29'b0_010100011000_010_0_101000110000;
      patterns[10435] = 29'b0_010100011000_011_1_010001100000;
      patterns[10436] = 29'b0_010100011000_100_0_001010001100;
      patterns[10437] = 29'b0_010100011000_101_0_000101000110;
      patterns[10438] = 29'b0_010100011000_110_0_010100011000;
      patterns[10439] = 29'b0_010100011000_111_0_010100011000;
      patterns[10440] = 29'b0_010100011001_000_0_010100011001;
      patterns[10441] = 29'b0_010100011001_001_0_011001010100;
      patterns[10442] = 29'b0_010100011001_010_0_101000110010;
      patterns[10443] = 29'b0_010100011001_011_1_010001100100;
      patterns[10444] = 29'b0_010100011001_100_1_001010001100;
      patterns[10445] = 29'b0_010100011001_101_0_100101000110;
      patterns[10446] = 29'b0_010100011001_110_0_010100011001;
      patterns[10447] = 29'b0_010100011001_111_0_010100011001;
      patterns[10448] = 29'b0_010100011010_000_0_010100011010;
      patterns[10449] = 29'b0_010100011010_001_0_011010010100;
      patterns[10450] = 29'b0_010100011010_010_0_101000110100;
      patterns[10451] = 29'b0_010100011010_011_1_010001101000;
      patterns[10452] = 29'b0_010100011010_100_0_001010001101;
      patterns[10453] = 29'b0_010100011010_101_1_000101000110;
      patterns[10454] = 29'b0_010100011010_110_0_010100011010;
      patterns[10455] = 29'b0_010100011010_111_0_010100011010;
      patterns[10456] = 29'b0_010100011011_000_0_010100011011;
      patterns[10457] = 29'b0_010100011011_001_0_011011010100;
      patterns[10458] = 29'b0_010100011011_010_0_101000110110;
      patterns[10459] = 29'b0_010100011011_011_1_010001101100;
      patterns[10460] = 29'b0_010100011011_100_1_001010001101;
      patterns[10461] = 29'b0_010100011011_101_1_100101000110;
      patterns[10462] = 29'b0_010100011011_110_0_010100011011;
      patterns[10463] = 29'b0_010100011011_111_0_010100011011;
      patterns[10464] = 29'b0_010100011100_000_0_010100011100;
      patterns[10465] = 29'b0_010100011100_001_0_011100010100;
      patterns[10466] = 29'b0_010100011100_010_0_101000111000;
      patterns[10467] = 29'b0_010100011100_011_1_010001110000;
      patterns[10468] = 29'b0_010100011100_100_0_001010001110;
      patterns[10469] = 29'b0_010100011100_101_0_000101000111;
      patterns[10470] = 29'b0_010100011100_110_0_010100011100;
      patterns[10471] = 29'b0_010100011100_111_0_010100011100;
      patterns[10472] = 29'b0_010100011101_000_0_010100011101;
      patterns[10473] = 29'b0_010100011101_001_0_011101010100;
      patterns[10474] = 29'b0_010100011101_010_0_101000111010;
      patterns[10475] = 29'b0_010100011101_011_1_010001110100;
      patterns[10476] = 29'b0_010100011101_100_1_001010001110;
      patterns[10477] = 29'b0_010100011101_101_0_100101000111;
      patterns[10478] = 29'b0_010100011101_110_0_010100011101;
      patterns[10479] = 29'b0_010100011101_111_0_010100011101;
      patterns[10480] = 29'b0_010100011110_000_0_010100011110;
      patterns[10481] = 29'b0_010100011110_001_0_011110010100;
      patterns[10482] = 29'b0_010100011110_010_0_101000111100;
      patterns[10483] = 29'b0_010100011110_011_1_010001111000;
      patterns[10484] = 29'b0_010100011110_100_0_001010001111;
      patterns[10485] = 29'b0_010100011110_101_1_000101000111;
      patterns[10486] = 29'b0_010100011110_110_0_010100011110;
      patterns[10487] = 29'b0_010100011110_111_0_010100011110;
      patterns[10488] = 29'b0_010100011111_000_0_010100011111;
      patterns[10489] = 29'b0_010100011111_001_0_011111010100;
      patterns[10490] = 29'b0_010100011111_010_0_101000111110;
      patterns[10491] = 29'b0_010100011111_011_1_010001111100;
      patterns[10492] = 29'b0_010100011111_100_1_001010001111;
      patterns[10493] = 29'b0_010100011111_101_1_100101000111;
      patterns[10494] = 29'b0_010100011111_110_0_010100011111;
      patterns[10495] = 29'b0_010100011111_111_0_010100011111;
      patterns[10496] = 29'b0_010100100000_000_0_010100100000;
      patterns[10497] = 29'b0_010100100000_001_0_100000010100;
      patterns[10498] = 29'b0_010100100000_010_0_101001000000;
      patterns[10499] = 29'b0_010100100000_011_1_010010000000;
      patterns[10500] = 29'b0_010100100000_100_0_001010010000;
      patterns[10501] = 29'b0_010100100000_101_0_000101001000;
      patterns[10502] = 29'b0_010100100000_110_0_010100100000;
      patterns[10503] = 29'b0_010100100000_111_0_010100100000;
      patterns[10504] = 29'b0_010100100001_000_0_010100100001;
      patterns[10505] = 29'b0_010100100001_001_0_100001010100;
      patterns[10506] = 29'b0_010100100001_010_0_101001000010;
      patterns[10507] = 29'b0_010100100001_011_1_010010000100;
      patterns[10508] = 29'b0_010100100001_100_1_001010010000;
      patterns[10509] = 29'b0_010100100001_101_0_100101001000;
      patterns[10510] = 29'b0_010100100001_110_0_010100100001;
      patterns[10511] = 29'b0_010100100001_111_0_010100100001;
      patterns[10512] = 29'b0_010100100010_000_0_010100100010;
      patterns[10513] = 29'b0_010100100010_001_0_100010010100;
      patterns[10514] = 29'b0_010100100010_010_0_101001000100;
      patterns[10515] = 29'b0_010100100010_011_1_010010001000;
      patterns[10516] = 29'b0_010100100010_100_0_001010010001;
      patterns[10517] = 29'b0_010100100010_101_1_000101001000;
      patterns[10518] = 29'b0_010100100010_110_0_010100100010;
      patterns[10519] = 29'b0_010100100010_111_0_010100100010;
      patterns[10520] = 29'b0_010100100011_000_0_010100100011;
      patterns[10521] = 29'b0_010100100011_001_0_100011010100;
      patterns[10522] = 29'b0_010100100011_010_0_101001000110;
      patterns[10523] = 29'b0_010100100011_011_1_010010001100;
      patterns[10524] = 29'b0_010100100011_100_1_001010010001;
      patterns[10525] = 29'b0_010100100011_101_1_100101001000;
      patterns[10526] = 29'b0_010100100011_110_0_010100100011;
      patterns[10527] = 29'b0_010100100011_111_0_010100100011;
      patterns[10528] = 29'b0_010100100100_000_0_010100100100;
      patterns[10529] = 29'b0_010100100100_001_0_100100010100;
      patterns[10530] = 29'b0_010100100100_010_0_101001001000;
      patterns[10531] = 29'b0_010100100100_011_1_010010010000;
      patterns[10532] = 29'b0_010100100100_100_0_001010010010;
      patterns[10533] = 29'b0_010100100100_101_0_000101001001;
      patterns[10534] = 29'b0_010100100100_110_0_010100100100;
      patterns[10535] = 29'b0_010100100100_111_0_010100100100;
      patterns[10536] = 29'b0_010100100101_000_0_010100100101;
      patterns[10537] = 29'b0_010100100101_001_0_100101010100;
      patterns[10538] = 29'b0_010100100101_010_0_101001001010;
      patterns[10539] = 29'b0_010100100101_011_1_010010010100;
      patterns[10540] = 29'b0_010100100101_100_1_001010010010;
      patterns[10541] = 29'b0_010100100101_101_0_100101001001;
      patterns[10542] = 29'b0_010100100101_110_0_010100100101;
      patterns[10543] = 29'b0_010100100101_111_0_010100100101;
      patterns[10544] = 29'b0_010100100110_000_0_010100100110;
      patterns[10545] = 29'b0_010100100110_001_0_100110010100;
      patterns[10546] = 29'b0_010100100110_010_0_101001001100;
      patterns[10547] = 29'b0_010100100110_011_1_010010011000;
      patterns[10548] = 29'b0_010100100110_100_0_001010010011;
      patterns[10549] = 29'b0_010100100110_101_1_000101001001;
      patterns[10550] = 29'b0_010100100110_110_0_010100100110;
      patterns[10551] = 29'b0_010100100110_111_0_010100100110;
      patterns[10552] = 29'b0_010100100111_000_0_010100100111;
      patterns[10553] = 29'b0_010100100111_001_0_100111010100;
      patterns[10554] = 29'b0_010100100111_010_0_101001001110;
      patterns[10555] = 29'b0_010100100111_011_1_010010011100;
      patterns[10556] = 29'b0_010100100111_100_1_001010010011;
      patterns[10557] = 29'b0_010100100111_101_1_100101001001;
      patterns[10558] = 29'b0_010100100111_110_0_010100100111;
      patterns[10559] = 29'b0_010100100111_111_0_010100100111;
      patterns[10560] = 29'b0_010100101000_000_0_010100101000;
      patterns[10561] = 29'b0_010100101000_001_0_101000010100;
      patterns[10562] = 29'b0_010100101000_010_0_101001010000;
      patterns[10563] = 29'b0_010100101000_011_1_010010100000;
      patterns[10564] = 29'b0_010100101000_100_0_001010010100;
      patterns[10565] = 29'b0_010100101000_101_0_000101001010;
      patterns[10566] = 29'b0_010100101000_110_0_010100101000;
      patterns[10567] = 29'b0_010100101000_111_0_010100101000;
      patterns[10568] = 29'b0_010100101001_000_0_010100101001;
      patterns[10569] = 29'b0_010100101001_001_0_101001010100;
      patterns[10570] = 29'b0_010100101001_010_0_101001010010;
      patterns[10571] = 29'b0_010100101001_011_1_010010100100;
      patterns[10572] = 29'b0_010100101001_100_1_001010010100;
      patterns[10573] = 29'b0_010100101001_101_0_100101001010;
      patterns[10574] = 29'b0_010100101001_110_0_010100101001;
      patterns[10575] = 29'b0_010100101001_111_0_010100101001;
      patterns[10576] = 29'b0_010100101010_000_0_010100101010;
      patterns[10577] = 29'b0_010100101010_001_0_101010010100;
      patterns[10578] = 29'b0_010100101010_010_0_101001010100;
      patterns[10579] = 29'b0_010100101010_011_1_010010101000;
      patterns[10580] = 29'b0_010100101010_100_0_001010010101;
      patterns[10581] = 29'b0_010100101010_101_1_000101001010;
      patterns[10582] = 29'b0_010100101010_110_0_010100101010;
      patterns[10583] = 29'b0_010100101010_111_0_010100101010;
      patterns[10584] = 29'b0_010100101011_000_0_010100101011;
      patterns[10585] = 29'b0_010100101011_001_0_101011010100;
      patterns[10586] = 29'b0_010100101011_010_0_101001010110;
      patterns[10587] = 29'b0_010100101011_011_1_010010101100;
      patterns[10588] = 29'b0_010100101011_100_1_001010010101;
      patterns[10589] = 29'b0_010100101011_101_1_100101001010;
      patterns[10590] = 29'b0_010100101011_110_0_010100101011;
      patterns[10591] = 29'b0_010100101011_111_0_010100101011;
      patterns[10592] = 29'b0_010100101100_000_0_010100101100;
      patterns[10593] = 29'b0_010100101100_001_0_101100010100;
      patterns[10594] = 29'b0_010100101100_010_0_101001011000;
      patterns[10595] = 29'b0_010100101100_011_1_010010110000;
      patterns[10596] = 29'b0_010100101100_100_0_001010010110;
      patterns[10597] = 29'b0_010100101100_101_0_000101001011;
      patterns[10598] = 29'b0_010100101100_110_0_010100101100;
      patterns[10599] = 29'b0_010100101100_111_0_010100101100;
      patterns[10600] = 29'b0_010100101101_000_0_010100101101;
      patterns[10601] = 29'b0_010100101101_001_0_101101010100;
      patterns[10602] = 29'b0_010100101101_010_0_101001011010;
      patterns[10603] = 29'b0_010100101101_011_1_010010110100;
      patterns[10604] = 29'b0_010100101101_100_1_001010010110;
      patterns[10605] = 29'b0_010100101101_101_0_100101001011;
      patterns[10606] = 29'b0_010100101101_110_0_010100101101;
      patterns[10607] = 29'b0_010100101101_111_0_010100101101;
      patterns[10608] = 29'b0_010100101110_000_0_010100101110;
      patterns[10609] = 29'b0_010100101110_001_0_101110010100;
      patterns[10610] = 29'b0_010100101110_010_0_101001011100;
      patterns[10611] = 29'b0_010100101110_011_1_010010111000;
      patterns[10612] = 29'b0_010100101110_100_0_001010010111;
      patterns[10613] = 29'b0_010100101110_101_1_000101001011;
      patterns[10614] = 29'b0_010100101110_110_0_010100101110;
      patterns[10615] = 29'b0_010100101110_111_0_010100101110;
      patterns[10616] = 29'b0_010100101111_000_0_010100101111;
      patterns[10617] = 29'b0_010100101111_001_0_101111010100;
      patterns[10618] = 29'b0_010100101111_010_0_101001011110;
      patterns[10619] = 29'b0_010100101111_011_1_010010111100;
      patterns[10620] = 29'b0_010100101111_100_1_001010010111;
      patterns[10621] = 29'b0_010100101111_101_1_100101001011;
      patterns[10622] = 29'b0_010100101111_110_0_010100101111;
      patterns[10623] = 29'b0_010100101111_111_0_010100101111;
      patterns[10624] = 29'b0_010100110000_000_0_010100110000;
      patterns[10625] = 29'b0_010100110000_001_0_110000010100;
      patterns[10626] = 29'b0_010100110000_010_0_101001100000;
      patterns[10627] = 29'b0_010100110000_011_1_010011000000;
      patterns[10628] = 29'b0_010100110000_100_0_001010011000;
      patterns[10629] = 29'b0_010100110000_101_0_000101001100;
      patterns[10630] = 29'b0_010100110000_110_0_010100110000;
      patterns[10631] = 29'b0_010100110000_111_0_010100110000;
      patterns[10632] = 29'b0_010100110001_000_0_010100110001;
      patterns[10633] = 29'b0_010100110001_001_0_110001010100;
      patterns[10634] = 29'b0_010100110001_010_0_101001100010;
      patterns[10635] = 29'b0_010100110001_011_1_010011000100;
      patterns[10636] = 29'b0_010100110001_100_1_001010011000;
      patterns[10637] = 29'b0_010100110001_101_0_100101001100;
      patterns[10638] = 29'b0_010100110001_110_0_010100110001;
      patterns[10639] = 29'b0_010100110001_111_0_010100110001;
      patterns[10640] = 29'b0_010100110010_000_0_010100110010;
      patterns[10641] = 29'b0_010100110010_001_0_110010010100;
      patterns[10642] = 29'b0_010100110010_010_0_101001100100;
      patterns[10643] = 29'b0_010100110010_011_1_010011001000;
      patterns[10644] = 29'b0_010100110010_100_0_001010011001;
      patterns[10645] = 29'b0_010100110010_101_1_000101001100;
      patterns[10646] = 29'b0_010100110010_110_0_010100110010;
      patterns[10647] = 29'b0_010100110010_111_0_010100110010;
      patterns[10648] = 29'b0_010100110011_000_0_010100110011;
      patterns[10649] = 29'b0_010100110011_001_0_110011010100;
      patterns[10650] = 29'b0_010100110011_010_0_101001100110;
      patterns[10651] = 29'b0_010100110011_011_1_010011001100;
      patterns[10652] = 29'b0_010100110011_100_1_001010011001;
      patterns[10653] = 29'b0_010100110011_101_1_100101001100;
      patterns[10654] = 29'b0_010100110011_110_0_010100110011;
      patterns[10655] = 29'b0_010100110011_111_0_010100110011;
      patterns[10656] = 29'b0_010100110100_000_0_010100110100;
      patterns[10657] = 29'b0_010100110100_001_0_110100010100;
      patterns[10658] = 29'b0_010100110100_010_0_101001101000;
      patterns[10659] = 29'b0_010100110100_011_1_010011010000;
      patterns[10660] = 29'b0_010100110100_100_0_001010011010;
      patterns[10661] = 29'b0_010100110100_101_0_000101001101;
      patterns[10662] = 29'b0_010100110100_110_0_010100110100;
      patterns[10663] = 29'b0_010100110100_111_0_010100110100;
      patterns[10664] = 29'b0_010100110101_000_0_010100110101;
      patterns[10665] = 29'b0_010100110101_001_0_110101010100;
      patterns[10666] = 29'b0_010100110101_010_0_101001101010;
      patterns[10667] = 29'b0_010100110101_011_1_010011010100;
      patterns[10668] = 29'b0_010100110101_100_1_001010011010;
      patterns[10669] = 29'b0_010100110101_101_0_100101001101;
      patterns[10670] = 29'b0_010100110101_110_0_010100110101;
      patterns[10671] = 29'b0_010100110101_111_0_010100110101;
      patterns[10672] = 29'b0_010100110110_000_0_010100110110;
      patterns[10673] = 29'b0_010100110110_001_0_110110010100;
      patterns[10674] = 29'b0_010100110110_010_0_101001101100;
      patterns[10675] = 29'b0_010100110110_011_1_010011011000;
      patterns[10676] = 29'b0_010100110110_100_0_001010011011;
      patterns[10677] = 29'b0_010100110110_101_1_000101001101;
      patterns[10678] = 29'b0_010100110110_110_0_010100110110;
      patterns[10679] = 29'b0_010100110110_111_0_010100110110;
      patterns[10680] = 29'b0_010100110111_000_0_010100110111;
      patterns[10681] = 29'b0_010100110111_001_0_110111010100;
      patterns[10682] = 29'b0_010100110111_010_0_101001101110;
      patterns[10683] = 29'b0_010100110111_011_1_010011011100;
      patterns[10684] = 29'b0_010100110111_100_1_001010011011;
      patterns[10685] = 29'b0_010100110111_101_1_100101001101;
      patterns[10686] = 29'b0_010100110111_110_0_010100110111;
      patterns[10687] = 29'b0_010100110111_111_0_010100110111;
      patterns[10688] = 29'b0_010100111000_000_0_010100111000;
      patterns[10689] = 29'b0_010100111000_001_0_111000010100;
      patterns[10690] = 29'b0_010100111000_010_0_101001110000;
      patterns[10691] = 29'b0_010100111000_011_1_010011100000;
      patterns[10692] = 29'b0_010100111000_100_0_001010011100;
      patterns[10693] = 29'b0_010100111000_101_0_000101001110;
      patterns[10694] = 29'b0_010100111000_110_0_010100111000;
      patterns[10695] = 29'b0_010100111000_111_0_010100111000;
      patterns[10696] = 29'b0_010100111001_000_0_010100111001;
      patterns[10697] = 29'b0_010100111001_001_0_111001010100;
      patterns[10698] = 29'b0_010100111001_010_0_101001110010;
      patterns[10699] = 29'b0_010100111001_011_1_010011100100;
      patterns[10700] = 29'b0_010100111001_100_1_001010011100;
      patterns[10701] = 29'b0_010100111001_101_0_100101001110;
      patterns[10702] = 29'b0_010100111001_110_0_010100111001;
      patterns[10703] = 29'b0_010100111001_111_0_010100111001;
      patterns[10704] = 29'b0_010100111010_000_0_010100111010;
      patterns[10705] = 29'b0_010100111010_001_0_111010010100;
      patterns[10706] = 29'b0_010100111010_010_0_101001110100;
      patterns[10707] = 29'b0_010100111010_011_1_010011101000;
      patterns[10708] = 29'b0_010100111010_100_0_001010011101;
      patterns[10709] = 29'b0_010100111010_101_1_000101001110;
      patterns[10710] = 29'b0_010100111010_110_0_010100111010;
      patterns[10711] = 29'b0_010100111010_111_0_010100111010;
      patterns[10712] = 29'b0_010100111011_000_0_010100111011;
      patterns[10713] = 29'b0_010100111011_001_0_111011010100;
      patterns[10714] = 29'b0_010100111011_010_0_101001110110;
      patterns[10715] = 29'b0_010100111011_011_1_010011101100;
      patterns[10716] = 29'b0_010100111011_100_1_001010011101;
      patterns[10717] = 29'b0_010100111011_101_1_100101001110;
      patterns[10718] = 29'b0_010100111011_110_0_010100111011;
      patterns[10719] = 29'b0_010100111011_111_0_010100111011;
      patterns[10720] = 29'b0_010100111100_000_0_010100111100;
      patterns[10721] = 29'b0_010100111100_001_0_111100010100;
      patterns[10722] = 29'b0_010100111100_010_0_101001111000;
      patterns[10723] = 29'b0_010100111100_011_1_010011110000;
      patterns[10724] = 29'b0_010100111100_100_0_001010011110;
      patterns[10725] = 29'b0_010100111100_101_0_000101001111;
      patterns[10726] = 29'b0_010100111100_110_0_010100111100;
      patterns[10727] = 29'b0_010100111100_111_0_010100111100;
      patterns[10728] = 29'b0_010100111101_000_0_010100111101;
      patterns[10729] = 29'b0_010100111101_001_0_111101010100;
      patterns[10730] = 29'b0_010100111101_010_0_101001111010;
      patterns[10731] = 29'b0_010100111101_011_1_010011110100;
      patterns[10732] = 29'b0_010100111101_100_1_001010011110;
      patterns[10733] = 29'b0_010100111101_101_0_100101001111;
      patterns[10734] = 29'b0_010100111101_110_0_010100111101;
      patterns[10735] = 29'b0_010100111101_111_0_010100111101;
      patterns[10736] = 29'b0_010100111110_000_0_010100111110;
      patterns[10737] = 29'b0_010100111110_001_0_111110010100;
      patterns[10738] = 29'b0_010100111110_010_0_101001111100;
      patterns[10739] = 29'b0_010100111110_011_1_010011111000;
      patterns[10740] = 29'b0_010100111110_100_0_001010011111;
      patterns[10741] = 29'b0_010100111110_101_1_000101001111;
      patterns[10742] = 29'b0_010100111110_110_0_010100111110;
      patterns[10743] = 29'b0_010100111110_111_0_010100111110;
      patterns[10744] = 29'b0_010100111111_000_0_010100111111;
      patterns[10745] = 29'b0_010100111111_001_0_111111010100;
      patterns[10746] = 29'b0_010100111111_010_0_101001111110;
      patterns[10747] = 29'b0_010100111111_011_1_010011111100;
      patterns[10748] = 29'b0_010100111111_100_1_001010011111;
      patterns[10749] = 29'b0_010100111111_101_1_100101001111;
      patterns[10750] = 29'b0_010100111111_110_0_010100111111;
      patterns[10751] = 29'b0_010100111111_111_0_010100111111;
      patterns[10752] = 29'b0_010101000000_000_0_010101000000;
      patterns[10753] = 29'b0_010101000000_001_0_000000010101;
      patterns[10754] = 29'b0_010101000000_010_0_101010000000;
      patterns[10755] = 29'b0_010101000000_011_1_010100000000;
      patterns[10756] = 29'b0_010101000000_100_0_001010100000;
      patterns[10757] = 29'b0_010101000000_101_0_000101010000;
      patterns[10758] = 29'b0_010101000000_110_0_010101000000;
      patterns[10759] = 29'b0_010101000000_111_0_010101000000;
      patterns[10760] = 29'b0_010101000001_000_0_010101000001;
      patterns[10761] = 29'b0_010101000001_001_0_000001010101;
      patterns[10762] = 29'b0_010101000001_010_0_101010000010;
      patterns[10763] = 29'b0_010101000001_011_1_010100000100;
      patterns[10764] = 29'b0_010101000001_100_1_001010100000;
      patterns[10765] = 29'b0_010101000001_101_0_100101010000;
      patterns[10766] = 29'b0_010101000001_110_0_010101000001;
      patterns[10767] = 29'b0_010101000001_111_0_010101000001;
      patterns[10768] = 29'b0_010101000010_000_0_010101000010;
      patterns[10769] = 29'b0_010101000010_001_0_000010010101;
      patterns[10770] = 29'b0_010101000010_010_0_101010000100;
      patterns[10771] = 29'b0_010101000010_011_1_010100001000;
      patterns[10772] = 29'b0_010101000010_100_0_001010100001;
      patterns[10773] = 29'b0_010101000010_101_1_000101010000;
      patterns[10774] = 29'b0_010101000010_110_0_010101000010;
      patterns[10775] = 29'b0_010101000010_111_0_010101000010;
      patterns[10776] = 29'b0_010101000011_000_0_010101000011;
      patterns[10777] = 29'b0_010101000011_001_0_000011010101;
      patterns[10778] = 29'b0_010101000011_010_0_101010000110;
      patterns[10779] = 29'b0_010101000011_011_1_010100001100;
      patterns[10780] = 29'b0_010101000011_100_1_001010100001;
      patterns[10781] = 29'b0_010101000011_101_1_100101010000;
      patterns[10782] = 29'b0_010101000011_110_0_010101000011;
      patterns[10783] = 29'b0_010101000011_111_0_010101000011;
      patterns[10784] = 29'b0_010101000100_000_0_010101000100;
      patterns[10785] = 29'b0_010101000100_001_0_000100010101;
      patterns[10786] = 29'b0_010101000100_010_0_101010001000;
      patterns[10787] = 29'b0_010101000100_011_1_010100010000;
      patterns[10788] = 29'b0_010101000100_100_0_001010100010;
      patterns[10789] = 29'b0_010101000100_101_0_000101010001;
      patterns[10790] = 29'b0_010101000100_110_0_010101000100;
      patterns[10791] = 29'b0_010101000100_111_0_010101000100;
      patterns[10792] = 29'b0_010101000101_000_0_010101000101;
      patterns[10793] = 29'b0_010101000101_001_0_000101010101;
      patterns[10794] = 29'b0_010101000101_010_0_101010001010;
      patterns[10795] = 29'b0_010101000101_011_1_010100010100;
      patterns[10796] = 29'b0_010101000101_100_1_001010100010;
      patterns[10797] = 29'b0_010101000101_101_0_100101010001;
      patterns[10798] = 29'b0_010101000101_110_0_010101000101;
      patterns[10799] = 29'b0_010101000101_111_0_010101000101;
      patterns[10800] = 29'b0_010101000110_000_0_010101000110;
      patterns[10801] = 29'b0_010101000110_001_0_000110010101;
      patterns[10802] = 29'b0_010101000110_010_0_101010001100;
      patterns[10803] = 29'b0_010101000110_011_1_010100011000;
      patterns[10804] = 29'b0_010101000110_100_0_001010100011;
      patterns[10805] = 29'b0_010101000110_101_1_000101010001;
      patterns[10806] = 29'b0_010101000110_110_0_010101000110;
      patterns[10807] = 29'b0_010101000110_111_0_010101000110;
      patterns[10808] = 29'b0_010101000111_000_0_010101000111;
      patterns[10809] = 29'b0_010101000111_001_0_000111010101;
      patterns[10810] = 29'b0_010101000111_010_0_101010001110;
      patterns[10811] = 29'b0_010101000111_011_1_010100011100;
      patterns[10812] = 29'b0_010101000111_100_1_001010100011;
      patterns[10813] = 29'b0_010101000111_101_1_100101010001;
      patterns[10814] = 29'b0_010101000111_110_0_010101000111;
      patterns[10815] = 29'b0_010101000111_111_0_010101000111;
      patterns[10816] = 29'b0_010101001000_000_0_010101001000;
      patterns[10817] = 29'b0_010101001000_001_0_001000010101;
      patterns[10818] = 29'b0_010101001000_010_0_101010010000;
      patterns[10819] = 29'b0_010101001000_011_1_010100100000;
      patterns[10820] = 29'b0_010101001000_100_0_001010100100;
      patterns[10821] = 29'b0_010101001000_101_0_000101010010;
      patterns[10822] = 29'b0_010101001000_110_0_010101001000;
      patterns[10823] = 29'b0_010101001000_111_0_010101001000;
      patterns[10824] = 29'b0_010101001001_000_0_010101001001;
      patterns[10825] = 29'b0_010101001001_001_0_001001010101;
      patterns[10826] = 29'b0_010101001001_010_0_101010010010;
      patterns[10827] = 29'b0_010101001001_011_1_010100100100;
      patterns[10828] = 29'b0_010101001001_100_1_001010100100;
      patterns[10829] = 29'b0_010101001001_101_0_100101010010;
      patterns[10830] = 29'b0_010101001001_110_0_010101001001;
      patterns[10831] = 29'b0_010101001001_111_0_010101001001;
      patterns[10832] = 29'b0_010101001010_000_0_010101001010;
      patterns[10833] = 29'b0_010101001010_001_0_001010010101;
      patterns[10834] = 29'b0_010101001010_010_0_101010010100;
      patterns[10835] = 29'b0_010101001010_011_1_010100101000;
      patterns[10836] = 29'b0_010101001010_100_0_001010100101;
      patterns[10837] = 29'b0_010101001010_101_1_000101010010;
      patterns[10838] = 29'b0_010101001010_110_0_010101001010;
      patterns[10839] = 29'b0_010101001010_111_0_010101001010;
      patterns[10840] = 29'b0_010101001011_000_0_010101001011;
      patterns[10841] = 29'b0_010101001011_001_0_001011010101;
      patterns[10842] = 29'b0_010101001011_010_0_101010010110;
      patterns[10843] = 29'b0_010101001011_011_1_010100101100;
      patterns[10844] = 29'b0_010101001011_100_1_001010100101;
      patterns[10845] = 29'b0_010101001011_101_1_100101010010;
      patterns[10846] = 29'b0_010101001011_110_0_010101001011;
      patterns[10847] = 29'b0_010101001011_111_0_010101001011;
      patterns[10848] = 29'b0_010101001100_000_0_010101001100;
      patterns[10849] = 29'b0_010101001100_001_0_001100010101;
      patterns[10850] = 29'b0_010101001100_010_0_101010011000;
      patterns[10851] = 29'b0_010101001100_011_1_010100110000;
      patterns[10852] = 29'b0_010101001100_100_0_001010100110;
      patterns[10853] = 29'b0_010101001100_101_0_000101010011;
      patterns[10854] = 29'b0_010101001100_110_0_010101001100;
      patterns[10855] = 29'b0_010101001100_111_0_010101001100;
      patterns[10856] = 29'b0_010101001101_000_0_010101001101;
      patterns[10857] = 29'b0_010101001101_001_0_001101010101;
      patterns[10858] = 29'b0_010101001101_010_0_101010011010;
      patterns[10859] = 29'b0_010101001101_011_1_010100110100;
      patterns[10860] = 29'b0_010101001101_100_1_001010100110;
      patterns[10861] = 29'b0_010101001101_101_0_100101010011;
      patterns[10862] = 29'b0_010101001101_110_0_010101001101;
      patterns[10863] = 29'b0_010101001101_111_0_010101001101;
      patterns[10864] = 29'b0_010101001110_000_0_010101001110;
      patterns[10865] = 29'b0_010101001110_001_0_001110010101;
      patterns[10866] = 29'b0_010101001110_010_0_101010011100;
      patterns[10867] = 29'b0_010101001110_011_1_010100111000;
      patterns[10868] = 29'b0_010101001110_100_0_001010100111;
      patterns[10869] = 29'b0_010101001110_101_1_000101010011;
      patterns[10870] = 29'b0_010101001110_110_0_010101001110;
      patterns[10871] = 29'b0_010101001110_111_0_010101001110;
      patterns[10872] = 29'b0_010101001111_000_0_010101001111;
      patterns[10873] = 29'b0_010101001111_001_0_001111010101;
      patterns[10874] = 29'b0_010101001111_010_0_101010011110;
      patterns[10875] = 29'b0_010101001111_011_1_010100111100;
      patterns[10876] = 29'b0_010101001111_100_1_001010100111;
      patterns[10877] = 29'b0_010101001111_101_1_100101010011;
      patterns[10878] = 29'b0_010101001111_110_0_010101001111;
      patterns[10879] = 29'b0_010101001111_111_0_010101001111;
      patterns[10880] = 29'b0_010101010000_000_0_010101010000;
      patterns[10881] = 29'b0_010101010000_001_0_010000010101;
      patterns[10882] = 29'b0_010101010000_010_0_101010100000;
      patterns[10883] = 29'b0_010101010000_011_1_010101000000;
      patterns[10884] = 29'b0_010101010000_100_0_001010101000;
      patterns[10885] = 29'b0_010101010000_101_0_000101010100;
      patterns[10886] = 29'b0_010101010000_110_0_010101010000;
      patterns[10887] = 29'b0_010101010000_111_0_010101010000;
      patterns[10888] = 29'b0_010101010001_000_0_010101010001;
      patterns[10889] = 29'b0_010101010001_001_0_010001010101;
      patterns[10890] = 29'b0_010101010001_010_0_101010100010;
      patterns[10891] = 29'b0_010101010001_011_1_010101000100;
      patterns[10892] = 29'b0_010101010001_100_1_001010101000;
      patterns[10893] = 29'b0_010101010001_101_0_100101010100;
      patterns[10894] = 29'b0_010101010001_110_0_010101010001;
      patterns[10895] = 29'b0_010101010001_111_0_010101010001;
      patterns[10896] = 29'b0_010101010010_000_0_010101010010;
      patterns[10897] = 29'b0_010101010010_001_0_010010010101;
      patterns[10898] = 29'b0_010101010010_010_0_101010100100;
      patterns[10899] = 29'b0_010101010010_011_1_010101001000;
      patterns[10900] = 29'b0_010101010010_100_0_001010101001;
      patterns[10901] = 29'b0_010101010010_101_1_000101010100;
      patterns[10902] = 29'b0_010101010010_110_0_010101010010;
      patterns[10903] = 29'b0_010101010010_111_0_010101010010;
      patterns[10904] = 29'b0_010101010011_000_0_010101010011;
      patterns[10905] = 29'b0_010101010011_001_0_010011010101;
      patterns[10906] = 29'b0_010101010011_010_0_101010100110;
      patterns[10907] = 29'b0_010101010011_011_1_010101001100;
      patterns[10908] = 29'b0_010101010011_100_1_001010101001;
      patterns[10909] = 29'b0_010101010011_101_1_100101010100;
      patterns[10910] = 29'b0_010101010011_110_0_010101010011;
      patterns[10911] = 29'b0_010101010011_111_0_010101010011;
      patterns[10912] = 29'b0_010101010100_000_0_010101010100;
      patterns[10913] = 29'b0_010101010100_001_0_010100010101;
      patterns[10914] = 29'b0_010101010100_010_0_101010101000;
      patterns[10915] = 29'b0_010101010100_011_1_010101010000;
      patterns[10916] = 29'b0_010101010100_100_0_001010101010;
      patterns[10917] = 29'b0_010101010100_101_0_000101010101;
      patterns[10918] = 29'b0_010101010100_110_0_010101010100;
      patterns[10919] = 29'b0_010101010100_111_0_010101010100;
      patterns[10920] = 29'b0_010101010101_000_0_010101010101;
      patterns[10921] = 29'b0_010101010101_001_0_010101010101;
      patterns[10922] = 29'b0_010101010101_010_0_101010101010;
      patterns[10923] = 29'b0_010101010101_011_1_010101010100;
      patterns[10924] = 29'b0_010101010101_100_1_001010101010;
      patterns[10925] = 29'b0_010101010101_101_0_100101010101;
      patterns[10926] = 29'b0_010101010101_110_0_010101010101;
      patterns[10927] = 29'b0_010101010101_111_0_010101010101;
      patterns[10928] = 29'b0_010101010110_000_0_010101010110;
      patterns[10929] = 29'b0_010101010110_001_0_010110010101;
      patterns[10930] = 29'b0_010101010110_010_0_101010101100;
      patterns[10931] = 29'b0_010101010110_011_1_010101011000;
      patterns[10932] = 29'b0_010101010110_100_0_001010101011;
      patterns[10933] = 29'b0_010101010110_101_1_000101010101;
      patterns[10934] = 29'b0_010101010110_110_0_010101010110;
      patterns[10935] = 29'b0_010101010110_111_0_010101010110;
      patterns[10936] = 29'b0_010101010111_000_0_010101010111;
      patterns[10937] = 29'b0_010101010111_001_0_010111010101;
      patterns[10938] = 29'b0_010101010111_010_0_101010101110;
      patterns[10939] = 29'b0_010101010111_011_1_010101011100;
      patterns[10940] = 29'b0_010101010111_100_1_001010101011;
      patterns[10941] = 29'b0_010101010111_101_1_100101010101;
      patterns[10942] = 29'b0_010101010111_110_0_010101010111;
      patterns[10943] = 29'b0_010101010111_111_0_010101010111;
      patterns[10944] = 29'b0_010101011000_000_0_010101011000;
      patterns[10945] = 29'b0_010101011000_001_0_011000010101;
      patterns[10946] = 29'b0_010101011000_010_0_101010110000;
      patterns[10947] = 29'b0_010101011000_011_1_010101100000;
      patterns[10948] = 29'b0_010101011000_100_0_001010101100;
      patterns[10949] = 29'b0_010101011000_101_0_000101010110;
      patterns[10950] = 29'b0_010101011000_110_0_010101011000;
      patterns[10951] = 29'b0_010101011000_111_0_010101011000;
      patterns[10952] = 29'b0_010101011001_000_0_010101011001;
      patterns[10953] = 29'b0_010101011001_001_0_011001010101;
      patterns[10954] = 29'b0_010101011001_010_0_101010110010;
      patterns[10955] = 29'b0_010101011001_011_1_010101100100;
      patterns[10956] = 29'b0_010101011001_100_1_001010101100;
      patterns[10957] = 29'b0_010101011001_101_0_100101010110;
      patterns[10958] = 29'b0_010101011001_110_0_010101011001;
      patterns[10959] = 29'b0_010101011001_111_0_010101011001;
      patterns[10960] = 29'b0_010101011010_000_0_010101011010;
      patterns[10961] = 29'b0_010101011010_001_0_011010010101;
      patterns[10962] = 29'b0_010101011010_010_0_101010110100;
      patterns[10963] = 29'b0_010101011010_011_1_010101101000;
      patterns[10964] = 29'b0_010101011010_100_0_001010101101;
      patterns[10965] = 29'b0_010101011010_101_1_000101010110;
      patterns[10966] = 29'b0_010101011010_110_0_010101011010;
      patterns[10967] = 29'b0_010101011010_111_0_010101011010;
      patterns[10968] = 29'b0_010101011011_000_0_010101011011;
      patterns[10969] = 29'b0_010101011011_001_0_011011010101;
      patterns[10970] = 29'b0_010101011011_010_0_101010110110;
      patterns[10971] = 29'b0_010101011011_011_1_010101101100;
      patterns[10972] = 29'b0_010101011011_100_1_001010101101;
      patterns[10973] = 29'b0_010101011011_101_1_100101010110;
      patterns[10974] = 29'b0_010101011011_110_0_010101011011;
      patterns[10975] = 29'b0_010101011011_111_0_010101011011;
      patterns[10976] = 29'b0_010101011100_000_0_010101011100;
      patterns[10977] = 29'b0_010101011100_001_0_011100010101;
      patterns[10978] = 29'b0_010101011100_010_0_101010111000;
      patterns[10979] = 29'b0_010101011100_011_1_010101110000;
      patterns[10980] = 29'b0_010101011100_100_0_001010101110;
      patterns[10981] = 29'b0_010101011100_101_0_000101010111;
      patterns[10982] = 29'b0_010101011100_110_0_010101011100;
      patterns[10983] = 29'b0_010101011100_111_0_010101011100;
      patterns[10984] = 29'b0_010101011101_000_0_010101011101;
      patterns[10985] = 29'b0_010101011101_001_0_011101010101;
      patterns[10986] = 29'b0_010101011101_010_0_101010111010;
      patterns[10987] = 29'b0_010101011101_011_1_010101110100;
      patterns[10988] = 29'b0_010101011101_100_1_001010101110;
      patterns[10989] = 29'b0_010101011101_101_0_100101010111;
      patterns[10990] = 29'b0_010101011101_110_0_010101011101;
      patterns[10991] = 29'b0_010101011101_111_0_010101011101;
      patterns[10992] = 29'b0_010101011110_000_0_010101011110;
      patterns[10993] = 29'b0_010101011110_001_0_011110010101;
      patterns[10994] = 29'b0_010101011110_010_0_101010111100;
      patterns[10995] = 29'b0_010101011110_011_1_010101111000;
      patterns[10996] = 29'b0_010101011110_100_0_001010101111;
      patterns[10997] = 29'b0_010101011110_101_1_000101010111;
      patterns[10998] = 29'b0_010101011110_110_0_010101011110;
      patterns[10999] = 29'b0_010101011110_111_0_010101011110;
      patterns[11000] = 29'b0_010101011111_000_0_010101011111;
      patterns[11001] = 29'b0_010101011111_001_0_011111010101;
      patterns[11002] = 29'b0_010101011111_010_0_101010111110;
      patterns[11003] = 29'b0_010101011111_011_1_010101111100;
      patterns[11004] = 29'b0_010101011111_100_1_001010101111;
      patterns[11005] = 29'b0_010101011111_101_1_100101010111;
      patterns[11006] = 29'b0_010101011111_110_0_010101011111;
      patterns[11007] = 29'b0_010101011111_111_0_010101011111;
      patterns[11008] = 29'b0_010101100000_000_0_010101100000;
      patterns[11009] = 29'b0_010101100000_001_0_100000010101;
      patterns[11010] = 29'b0_010101100000_010_0_101011000000;
      patterns[11011] = 29'b0_010101100000_011_1_010110000000;
      patterns[11012] = 29'b0_010101100000_100_0_001010110000;
      patterns[11013] = 29'b0_010101100000_101_0_000101011000;
      patterns[11014] = 29'b0_010101100000_110_0_010101100000;
      patterns[11015] = 29'b0_010101100000_111_0_010101100000;
      patterns[11016] = 29'b0_010101100001_000_0_010101100001;
      patterns[11017] = 29'b0_010101100001_001_0_100001010101;
      patterns[11018] = 29'b0_010101100001_010_0_101011000010;
      patterns[11019] = 29'b0_010101100001_011_1_010110000100;
      patterns[11020] = 29'b0_010101100001_100_1_001010110000;
      patterns[11021] = 29'b0_010101100001_101_0_100101011000;
      patterns[11022] = 29'b0_010101100001_110_0_010101100001;
      patterns[11023] = 29'b0_010101100001_111_0_010101100001;
      patterns[11024] = 29'b0_010101100010_000_0_010101100010;
      patterns[11025] = 29'b0_010101100010_001_0_100010010101;
      patterns[11026] = 29'b0_010101100010_010_0_101011000100;
      patterns[11027] = 29'b0_010101100010_011_1_010110001000;
      patterns[11028] = 29'b0_010101100010_100_0_001010110001;
      patterns[11029] = 29'b0_010101100010_101_1_000101011000;
      patterns[11030] = 29'b0_010101100010_110_0_010101100010;
      patterns[11031] = 29'b0_010101100010_111_0_010101100010;
      patterns[11032] = 29'b0_010101100011_000_0_010101100011;
      patterns[11033] = 29'b0_010101100011_001_0_100011010101;
      patterns[11034] = 29'b0_010101100011_010_0_101011000110;
      patterns[11035] = 29'b0_010101100011_011_1_010110001100;
      patterns[11036] = 29'b0_010101100011_100_1_001010110001;
      patterns[11037] = 29'b0_010101100011_101_1_100101011000;
      patterns[11038] = 29'b0_010101100011_110_0_010101100011;
      patterns[11039] = 29'b0_010101100011_111_0_010101100011;
      patterns[11040] = 29'b0_010101100100_000_0_010101100100;
      patterns[11041] = 29'b0_010101100100_001_0_100100010101;
      patterns[11042] = 29'b0_010101100100_010_0_101011001000;
      patterns[11043] = 29'b0_010101100100_011_1_010110010000;
      patterns[11044] = 29'b0_010101100100_100_0_001010110010;
      patterns[11045] = 29'b0_010101100100_101_0_000101011001;
      patterns[11046] = 29'b0_010101100100_110_0_010101100100;
      patterns[11047] = 29'b0_010101100100_111_0_010101100100;
      patterns[11048] = 29'b0_010101100101_000_0_010101100101;
      patterns[11049] = 29'b0_010101100101_001_0_100101010101;
      patterns[11050] = 29'b0_010101100101_010_0_101011001010;
      patterns[11051] = 29'b0_010101100101_011_1_010110010100;
      patterns[11052] = 29'b0_010101100101_100_1_001010110010;
      patterns[11053] = 29'b0_010101100101_101_0_100101011001;
      patterns[11054] = 29'b0_010101100101_110_0_010101100101;
      patterns[11055] = 29'b0_010101100101_111_0_010101100101;
      patterns[11056] = 29'b0_010101100110_000_0_010101100110;
      patterns[11057] = 29'b0_010101100110_001_0_100110010101;
      patterns[11058] = 29'b0_010101100110_010_0_101011001100;
      patterns[11059] = 29'b0_010101100110_011_1_010110011000;
      patterns[11060] = 29'b0_010101100110_100_0_001010110011;
      patterns[11061] = 29'b0_010101100110_101_1_000101011001;
      patterns[11062] = 29'b0_010101100110_110_0_010101100110;
      patterns[11063] = 29'b0_010101100110_111_0_010101100110;
      patterns[11064] = 29'b0_010101100111_000_0_010101100111;
      patterns[11065] = 29'b0_010101100111_001_0_100111010101;
      patterns[11066] = 29'b0_010101100111_010_0_101011001110;
      patterns[11067] = 29'b0_010101100111_011_1_010110011100;
      patterns[11068] = 29'b0_010101100111_100_1_001010110011;
      patterns[11069] = 29'b0_010101100111_101_1_100101011001;
      patterns[11070] = 29'b0_010101100111_110_0_010101100111;
      patterns[11071] = 29'b0_010101100111_111_0_010101100111;
      patterns[11072] = 29'b0_010101101000_000_0_010101101000;
      patterns[11073] = 29'b0_010101101000_001_0_101000010101;
      patterns[11074] = 29'b0_010101101000_010_0_101011010000;
      patterns[11075] = 29'b0_010101101000_011_1_010110100000;
      patterns[11076] = 29'b0_010101101000_100_0_001010110100;
      patterns[11077] = 29'b0_010101101000_101_0_000101011010;
      patterns[11078] = 29'b0_010101101000_110_0_010101101000;
      patterns[11079] = 29'b0_010101101000_111_0_010101101000;
      patterns[11080] = 29'b0_010101101001_000_0_010101101001;
      patterns[11081] = 29'b0_010101101001_001_0_101001010101;
      patterns[11082] = 29'b0_010101101001_010_0_101011010010;
      patterns[11083] = 29'b0_010101101001_011_1_010110100100;
      patterns[11084] = 29'b0_010101101001_100_1_001010110100;
      patterns[11085] = 29'b0_010101101001_101_0_100101011010;
      patterns[11086] = 29'b0_010101101001_110_0_010101101001;
      patterns[11087] = 29'b0_010101101001_111_0_010101101001;
      patterns[11088] = 29'b0_010101101010_000_0_010101101010;
      patterns[11089] = 29'b0_010101101010_001_0_101010010101;
      patterns[11090] = 29'b0_010101101010_010_0_101011010100;
      patterns[11091] = 29'b0_010101101010_011_1_010110101000;
      patterns[11092] = 29'b0_010101101010_100_0_001010110101;
      patterns[11093] = 29'b0_010101101010_101_1_000101011010;
      patterns[11094] = 29'b0_010101101010_110_0_010101101010;
      patterns[11095] = 29'b0_010101101010_111_0_010101101010;
      patterns[11096] = 29'b0_010101101011_000_0_010101101011;
      patterns[11097] = 29'b0_010101101011_001_0_101011010101;
      patterns[11098] = 29'b0_010101101011_010_0_101011010110;
      patterns[11099] = 29'b0_010101101011_011_1_010110101100;
      patterns[11100] = 29'b0_010101101011_100_1_001010110101;
      patterns[11101] = 29'b0_010101101011_101_1_100101011010;
      patterns[11102] = 29'b0_010101101011_110_0_010101101011;
      patterns[11103] = 29'b0_010101101011_111_0_010101101011;
      patterns[11104] = 29'b0_010101101100_000_0_010101101100;
      patterns[11105] = 29'b0_010101101100_001_0_101100010101;
      patterns[11106] = 29'b0_010101101100_010_0_101011011000;
      patterns[11107] = 29'b0_010101101100_011_1_010110110000;
      patterns[11108] = 29'b0_010101101100_100_0_001010110110;
      patterns[11109] = 29'b0_010101101100_101_0_000101011011;
      patterns[11110] = 29'b0_010101101100_110_0_010101101100;
      patterns[11111] = 29'b0_010101101100_111_0_010101101100;
      patterns[11112] = 29'b0_010101101101_000_0_010101101101;
      patterns[11113] = 29'b0_010101101101_001_0_101101010101;
      patterns[11114] = 29'b0_010101101101_010_0_101011011010;
      patterns[11115] = 29'b0_010101101101_011_1_010110110100;
      patterns[11116] = 29'b0_010101101101_100_1_001010110110;
      patterns[11117] = 29'b0_010101101101_101_0_100101011011;
      patterns[11118] = 29'b0_010101101101_110_0_010101101101;
      patterns[11119] = 29'b0_010101101101_111_0_010101101101;
      patterns[11120] = 29'b0_010101101110_000_0_010101101110;
      patterns[11121] = 29'b0_010101101110_001_0_101110010101;
      patterns[11122] = 29'b0_010101101110_010_0_101011011100;
      patterns[11123] = 29'b0_010101101110_011_1_010110111000;
      patterns[11124] = 29'b0_010101101110_100_0_001010110111;
      patterns[11125] = 29'b0_010101101110_101_1_000101011011;
      patterns[11126] = 29'b0_010101101110_110_0_010101101110;
      patterns[11127] = 29'b0_010101101110_111_0_010101101110;
      patterns[11128] = 29'b0_010101101111_000_0_010101101111;
      patterns[11129] = 29'b0_010101101111_001_0_101111010101;
      patterns[11130] = 29'b0_010101101111_010_0_101011011110;
      patterns[11131] = 29'b0_010101101111_011_1_010110111100;
      patterns[11132] = 29'b0_010101101111_100_1_001010110111;
      patterns[11133] = 29'b0_010101101111_101_1_100101011011;
      patterns[11134] = 29'b0_010101101111_110_0_010101101111;
      patterns[11135] = 29'b0_010101101111_111_0_010101101111;
      patterns[11136] = 29'b0_010101110000_000_0_010101110000;
      patterns[11137] = 29'b0_010101110000_001_0_110000010101;
      patterns[11138] = 29'b0_010101110000_010_0_101011100000;
      patterns[11139] = 29'b0_010101110000_011_1_010111000000;
      patterns[11140] = 29'b0_010101110000_100_0_001010111000;
      patterns[11141] = 29'b0_010101110000_101_0_000101011100;
      patterns[11142] = 29'b0_010101110000_110_0_010101110000;
      patterns[11143] = 29'b0_010101110000_111_0_010101110000;
      patterns[11144] = 29'b0_010101110001_000_0_010101110001;
      patterns[11145] = 29'b0_010101110001_001_0_110001010101;
      patterns[11146] = 29'b0_010101110001_010_0_101011100010;
      patterns[11147] = 29'b0_010101110001_011_1_010111000100;
      patterns[11148] = 29'b0_010101110001_100_1_001010111000;
      patterns[11149] = 29'b0_010101110001_101_0_100101011100;
      patterns[11150] = 29'b0_010101110001_110_0_010101110001;
      patterns[11151] = 29'b0_010101110001_111_0_010101110001;
      patterns[11152] = 29'b0_010101110010_000_0_010101110010;
      patterns[11153] = 29'b0_010101110010_001_0_110010010101;
      patterns[11154] = 29'b0_010101110010_010_0_101011100100;
      patterns[11155] = 29'b0_010101110010_011_1_010111001000;
      patterns[11156] = 29'b0_010101110010_100_0_001010111001;
      patterns[11157] = 29'b0_010101110010_101_1_000101011100;
      patterns[11158] = 29'b0_010101110010_110_0_010101110010;
      patterns[11159] = 29'b0_010101110010_111_0_010101110010;
      patterns[11160] = 29'b0_010101110011_000_0_010101110011;
      patterns[11161] = 29'b0_010101110011_001_0_110011010101;
      patterns[11162] = 29'b0_010101110011_010_0_101011100110;
      patterns[11163] = 29'b0_010101110011_011_1_010111001100;
      patterns[11164] = 29'b0_010101110011_100_1_001010111001;
      patterns[11165] = 29'b0_010101110011_101_1_100101011100;
      patterns[11166] = 29'b0_010101110011_110_0_010101110011;
      patterns[11167] = 29'b0_010101110011_111_0_010101110011;
      patterns[11168] = 29'b0_010101110100_000_0_010101110100;
      patterns[11169] = 29'b0_010101110100_001_0_110100010101;
      patterns[11170] = 29'b0_010101110100_010_0_101011101000;
      patterns[11171] = 29'b0_010101110100_011_1_010111010000;
      patterns[11172] = 29'b0_010101110100_100_0_001010111010;
      patterns[11173] = 29'b0_010101110100_101_0_000101011101;
      patterns[11174] = 29'b0_010101110100_110_0_010101110100;
      patterns[11175] = 29'b0_010101110100_111_0_010101110100;
      patterns[11176] = 29'b0_010101110101_000_0_010101110101;
      patterns[11177] = 29'b0_010101110101_001_0_110101010101;
      patterns[11178] = 29'b0_010101110101_010_0_101011101010;
      patterns[11179] = 29'b0_010101110101_011_1_010111010100;
      patterns[11180] = 29'b0_010101110101_100_1_001010111010;
      patterns[11181] = 29'b0_010101110101_101_0_100101011101;
      patterns[11182] = 29'b0_010101110101_110_0_010101110101;
      patterns[11183] = 29'b0_010101110101_111_0_010101110101;
      patterns[11184] = 29'b0_010101110110_000_0_010101110110;
      patterns[11185] = 29'b0_010101110110_001_0_110110010101;
      patterns[11186] = 29'b0_010101110110_010_0_101011101100;
      patterns[11187] = 29'b0_010101110110_011_1_010111011000;
      patterns[11188] = 29'b0_010101110110_100_0_001010111011;
      patterns[11189] = 29'b0_010101110110_101_1_000101011101;
      patterns[11190] = 29'b0_010101110110_110_0_010101110110;
      patterns[11191] = 29'b0_010101110110_111_0_010101110110;
      patterns[11192] = 29'b0_010101110111_000_0_010101110111;
      patterns[11193] = 29'b0_010101110111_001_0_110111010101;
      patterns[11194] = 29'b0_010101110111_010_0_101011101110;
      patterns[11195] = 29'b0_010101110111_011_1_010111011100;
      patterns[11196] = 29'b0_010101110111_100_1_001010111011;
      patterns[11197] = 29'b0_010101110111_101_1_100101011101;
      patterns[11198] = 29'b0_010101110111_110_0_010101110111;
      patterns[11199] = 29'b0_010101110111_111_0_010101110111;
      patterns[11200] = 29'b0_010101111000_000_0_010101111000;
      patterns[11201] = 29'b0_010101111000_001_0_111000010101;
      patterns[11202] = 29'b0_010101111000_010_0_101011110000;
      patterns[11203] = 29'b0_010101111000_011_1_010111100000;
      patterns[11204] = 29'b0_010101111000_100_0_001010111100;
      patterns[11205] = 29'b0_010101111000_101_0_000101011110;
      patterns[11206] = 29'b0_010101111000_110_0_010101111000;
      patterns[11207] = 29'b0_010101111000_111_0_010101111000;
      patterns[11208] = 29'b0_010101111001_000_0_010101111001;
      patterns[11209] = 29'b0_010101111001_001_0_111001010101;
      patterns[11210] = 29'b0_010101111001_010_0_101011110010;
      patterns[11211] = 29'b0_010101111001_011_1_010111100100;
      patterns[11212] = 29'b0_010101111001_100_1_001010111100;
      patterns[11213] = 29'b0_010101111001_101_0_100101011110;
      patterns[11214] = 29'b0_010101111001_110_0_010101111001;
      patterns[11215] = 29'b0_010101111001_111_0_010101111001;
      patterns[11216] = 29'b0_010101111010_000_0_010101111010;
      patterns[11217] = 29'b0_010101111010_001_0_111010010101;
      patterns[11218] = 29'b0_010101111010_010_0_101011110100;
      patterns[11219] = 29'b0_010101111010_011_1_010111101000;
      patterns[11220] = 29'b0_010101111010_100_0_001010111101;
      patterns[11221] = 29'b0_010101111010_101_1_000101011110;
      patterns[11222] = 29'b0_010101111010_110_0_010101111010;
      patterns[11223] = 29'b0_010101111010_111_0_010101111010;
      patterns[11224] = 29'b0_010101111011_000_0_010101111011;
      patterns[11225] = 29'b0_010101111011_001_0_111011010101;
      patterns[11226] = 29'b0_010101111011_010_0_101011110110;
      patterns[11227] = 29'b0_010101111011_011_1_010111101100;
      patterns[11228] = 29'b0_010101111011_100_1_001010111101;
      patterns[11229] = 29'b0_010101111011_101_1_100101011110;
      patterns[11230] = 29'b0_010101111011_110_0_010101111011;
      patterns[11231] = 29'b0_010101111011_111_0_010101111011;
      patterns[11232] = 29'b0_010101111100_000_0_010101111100;
      patterns[11233] = 29'b0_010101111100_001_0_111100010101;
      patterns[11234] = 29'b0_010101111100_010_0_101011111000;
      patterns[11235] = 29'b0_010101111100_011_1_010111110000;
      patterns[11236] = 29'b0_010101111100_100_0_001010111110;
      patterns[11237] = 29'b0_010101111100_101_0_000101011111;
      patterns[11238] = 29'b0_010101111100_110_0_010101111100;
      patterns[11239] = 29'b0_010101111100_111_0_010101111100;
      patterns[11240] = 29'b0_010101111101_000_0_010101111101;
      patterns[11241] = 29'b0_010101111101_001_0_111101010101;
      patterns[11242] = 29'b0_010101111101_010_0_101011111010;
      patterns[11243] = 29'b0_010101111101_011_1_010111110100;
      patterns[11244] = 29'b0_010101111101_100_1_001010111110;
      patterns[11245] = 29'b0_010101111101_101_0_100101011111;
      patterns[11246] = 29'b0_010101111101_110_0_010101111101;
      patterns[11247] = 29'b0_010101111101_111_0_010101111101;
      patterns[11248] = 29'b0_010101111110_000_0_010101111110;
      patterns[11249] = 29'b0_010101111110_001_0_111110010101;
      patterns[11250] = 29'b0_010101111110_010_0_101011111100;
      patterns[11251] = 29'b0_010101111110_011_1_010111111000;
      patterns[11252] = 29'b0_010101111110_100_0_001010111111;
      patterns[11253] = 29'b0_010101111110_101_1_000101011111;
      patterns[11254] = 29'b0_010101111110_110_0_010101111110;
      patterns[11255] = 29'b0_010101111110_111_0_010101111110;
      patterns[11256] = 29'b0_010101111111_000_0_010101111111;
      patterns[11257] = 29'b0_010101111111_001_0_111111010101;
      patterns[11258] = 29'b0_010101111111_010_0_101011111110;
      patterns[11259] = 29'b0_010101111111_011_1_010111111100;
      patterns[11260] = 29'b0_010101111111_100_1_001010111111;
      patterns[11261] = 29'b0_010101111111_101_1_100101011111;
      patterns[11262] = 29'b0_010101111111_110_0_010101111111;
      patterns[11263] = 29'b0_010101111111_111_0_010101111111;
      patterns[11264] = 29'b0_010110000000_000_0_010110000000;
      patterns[11265] = 29'b0_010110000000_001_0_000000010110;
      patterns[11266] = 29'b0_010110000000_010_0_101100000000;
      patterns[11267] = 29'b0_010110000000_011_1_011000000000;
      patterns[11268] = 29'b0_010110000000_100_0_001011000000;
      patterns[11269] = 29'b0_010110000000_101_0_000101100000;
      patterns[11270] = 29'b0_010110000000_110_0_010110000000;
      patterns[11271] = 29'b0_010110000000_111_0_010110000000;
      patterns[11272] = 29'b0_010110000001_000_0_010110000001;
      patterns[11273] = 29'b0_010110000001_001_0_000001010110;
      patterns[11274] = 29'b0_010110000001_010_0_101100000010;
      patterns[11275] = 29'b0_010110000001_011_1_011000000100;
      patterns[11276] = 29'b0_010110000001_100_1_001011000000;
      patterns[11277] = 29'b0_010110000001_101_0_100101100000;
      patterns[11278] = 29'b0_010110000001_110_0_010110000001;
      patterns[11279] = 29'b0_010110000001_111_0_010110000001;
      patterns[11280] = 29'b0_010110000010_000_0_010110000010;
      patterns[11281] = 29'b0_010110000010_001_0_000010010110;
      patterns[11282] = 29'b0_010110000010_010_0_101100000100;
      patterns[11283] = 29'b0_010110000010_011_1_011000001000;
      patterns[11284] = 29'b0_010110000010_100_0_001011000001;
      patterns[11285] = 29'b0_010110000010_101_1_000101100000;
      patterns[11286] = 29'b0_010110000010_110_0_010110000010;
      patterns[11287] = 29'b0_010110000010_111_0_010110000010;
      patterns[11288] = 29'b0_010110000011_000_0_010110000011;
      patterns[11289] = 29'b0_010110000011_001_0_000011010110;
      patterns[11290] = 29'b0_010110000011_010_0_101100000110;
      patterns[11291] = 29'b0_010110000011_011_1_011000001100;
      patterns[11292] = 29'b0_010110000011_100_1_001011000001;
      patterns[11293] = 29'b0_010110000011_101_1_100101100000;
      patterns[11294] = 29'b0_010110000011_110_0_010110000011;
      patterns[11295] = 29'b0_010110000011_111_0_010110000011;
      patterns[11296] = 29'b0_010110000100_000_0_010110000100;
      patterns[11297] = 29'b0_010110000100_001_0_000100010110;
      patterns[11298] = 29'b0_010110000100_010_0_101100001000;
      patterns[11299] = 29'b0_010110000100_011_1_011000010000;
      patterns[11300] = 29'b0_010110000100_100_0_001011000010;
      patterns[11301] = 29'b0_010110000100_101_0_000101100001;
      patterns[11302] = 29'b0_010110000100_110_0_010110000100;
      patterns[11303] = 29'b0_010110000100_111_0_010110000100;
      patterns[11304] = 29'b0_010110000101_000_0_010110000101;
      patterns[11305] = 29'b0_010110000101_001_0_000101010110;
      patterns[11306] = 29'b0_010110000101_010_0_101100001010;
      patterns[11307] = 29'b0_010110000101_011_1_011000010100;
      patterns[11308] = 29'b0_010110000101_100_1_001011000010;
      patterns[11309] = 29'b0_010110000101_101_0_100101100001;
      patterns[11310] = 29'b0_010110000101_110_0_010110000101;
      patterns[11311] = 29'b0_010110000101_111_0_010110000101;
      patterns[11312] = 29'b0_010110000110_000_0_010110000110;
      patterns[11313] = 29'b0_010110000110_001_0_000110010110;
      patterns[11314] = 29'b0_010110000110_010_0_101100001100;
      patterns[11315] = 29'b0_010110000110_011_1_011000011000;
      patterns[11316] = 29'b0_010110000110_100_0_001011000011;
      patterns[11317] = 29'b0_010110000110_101_1_000101100001;
      patterns[11318] = 29'b0_010110000110_110_0_010110000110;
      patterns[11319] = 29'b0_010110000110_111_0_010110000110;
      patterns[11320] = 29'b0_010110000111_000_0_010110000111;
      patterns[11321] = 29'b0_010110000111_001_0_000111010110;
      patterns[11322] = 29'b0_010110000111_010_0_101100001110;
      patterns[11323] = 29'b0_010110000111_011_1_011000011100;
      patterns[11324] = 29'b0_010110000111_100_1_001011000011;
      patterns[11325] = 29'b0_010110000111_101_1_100101100001;
      patterns[11326] = 29'b0_010110000111_110_0_010110000111;
      patterns[11327] = 29'b0_010110000111_111_0_010110000111;
      patterns[11328] = 29'b0_010110001000_000_0_010110001000;
      patterns[11329] = 29'b0_010110001000_001_0_001000010110;
      patterns[11330] = 29'b0_010110001000_010_0_101100010000;
      patterns[11331] = 29'b0_010110001000_011_1_011000100000;
      patterns[11332] = 29'b0_010110001000_100_0_001011000100;
      patterns[11333] = 29'b0_010110001000_101_0_000101100010;
      patterns[11334] = 29'b0_010110001000_110_0_010110001000;
      patterns[11335] = 29'b0_010110001000_111_0_010110001000;
      patterns[11336] = 29'b0_010110001001_000_0_010110001001;
      patterns[11337] = 29'b0_010110001001_001_0_001001010110;
      patterns[11338] = 29'b0_010110001001_010_0_101100010010;
      patterns[11339] = 29'b0_010110001001_011_1_011000100100;
      patterns[11340] = 29'b0_010110001001_100_1_001011000100;
      patterns[11341] = 29'b0_010110001001_101_0_100101100010;
      patterns[11342] = 29'b0_010110001001_110_0_010110001001;
      patterns[11343] = 29'b0_010110001001_111_0_010110001001;
      patterns[11344] = 29'b0_010110001010_000_0_010110001010;
      patterns[11345] = 29'b0_010110001010_001_0_001010010110;
      patterns[11346] = 29'b0_010110001010_010_0_101100010100;
      patterns[11347] = 29'b0_010110001010_011_1_011000101000;
      patterns[11348] = 29'b0_010110001010_100_0_001011000101;
      patterns[11349] = 29'b0_010110001010_101_1_000101100010;
      patterns[11350] = 29'b0_010110001010_110_0_010110001010;
      patterns[11351] = 29'b0_010110001010_111_0_010110001010;
      patterns[11352] = 29'b0_010110001011_000_0_010110001011;
      patterns[11353] = 29'b0_010110001011_001_0_001011010110;
      patterns[11354] = 29'b0_010110001011_010_0_101100010110;
      patterns[11355] = 29'b0_010110001011_011_1_011000101100;
      patterns[11356] = 29'b0_010110001011_100_1_001011000101;
      patterns[11357] = 29'b0_010110001011_101_1_100101100010;
      patterns[11358] = 29'b0_010110001011_110_0_010110001011;
      patterns[11359] = 29'b0_010110001011_111_0_010110001011;
      patterns[11360] = 29'b0_010110001100_000_0_010110001100;
      patterns[11361] = 29'b0_010110001100_001_0_001100010110;
      patterns[11362] = 29'b0_010110001100_010_0_101100011000;
      patterns[11363] = 29'b0_010110001100_011_1_011000110000;
      patterns[11364] = 29'b0_010110001100_100_0_001011000110;
      patterns[11365] = 29'b0_010110001100_101_0_000101100011;
      patterns[11366] = 29'b0_010110001100_110_0_010110001100;
      patterns[11367] = 29'b0_010110001100_111_0_010110001100;
      patterns[11368] = 29'b0_010110001101_000_0_010110001101;
      patterns[11369] = 29'b0_010110001101_001_0_001101010110;
      patterns[11370] = 29'b0_010110001101_010_0_101100011010;
      patterns[11371] = 29'b0_010110001101_011_1_011000110100;
      patterns[11372] = 29'b0_010110001101_100_1_001011000110;
      patterns[11373] = 29'b0_010110001101_101_0_100101100011;
      patterns[11374] = 29'b0_010110001101_110_0_010110001101;
      patterns[11375] = 29'b0_010110001101_111_0_010110001101;
      patterns[11376] = 29'b0_010110001110_000_0_010110001110;
      patterns[11377] = 29'b0_010110001110_001_0_001110010110;
      patterns[11378] = 29'b0_010110001110_010_0_101100011100;
      patterns[11379] = 29'b0_010110001110_011_1_011000111000;
      patterns[11380] = 29'b0_010110001110_100_0_001011000111;
      patterns[11381] = 29'b0_010110001110_101_1_000101100011;
      patterns[11382] = 29'b0_010110001110_110_0_010110001110;
      patterns[11383] = 29'b0_010110001110_111_0_010110001110;
      patterns[11384] = 29'b0_010110001111_000_0_010110001111;
      patterns[11385] = 29'b0_010110001111_001_0_001111010110;
      patterns[11386] = 29'b0_010110001111_010_0_101100011110;
      patterns[11387] = 29'b0_010110001111_011_1_011000111100;
      patterns[11388] = 29'b0_010110001111_100_1_001011000111;
      patterns[11389] = 29'b0_010110001111_101_1_100101100011;
      patterns[11390] = 29'b0_010110001111_110_0_010110001111;
      patterns[11391] = 29'b0_010110001111_111_0_010110001111;
      patterns[11392] = 29'b0_010110010000_000_0_010110010000;
      patterns[11393] = 29'b0_010110010000_001_0_010000010110;
      patterns[11394] = 29'b0_010110010000_010_0_101100100000;
      patterns[11395] = 29'b0_010110010000_011_1_011001000000;
      patterns[11396] = 29'b0_010110010000_100_0_001011001000;
      patterns[11397] = 29'b0_010110010000_101_0_000101100100;
      patterns[11398] = 29'b0_010110010000_110_0_010110010000;
      patterns[11399] = 29'b0_010110010000_111_0_010110010000;
      patterns[11400] = 29'b0_010110010001_000_0_010110010001;
      patterns[11401] = 29'b0_010110010001_001_0_010001010110;
      patterns[11402] = 29'b0_010110010001_010_0_101100100010;
      patterns[11403] = 29'b0_010110010001_011_1_011001000100;
      patterns[11404] = 29'b0_010110010001_100_1_001011001000;
      patterns[11405] = 29'b0_010110010001_101_0_100101100100;
      patterns[11406] = 29'b0_010110010001_110_0_010110010001;
      patterns[11407] = 29'b0_010110010001_111_0_010110010001;
      patterns[11408] = 29'b0_010110010010_000_0_010110010010;
      patterns[11409] = 29'b0_010110010010_001_0_010010010110;
      patterns[11410] = 29'b0_010110010010_010_0_101100100100;
      patterns[11411] = 29'b0_010110010010_011_1_011001001000;
      patterns[11412] = 29'b0_010110010010_100_0_001011001001;
      patterns[11413] = 29'b0_010110010010_101_1_000101100100;
      patterns[11414] = 29'b0_010110010010_110_0_010110010010;
      patterns[11415] = 29'b0_010110010010_111_0_010110010010;
      patterns[11416] = 29'b0_010110010011_000_0_010110010011;
      patterns[11417] = 29'b0_010110010011_001_0_010011010110;
      patterns[11418] = 29'b0_010110010011_010_0_101100100110;
      patterns[11419] = 29'b0_010110010011_011_1_011001001100;
      patterns[11420] = 29'b0_010110010011_100_1_001011001001;
      patterns[11421] = 29'b0_010110010011_101_1_100101100100;
      patterns[11422] = 29'b0_010110010011_110_0_010110010011;
      patterns[11423] = 29'b0_010110010011_111_0_010110010011;
      patterns[11424] = 29'b0_010110010100_000_0_010110010100;
      patterns[11425] = 29'b0_010110010100_001_0_010100010110;
      patterns[11426] = 29'b0_010110010100_010_0_101100101000;
      patterns[11427] = 29'b0_010110010100_011_1_011001010000;
      patterns[11428] = 29'b0_010110010100_100_0_001011001010;
      patterns[11429] = 29'b0_010110010100_101_0_000101100101;
      patterns[11430] = 29'b0_010110010100_110_0_010110010100;
      patterns[11431] = 29'b0_010110010100_111_0_010110010100;
      patterns[11432] = 29'b0_010110010101_000_0_010110010101;
      patterns[11433] = 29'b0_010110010101_001_0_010101010110;
      patterns[11434] = 29'b0_010110010101_010_0_101100101010;
      patterns[11435] = 29'b0_010110010101_011_1_011001010100;
      patterns[11436] = 29'b0_010110010101_100_1_001011001010;
      patterns[11437] = 29'b0_010110010101_101_0_100101100101;
      patterns[11438] = 29'b0_010110010101_110_0_010110010101;
      patterns[11439] = 29'b0_010110010101_111_0_010110010101;
      patterns[11440] = 29'b0_010110010110_000_0_010110010110;
      patterns[11441] = 29'b0_010110010110_001_0_010110010110;
      patterns[11442] = 29'b0_010110010110_010_0_101100101100;
      patterns[11443] = 29'b0_010110010110_011_1_011001011000;
      patterns[11444] = 29'b0_010110010110_100_0_001011001011;
      patterns[11445] = 29'b0_010110010110_101_1_000101100101;
      patterns[11446] = 29'b0_010110010110_110_0_010110010110;
      patterns[11447] = 29'b0_010110010110_111_0_010110010110;
      patterns[11448] = 29'b0_010110010111_000_0_010110010111;
      patterns[11449] = 29'b0_010110010111_001_0_010111010110;
      patterns[11450] = 29'b0_010110010111_010_0_101100101110;
      patterns[11451] = 29'b0_010110010111_011_1_011001011100;
      patterns[11452] = 29'b0_010110010111_100_1_001011001011;
      patterns[11453] = 29'b0_010110010111_101_1_100101100101;
      patterns[11454] = 29'b0_010110010111_110_0_010110010111;
      patterns[11455] = 29'b0_010110010111_111_0_010110010111;
      patterns[11456] = 29'b0_010110011000_000_0_010110011000;
      patterns[11457] = 29'b0_010110011000_001_0_011000010110;
      patterns[11458] = 29'b0_010110011000_010_0_101100110000;
      patterns[11459] = 29'b0_010110011000_011_1_011001100000;
      patterns[11460] = 29'b0_010110011000_100_0_001011001100;
      patterns[11461] = 29'b0_010110011000_101_0_000101100110;
      patterns[11462] = 29'b0_010110011000_110_0_010110011000;
      patterns[11463] = 29'b0_010110011000_111_0_010110011000;
      patterns[11464] = 29'b0_010110011001_000_0_010110011001;
      patterns[11465] = 29'b0_010110011001_001_0_011001010110;
      patterns[11466] = 29'b0_010110011001_010_0_101100110010;
      patterns[11467] = 29'b0_010110011001_011_1_011001100100;
      patterns[11468] = 29'b0_010110011001_100_1_001011001100;
      patterns[11469] = 29'b0_010110011001_101_0_100101100110;
      patterns[11470] = 29'b0_010110011001_110_0_010110011001;
      patterns[11471] = 29'b0_010110011001_111_0_010110011001;
      patterns[11472] = 29'b0_010110011010_000_0_010110011010;
      patterns[11473] = 29'b0_010110011010_001_0_011010010110;
      patterns[11474] = 29'b0_010110011010_010_0_101100110100;
      patterns[11475] = 29'b0_010110011010_011_1_011001101000;
      patterns[11476] = 29'b0_010110011010_100_0_001011001101;
      patterns[11477] = 29'b0_010110011010_101_1_000101100110;
      patterns[11478] = 29'b0_010110011010_110_0_010110011010;
      patterns[11479] = 29'b0_010110011010_111_0_010110011010;
      patterns[11480] = 29'b0_010110011011_000_0_010110011011;
      patterns[11481] = 29'b0_010110011011_001_0_011011010110;
      patterns[11482] = 29'b0_010110011011_010_0_101100110110;
      patterns[11483] = 29'b0_010110011011_011_1_011001101100;
      patterns[11484] = 29'b0_010110011011_100_1_001011001101;
      patterns[11485] = 29'b0_010110011011_101_1_100101100110;
      patterns[11486] = 29'b0_010110011011_110_0_010110011011;
      patterns[11487] = 29'b0_010110011011_111_0_010110011011;
      patterns[11488] = 29'b0_010110011100_000_0_010110011100;
      patterns[11489] = 29'b0_010110011100_001_0_011100010110;
      patterns[11490] = 29'b0_010110011100_010_0_101100111000;
      patterns[11491] = 29'b0_010110011100_011_1_011001110000;
      patterns[11492] = 29'b0_010110011100_100_0_001011001110;
      patterns[11493] = 29'b0_010110011100_101_0_000101100111;
      patterns[11494] = 29'b0_010110011100_110_0_010110011100;
      patterns[11495] = 29'b0_010110011100_111_0_010110011100;
      patterns[11496] = 29'b0_010110011101_000_0_010110011101;
      patterns[11497] = 29'b0_010110011101_001_0_011101010110;
      patterns[11498] = 29'b0_010110011101_010_0_101100111010;
      patterns[11499] = 29'b0_010110011101_011_1_011001110100;
      patterns[11500] = 29'b0_010110011101_100_1_001011001110;
      patterns[11501] = 29'b0_010110011101_101_0_100101100111;
      patterns[11502] = 29'b0_010110011101_110_0_010110011101;
      patterns[11503] = 29'b0_010110011101_111_0_010110011101;
      patterns[11504] = 29'b0_010110011110_000_0_010110011110;
      patterns[11505] = 29'b0_010110011110_001_0_011110010110;
      patterns[11506] = 29'b0_010110011110_010_0_101100111100;
      patterns[11507] = 29'b0_010110011110_011_1_011001111000;
      patterns[11508] = 29'b0_010110011110_100_0_001011001111;
      patterns[11509] = 29'b0_010110011110_101_1_000101100111;
      patterns[11510] = 29'b0_010110011110_110_0_010110011110;
      patterns[11511] = 29'b0_010110011110_111_0_010110011110;
      patterns[11512] = 29'b0_010110011111_000_0_010110011111;
      patterns[11513] = 29'b0_010110011111_001_0_011111010110;
      patterns[11514] = 29'b0_010110011111_010_0_101100111110;
      patterns[11515] = 29'b0_010110011111_011_1_011001111100;
      patterns[11516] = 29'b0_010110011111_100_1_001011001111;
      patterns[11517] = 29'b0_010110011111_101_1_100101100111;
      patterns[11518] = 29'b0_010110011111_110_0_010110011111;
      patterns[11519] = 29'b0_010110011111_111_0_010110011111;
      patterns[11520] = 29'b0_010110100000_000_0_010110100000;
      patterns[11521] = 29'b0_010110100000_001_0_100000010110;
      patterns[11522] = 29'b0_010110100000_010_0_101101000000;
      patterns[11523] = 29'b0_010110100000_011_1_011010000000;
      patterns[11524] = 29'b0_010110100000_100_0_001011010000;
      patterns[11525] = 29'b0_010110100000_101_0_000101101000;
      patterns[11526] = 29'b0_010110100000_110_0_010110100000;
      patterns[11527] = 29'b0_010110100000_111_0_010110100000;
      patterns[11528] = 29'b0_010110100001_000_0_010110100001;
      patterns[11529] = 29'b0_010110100001_001_0_100001010110;
      patterns[11530] = 29'b0_010110100001_010_0_101101000010;
      patterns[11531] = 29'b0_010110100001_011_1_011010000100;
      patterns[11532] = 29'b0_010110100001_100_1_001011010000;
      patterns[11533] = 29'b0_010110100001_101_0_100101101000;
      patterns[11534] = 29'b0_010110100001_110_0_010110100001;
      patterns[11535] = 29'b0_010110100001_111_0_010110100001;
      patterns[11536] = 29'b0_010110100010_000_0_010110100010;
      patterns[11537] = 29'b0_010110100010_001_0_100010010110;
      patterns[11538] = 29'b0_010110100010_010_0_101101000100;
      patterns[11539] = 29'b0_010110100010_011_1_011010001000;
      patterns[11540] = 29'b0_010110100010_100_0_001011010001;
      patterns[11541] = 29'b0_010110100010_101_1_000101101000;
      patterns[11542] = 29'b0_010110100010_110_0_010110100010;
      patterns[11543] = 29'b0_010110100010_111_0_010110100010;
      patterns[11544] = 29'b0_010110100011_000_0_010110100011;
      patterns[11545] = 29'b0_010110100011_001_0_100011010110;
      patterns[11546] = 29'b0_010110100011_010_0_101101000110;
      patterns[11547] = 29'b0_010110100011_011_1_011010001100;
      patterns[11548] = 29'b0_010110100011_100_1_001011010001;
      patterns[11549] = 29'b0_010110100011_101_1_100101101000;
      patterns[11550] = 29'b0_010110100011_110_0_010110100011;
      patterns[11551] = 29'b0_010110100011_111_0_010110100011;
      patterns[11552] = 29'b0_010110100100_000_0_010110100100;
      patterns[11553] = 29'b0_010110100100_001_0_100100010110;
      patterns[11554] = 29'b0_010110100100_010_0_101101001000;
      patterns[11555] = 29'b0_010110100100_011_1_011010010000;
      patterns[11556] = 29'b0_010110100100_100_0_001011010010;
      patterns[11557] = 29'b0_010110100100_101_0_000101101001;
      patterns[11558] = 29'b0_010110100100_110_0_010110100100;
      patterns[11559] = 29'b0_010110100100_111_0_010110100100;
      patterns[11560] = 29'b0_010110100101_000_0_010110100101;
      patterns[11561] = 29'b0_010110100101_001_0_100101010110;
      patterns[11562] = 29'b0_010110100101_010_0_101101001010;
      patterns[11563] = 29'b0_010110100101_011_1_011010010100;
      patterns[11564] = 29'b0_010110100101_100_1_001011010010;
      patterns[11565] = 29'b0_010110100101_101_0_100101101001;
      patterns[11566] = 29'b0_010110100101_110_0_010110100101;
      patterns[11567] = 29'b0_010110100101_111_0_010110100101;
      patterns[11568] = 29'b0_010110100110_000_0_010110100110;
      patterns[11569] = 29'b0_010110100110_001_0_100110010110;
      patterns[11570] = 29'b0_010110100110_010_0_101101001100;
      patterns[11571] = 29'b0_010110100110_011_1_011010011000;
      patterns[11572] = 29'b0_010110100110_100_0_001011010011;
      patterns[11573] = 29'b0_010110100110_101_1_000101101001;
      patterns[11574] = 29'b0_010110100110_110_0_010110100110;
      patterns[11575] = 29'b0_010110100110_111_0_010110100110;
      patterns[11576] = 29'b0_010110100111_000_0_010110100111;
      patterns[11577] = 29'b0_010110100111_001_0_100111010110;
      patterns[11578] = 29'b0_010110100111_010_0_101101001110;
      patterns[11579] = 29'b0_010110100111_011_1_011010011100;
      patterns[11580] = 29'b0_010110100111_100_1_001011010011;
      patterns[11581] = 29'b0_010110100111_101_1_100101101001;
      patterns[11582] = 29'b0_010110100111_110_0_010110100111;
      patterns[11583] = 29'b0_010110100111_111_0_010110100111;
      patterns[11584] = 29'b0_010110101000_000_0_010110101000;
      patterns[11585] = 29'b0_010110101000_001_0_101000010110;
      patterns[11586] = 29'b0_010110101000_010_0_101101010000;
      patterns[11587] = 29'b0_010110101000_011_1_011010100000;
      patterns[11588] = 29'b0_010110101000_100_0_001011010100;
      patterns[11589] = 29'b0_010110101000_101_0_000101101010;
      patterns[11590] = 29'b0_010110101000_110_0_010110101000;
      patterns[11591] = 29'b0_010110101000_111_0_010110101000;
      patterns[11592] = 29'b0_010110101001_000_0_010110101001;
      patterns[11593] = 29'b0_010110101001_001_0_101001010110;
      patterns[11594] = 29'b0_010110101001_010_0_101101010010;
      patterns[11595] = 29'b0_010110101001_011_1_011010100100;
      patterns[11596] = 29'b0_010110101001_100_1_001011010100;
      patterns[11597] = 29'b0_010110101001_101_0_100101101010;
      patterns[11598] = 29'b0_010110101001_110_0_010110101001;
      patterns[11599] = 29'b0_010110101001_111_0_010110101001;
      patterns[11600] = 29'b0_010110101010_000_0_010110101010;
      patterns[11601] = 29'b0_010110101010_001_0_101010010110;
      patterns[11602] = 29'b0_010110101010_010_0_101101010100;
      patterns[11603] = 29'b0_010110101010_011_1_011010101000;
      patterns[11604] = 29'b0_010110101010_100_0_001011010101;
      patterns[11605] = 29'b0_010110101010_101_1_000101101010;
      patterns[11606] = 29'b0_010110101010_110_0_010110101010;
      patterns[11607] = 29'b0_010110101010_111_0_010110101010;
      patterns[11608] = 29'b0_010110101011_000_0_010110101011;
      patterns[11609] = 29'b0_010110101011_001_0_101011010110;
      patterns[11610] = 29'b0_010110101011_010_0_101101010110;
      patterns[11611] = 29'b0_010110101011_011_1_011010101100;
      patterns[11612] = 29'b0_010110101011_100_1_001011010101;
      patterns[11613] = 29'b0_010110101011_101_1_100101101010;
      patterns[11614] = 29'b0_010110101011_110_0_010110101011;
      patterns[11615] = 29'b0_010110101011_111_0_010110101011;
      patterns[11616] = 29'b0_010110101100_000_0_010110101100;
      patterns[11617] = 29'b0_010110101100_001_0_101100010110;
      patterns[11618] = 29'b0_010110101100_010_0_101101011000;
      patterns[11619] = 29'b0_010110101100_011_1_011010110000;
      patterns[11620] = 29'b0_010110101100_100_0_001011010110;
      patterns[11621] = 29'b0_010110101100_101_0_000101101011;
      patterns[11622] = 29'b0_010110101100_110_0_010110101100;
      patterns[11623] = 29'b0_010110101100_111_0_010110101100;
      patterns[11624] = 29'b0_010110101101_000_0_010110101101;
      patterns[11625] = 29'b0_010110101101_001_0_101101010110;
      patterns[11626] = 29'b0_010110101101_010_0_101101011010;
      patterns[11627] = 29'b0_010110101101_011_1_011010110100;
      patterns[11628] = 29'b0_010110101101_100_1_001011010110;
      patterns[11629] = 29'b0_010110101101_101_0_100101101011;
      patterns[11630] = 29'b0_010110101101_110_0_010110101101;
      patterns[11631] = 29'b0_010110101101_111_0_010110101101;
      patterns[11632] = 29'b0_010110101110_000_0_010110101110;
      patterns[11633] = 29'b0_010110101110_001_0_101110010110;
      patterns[11634] = 29'b0_010110101110_010_0_101101011100;
      patterns[11635] = 29'b0_010110101110_011_1_011010111000;
      patterns[11636] = 29'b0_010110101110_100_0_001011010111;
      patterns[11637] = 29'b0_010110101110_101_1_000101101011;
      patterns[11638] = 29'b0_010110101110_110_0_010110101110;
      patterns[11639] = 29'b0_010110101110_111_0_010110101110;
      patterns[11640] = 29'b0_010110101111_000_0_010110101111;
      patterns[11641] = 29'b0_010110101111_001_0_101111010110;
      patterns[11642] = 29'b0_010110101111_010_0_101101011110;
      patterns[11643] = 29'b0_010110101111_011_1_011010111100;
      patterns[11644] = 29'b0_010110101111_100_1_001011010111;
      patterns[11645] = 29'b0_010110101111_101_1_100101101011;
      patterns[11646] = 29'b0_010110101111_110_0_010110101111;
      patterns[11647] = 29'b0_010110101111_111_0_010110101111;
      patterns[11648] = 29'b0_010110110000_000_0_010110110000;
      patterns[11649] = 29'b0_010110110000_001_0_110000010110;
      patterns[11650] = 29'b0_010110110000_010_0_101101100000;
      patterns[11651] = 29'b0_010110110000_011_1_011011000000;
      patterns[11652] = 29'b0_010110110000_100_0_001011011000;
      patterns[11653] = 29'b0_010110110000_101_0_000101101100;
      patterns[11654] = 29'b0_010110110000_110_0_010110110000;
      patterns[11655] = 29'b0_010110110000_111_0_010110110000;
      patterns[11656] = 29'b0_010110110001_000_0_010110110001;
      patterns[11657] = 29'b0_010110110001_001_0_110001010110;
      patterns[11658] = 29'b0_010110110001_010_0_101101100010;
      patterns[11659] = 29'b0_010110110001_011_1_011011000100;
      patterns[11660] = 29'b0_010110110001_100_1_001011011000;
      patterns[11661] = 29'b0_010110110001_101_0_100101101100;
      patterns[11662] = 29'b0_010110110001_110_0_010110110001;
      patterns[11663] = 29'b0_010110110001_111_0_010110110001;
      patterns[11664] = 29'b0_010110110010_000_0_010110110010;
      patterns[11665] = 29'b0_010110110010_001_0_110010010110;
      patterns[11666] = 29'b0_010110110010_010_0_101101100100;
      patterns[11667] = 29'b0_010110110010_011_1_011011001000;
      patterns[11668] = 29'b0_010110110010_100_0_001011011001;
      patterns[11669] = 29'b0_010110110010_101_1_000101101100;
      patterns[11670] = 29'b0_010110110010_110_0_010110110010;
      patterns[11671] = 29'b0_010110110010_111_0_010110110010;
      patterns[11672] = 29'b0_010110110011_000_0_010110110011;
      patterns[11673] = 29'b0_010110110011_001_0_110011010110;
      patterns[11674] = 29'b0_010110110011_010_0_101101100110;
      patterns[11675] = 29'b0_010110110011_011_1_011011001100;
      patterns[11676] = 29'b0_010110110011_100_1_001011011001;
      patterns[11677] = 29'b0_010110110011_101_1_100101101100;
      patterns[11678] = 29'b0_010110110011_110_0_010110110011;
      patterns[11679] = 29'b0_010110110011_111_0_010110110011;
      patterns[11680] = 29'b0_010110110100_000_0_010110110100;
      patterns[11681] = 29'b0_010110110100_001_0_110100010110;
      patterns[11682] = 29'b0_010110110100_010_0_101101101000;
      patterns[11683] = 29'b0_010110110100_011_1_011011010000;
      patterns[11684] = 29'b0_010110110100_100_0_001011011010;
      patterns[11685] = 29'b0_010110110100_101_0_000101101101;
      patterns[11686] = 29'b0_010110110100_110_0_010110110100;
      patterns[11687] = 29'b0_010110110100_111_0_010110110100;
      patterns[11688] = 29'b0_010110110101_000_0_010110110101;
      patterns[11689] = 29'b0_010110110101_001_0_110101010110;
      patterns[11690] = 29'b0_010110110101_010_0_101101101010;
      patterns[11691] = 29'b0_010110110101_011_1_011011010100;
      patterns[11692] = 29'b0_010110110101_100_1_001011011010;
      patterns[11693] = 29'b0_010110110101_101_0_100101101101;
      patterns[11694] = 29'b0_010110110101_110_0_010110110101;
      patterns[11695] = 29'b0_010110110101_111_0_010110110101;
      patterns[11696] = 29'b0_010110110110_000_0_010110110110;
      patterns[11697] = 29'b0_010110110110_001_0_110110010110;
      patterns[11698] = 29'b0_010110110110_010_0_101101101100;
      patterns[11699] = 29'b0_010110110110_011_1_011011011000;
      patterns[11700] = 29'b0_010110110110_100_0_001011011011;
      patterns[11701] = 29'b0_010110110110_101_1_000101101101;
      patterns[11702] = 29'b0_010110110110_110_0_010110110110;
      patterns[11703] = 29'b0_010110110110_111_0_010110110110;
      patterns[11704] = 29'b0_010110110111_000_0_010110110111;
      patterns[11705] = 29'b0_010110110111_001_0_110111010110;
      patterns[11706] = 29'b0_010110110111_010_0_101101101110;
      patterns[11707] = 29'b0_010110110111_011_1_011011011100;
      patterns[11708] = 29'b0_010110110111_100_1_001011011011;
      patterns[11709] = 29'b0_010110110111_101_1_100101101101;
      patterns[11710] = 29'b0_010110110111_110_0_010110110111;
      patterns[11711] = 29'b0_010110110111_111_0_010110110111;
      patterns[11712] = 29'b0_010110111000_000_0_010110111000;
      patterns[11713] = 29'b0_010110111000_001_0_111000010110;
      patterns[11714] = 29'b0_010110111000_010_0_101101110000;
      patterns[11715] = 29'b0_010110111000_011_1_011011100000;
      patterns[11716] = 29'b0_010110111000_100_0_001011011100;
      patterns[11717] = 29'b0_010110111000_101_0_000101101110;
      patterns[11718] = 29'b0_010110111000_110_0_010110111000;
      patterns[11719] = 29'b0_010110111000_111_0_010110111000;
      patterns[11720] = 29'b0_010110111001_000_0_010110111001;
      patterns[11721] = 29'b0_010110111001_001_0_111001010110;
      patterns[11722] = 29'b0_010110111001_010_0_101101110010;
      patterns[11723] = 29'b0_010110111001_011_1_011011100100;
      patterns[11724] = 29'b0_010110111001_100_1_001011011100;
      patterns[11725] = 29'b0_010110111001_101_0_100101101110;
      patterns[11726] = 29'b0_010110111001_110_0_010110111001;
      patterns[11727] = 29'b0_010110111001_111_0_010110111001;
      patterns[11728] = 29'b0_010110111010_000_0_010110111010;
      patterns[11729] = 29'b0_010110111010_001_0_111010010110;
      patterns[11730] = 29'b0_010110111010_010_0_101101110100;
      patterns[11731] = 29'b0_010110111010_011_1_011011101000;
      patterns[11732] = 29'b0_010110111010_100_0_001011011101;
      patterns[11733] = 29'b0_010110111010_101_1_000101101110;
      patterns[11734] = 29'b0_010110111010_110_0_010110111010;
      patterns[11735] = 29'b0_010110111010_111_0_010110111010;
      patterns[11736] = 29'b0_010110111011_000_0_010110111011;
      patterns[11737] = 29'b0_010110111011_001_0_111011010110;
      patterns[11738] = 29'b0_010110111011_010_0_101101110110;
      patterns[11739] = 29'b0_010110111011_011_1_011011101100;
      patterns[11740] = 29'b0_010110111011_100_1_001011011101;
      patterns[11741] = 29'b0_010110111011_101_1_100101101110;
      patterns[11742] = 29'b0_010110111011_110_0_010110111011;
      patterns[11743] = 29'b0_010110111011_111_0_010110111011;
      patterns[11744] = 29'b0_010110111100_000_0_010110111100;
      patterns[11745] = 29'b0_010110111100_001_0_111100010110;
      patterns[11746] = 29'b0_010110111100_010_0_101101111000;
      patterns[11747] = 29'b0_010110111100_011_1_011011110000;
      patterns[11748] = 29'b0_010110111100_100_0_001011011110;
      patterns[11749] = 29'b0_010110111100_101_0_000101101111;
      patterns[11750] = 29'b0_010110111100_110_0_010110111100;
      patterns[11751] = 29'b0_010110111100_111_0_010110111100;
      patterns[11752] = 29'b0_010110111101_000_0_010110111101;
      patterns[11753] = 29'b0_010110111101_001_0_111101010110;
      patterns[11754] = 29'b0_010110111101_010_0_101101111010;
      patterns[11755] = 29'b0_010110111101_011_1_011011110100;
      patterns[11756] = 29'b0_010110111101_100_1_001011011110;
      patterns[11757] = 29'b0_010110111101_101_0_100101101111;
      patterns[11758] = 29'b0_010110111101_110_0_010110111101;
      patterns[11759] = 29'b0_010110111101_111_0_010110111101;
      patterns[11760] = 29'b0_010110111110_000_0_010110111110;
      patterns[11761] = 29'b0_010110111110_001_0_111110010110;
      patterns[11762] = 29'b0_010110111110_010_0_101101111100;
      patterns[11763] = 29'b0_010110111110_011_1_011011111000;
      patterns[11764] = 29'b0_010110111110_100_0_001011011111;
      patterns[11765] = 29'b0_010110111110_101_1_000101101111;
      patterns[11766] = 29'b0_010110111110_110_0_010110111110;
      patterns[11767] = 29'b0_010110111110_111_0_010110111110;
      patterns[11768] = 29'b0_010110111111_000_0_010110111111;
      patterns[11769] = 29'b0_010110111111_001_0_111111010110;
      patterns[11770] = 29'b0_010110111111_010_0_101101111110;
      patterns[11771] = 29'b0_010110111111_011_1_011011111100;
      patterns[11772] = 29'b0_010110111111_100_1_001011011111;
      patterns[11773] = 29'b0_010110111111_101_1_100101101111;
      patterns[11774] = 29'b0_010110111111_110_0_010110111111;
      patterns[11775] = 29'b0_010110111111_111_0_010110111111;
      patterns[11776] = 29'b0_010111000000_000_0_010111000000;
      patterns[11777] = 29'b0_010111000000_001_0_000000010111;
      patterns[11778] = 29'b0_010111000000_010_0_101110000000;
      patterns[11779] = 29'b0_010111000000_011_1_011100000000;
      patterns[11780] = 29'b0_010111000000_100_0_001011100000;
      patterns[11781] = 29'b0_010111000000_101_0_000101110000;
      patterns[11782] = 29'b0_010111000000_110_0_010111000000;
      patterns[11783] = 29'b0_010111000000_111_0_010111000000;
      patterns[11784] = 29'b0_010111000001_000_0_010111000001;
      patterns[11785] = 29'b0_010111000001_001_0_000001010111;
      patterns[11786] = 29'b0_010111000001_010_0_101110000010;
      patterns[11787] = 29'b0_010111000001_011_1_011100000100;
      patterns[11788] = 29'b0_010111000001_100_1_001011100000;
      patterns[11789] = 29'b0_010111000001_101_0_100101110000;
      patterns[11790] = 29'b0_010111000001_110_0_010111000001;
      patterns[11791] = 29'b0_010111000001_111_0_010111000001;
      patterns[11792] = 29'b0_010111000010_000_0_010111000010;
      patterns[11793] = 29'b0_010111000010_001_0_000010010111;
      patterns[11794] = 29'b0_010111000010_010_0_101110000100;
      patterns[11795] = 29'b0_010111000010_011_1_011100001000;
      patterns[11796] = 29'b0_010111000010_100_0_001011100001;
      patterns[11797] = 29'b0_010111000010_101_1_000101110000;
      patterns[11798] = 29'b0_010111000010_110_0_010111000010;
      patterns[11799] = 29'b0_010111000010_111_0_010111000010;
      patterns[11800] = 29'b0_010111000011_000_0_010111000011;
      patterns[11801] = 29'b0_010111000011_001_0_000011010111;
      patterns[11802] = 29'b0_010111000011_010_0_101110000110;
      patterns[11803] = 29'b0_010111000011_011_1_011100001100;
      patterns[11804] = 29'b0_010111000011_100_1_001011100001;
      patterns[11805] = 29'b0_010111000011_101_1_100101110000;
      patterns[11806] = 29'b0_010111000011_110_0_010111000011;
      patterns[11807] = 29'b0_010111000011_111_0_010111000011;
      patterns[11808] = 29'b0_010111000100_000_0_010111000100;
      patterns[11809] = 29'b0_010111000100_001_0_000100010111;
      patterns[11810] = 29'b0_010111000100_010_0_101110001000;
      patterns[11811] = 29'b0_010111000100_011_1_011100010000;
      patterns[11812] = 29'b0_010111000100_100_0_001011100010;
      patterns[11813] = 29'b0_010111000100_101_0_000101110001;
      patterns[11814] = 29'b0_010111000100_110_0_010111000100;
      patterns[11815] = 29'b0_010111000100_111_0_010111000100;
      patterns[11816] = 29'b0_010111000101_000_0_010111000101;
      patterns[11817] = 29'b0_010111000101_001_0_000101010111;
      patterns[11818] = 29'b0_010111000101_010_0_101110001010;
      patterns[11819] = 29'b0_010111000101_011_1_011100010100;
      patterns[11820] = 29'b0_010111000101_100_1_001011100010;
      patterns[11821] = 29'b0_010111000101_101_0_100101110001;
      patterns[11822] = 29'b0_010111000101_110_0_010111000101;
      patterns[11823] = 29'b0_010111000101_111_0_010111000101;
      patterns[11824] = 29'b0_010111000110_000_0_010111000110;
      patterns[11825] = 29'b0_010111000110_001_0_000110010111;
      patterns[11826] = 29'b0_010111000110_010_0_101110001100;
      patterns[11827] = 29'b0_010111000110_011_1_011100011000;
      patterns[11828] = 29'b0_010111000110_100_0_001011100011;
      patterns[11829] = 29'b0_010111000110_101_1_000101110001;
      patterns[11830] = 29'b0_010111000110_110_0_010111000110;
      patterns[11831] = 29'b0_010111000110_111_0_010111000110;
      patterns[11832] = 29'b0_010111000111_000_0_010111000111;
      patterns[11833] = 29'b0_010111000111_001_0_000111010111;
      patterns[11834] = 29'b0_010111000111_010_0_101110001110;
      patterns[11835] = 29'b0_010111000111_011_1_011100011100;
      patterns[11836] = 29'b0_010111000111_100_1_001011100011;
      patterns[11837] = 29'b0_010111000111_101_1_100101110001;
      patterns[11838] = 29'b0_010111000111_110_0_010111000111;
      patterns[11839] = 29'b0_010111000111_111_0_010111000111;
      patterns[11840] = 29'b0_010111001000_000_0_010111001000;
      patterns[11841] = 29'b0_010111001000_001_0_001000010111;
      patterns[11842] = 29'b0_010111001000_010_0_101110010000;
      patterns[11843] = 29'b0_010111001000_011_1_011100100000;
      patterns[11844] = 29'b0_010111001000_100_0_001011100100;
      patterns[11845] = 29'b0_010111001000_101_0_000101110010;
      patterns[11846] = 29'b0_010111001000_110_0_010111001000;
      patterns[11847] = 29'b0_010111001000_111_0_010111001000;
      patterns[11848] = 29'b0_010111001001_000_0_010111001001;
      patterns[11849] = 29'b0_010111001001_001_0_001001010111;
      patterns[11850] = 29'b0_010111001001_010_0_101110010010;
      patterns[11851] = 29'b0_010111001001_011_1_011100100100;
      patterns[11852] = 29'b0_010111001001_100_1_001011100100;
      patterns[11853] = 29'b0_010111001001_101_0_100101110010;
      patterns[11854] = 29'b0_010111001001_110_0_010111001001;
      patterns[11855] = 29'b0_010111001001_111_0_010111001001;
      patterns[11856] = 29'b0_010111001010_000_0_010111001010;
      patterns[11857] = 29'b0_010111001010_001_0_001010010111;
      patterns[11858] = 29'b0_010111001010_010_0_101110010100;
      patterns[11859] = 29'b0_010111001010_011_1_011100101000;
      patterns[11860] = 29'b0_010111001010_100_0_001011100101;
      patterns[11861] = 29'b0_010111001010_101_1_000101110010;
      patterns[11862] = 29'b0_010111001010_110_0_010111001010;
      patterns[11863] = 29'b0_010111001010_111_0_010111001010;
      patterns[11864] = 29'b0_010111001011_000_0_010111001011;
      patterns[11865] = 29'b0_010111001011_001_0_001011010111;
      patterns[11866] = 29'b0_010111001011_010_0_101110010110;
      patterns[11867] = 29'b0_010111001011_011_1_011100101100;
      patterns[11868] = 29'b0_010111001011_100_1_001011100101;
      patterns[11869] = 29'b0_010111001011_101_1_100101110010;
      patterns[11870] = 29'b0_010111001011_110_0_010111001011;
      patterns[11871] = 29'b0_010111001011_111_0_010111001011;
      patterns[11872] = 29'b0_010111001100_000_0_010111001100;
      patterns[11873] = 29'b0_010111001100_001_0_001100010111;
      patterns[11874] = 29'b0_010111001100_010_0_101110011000;
      patterns[11875] = 29'b0_010111001100_011_1_011100110000;
      patterns[11876] = 29'b0_010111001100_100_0_001011100110;
      patterns[11877] = 29'b0_010111001100_101_0_000101110011;
      patterns[11878] = 29'b0_010111001100_110_0_010111001100;
      patterns[11879] = 29'b0_010111001100_111_0_010111001100;
      patterns[11880] = 29'b0_010111001101_000_0_010111001101;
      patterns[11881] = 29'b0_010111001101_001_0_001101010111;
      patterns[11882] = 29'b0_010111001101_010_0_101110011010;
      patterns[11883] = 29'b0_010111001101_011_1_011100110100;
      patterns[11884] = 29'b0_010111001101_100_1_001011100110;
      patterns[11885] = 29'b0_010111001101_101_0_100101110011;
      patterns[11886] = 29'b0_010111001101_110_0_010111001101;
      patterns[11887] = 29'b0_010111001101_111_0_010111001101;
      patterns[11888] = 29'b0_010111001110_000_0_010111001110;
      patterns[11889] = 29'b0_010111001110_001_0_001110010111;
      patterns[11890] = 29'b0_010111001110_010_0_101110011100;
      patterns[11891] = 29'b0_010111001110_011_1_011100111000;
      patterns[11892] = 29'b0_010111001110_100_0_001011100111;
      patterns[11893] = 29'b0_010111001110_101_1_000101110011;
      patterns[11894] = 29'b0_010111001110_110_0_010111001110;
      patterns[11895] = 29'b0_010111001110_111_0_010111001110;
      patterns[11896] = 29'b0_010111001111_000_0_010111001111;
      patterns[11897] = 29'b0_010111001111_001_0_001111010111;
      patterns[11898] = 29'b0_010111001111_010_0_101110011110;
      patterns[11899] = 29'b0_010111001111_011_1_011100111100;
      patterns[11900] = 29'b0_010111001111_100_1_001011100111;
      patterns[11901] = 29'b0_010111001111_101_1_100101110011;
      patterns[11902] = 29'b0_010111001111_110_0_010111001111;
      patterns[11903] = 29'b0_010111001111_111_0_010111001111;
      patterns[11904] = 29'b0_010111010000_000_0_010111010000;
      patterns[11905] = 29'b0_010111010000_001_0_010000010111;
      patterns[11906] = 29'b0_010111010000_010_0_101110100000;
      patterns[11907] = 29'b0_010111010000_011_1_011101000000;
      patterns[11908] = 29'b0_010111010000_100_0_001011101000;
      patterns[11909] = 29'b0_010111010000_101_0_000101110100;
      patterns[11910] = 29'b0_010111010000_110_0_010111010000;
      patterns[11911] = 29'b0_010111010000_111_0_010111010000;
      patterns[11912] = 29'b0_010111010001_000_0_010111010001;
      patterns[11913] = 29'b0_010111010001_001_0_010001010111;
      patterns[11914] = 29'b0_010111010001_010_0_101110100010;
      patterns[11915] = 29'b0_010111010001_011_1_011101000100;
      patterns[11916] = 29'b0_010111010001_100_1_001011101000;
      patterns[11917] = 29'b0_010111010001_101_0_100101110100;
      patterns[11918] = 29'b0_010111010001_110_0_010111010001;
      patterns[11919] = 29'b0_010111010001_111_0_010111010001;
      patterns[11920] = 29'b0_010111010010_000_0_010111010010;
      patterns[11921] = 29'b0_010111010010_001_0_010010010111;
      patterns[11922] = 29'b0_010111010010_010_0_101110100100;
      patterns[11923] = 29'b0_010111010010_011_1_011101001000;
      patterns[11924] = 29'b0_010111010010_100_0_001011101001;
      patterns[11925] = 29'b0_010111010010_101_1_000101110100;
      patterns[11926] = 29'b0_010111010010_110_0_010111010010;
      patterns[11927] = 29'b0_010111010010_111_0_010111010010;
      patterns[11928] = 29'b0_010111010011_000_0_010111010011;
      patterns[11929] = 29'b0_010111010011_001_0_010011010111;
      patterns[11930] = 29'b0_010111010011_010_0_101110100110;
      patterns[11931] = 29'b0_010111010011_011_1_011101001100;
      patterns[11932] = 29'b0_010111010011_100_1_001011101001;
      patterns[11933] = 29'b0_010111010011_101_1_100101110100;
      patterns[11934] = 29'b0_010111010011_110_0_010111010011;
      patterns[11935] = 29'b0_010111010011_111_0_010111010011;
      patterns[11936] = 29'b0_010111010100_000_0_010111010100;
      patterns[11937] = 29'b0_010111010100_001_0_010100010111;
      patterns[11938] = 29'b0_010111010100_010_0_101110101000;
      patterns[11939] = 29'b0_010111010100_011_1_011101010000;
      patterns[11940] = 29'b0_010111010100_100_0_001011101010;
      patterns[11941] = 29'b0_010111010100_101_0_000101110101;
      patterns[11942] = 29'b0_010111010100_110_0_010111010100;
      patterns[11943] = 29'b0_010111010100_111_0_010111010100;
      patterns[11944] = 29'b0_010111010101_000_0_010111010101;
      patterns[11945] = 29'b0_010111010101_001_0_010101010111;
      patterns[11946] = 29'b0_010111010101_010_0_101110101010;
      patterns[11947] = 29'b0_010111010101_011_1_011101010100;
      patterns[11948] = 29'b0_010111010101_100_1_001011101010;
      patterns[11949] = 29'b0_010111010101_101_0_100101110101;
      patterns[11950] = 29'b0_010111010101_110_0_010111010101;
      patterns[11951] = 29'b0_010111010101_111_0_010111010101;
      patterns[11952] = 29'b0_010111010110_000_0_010111010110;
      patterns[11953] = 29'b0_010111010110_001_0_010110010111;
      patterns[11954] = 29'b0_010111010110_010_0_101110101100;
      patterns[11955] = 29'b0_010111010110_011_1_011101011000;
      patterns[11956] = 29'b0_010111010110_100_0_001011101011;
      patterns[11957] = 29'b0_010111010110_101_1_000101110101;
      patterns[11958] = 29'b0_010111010110_110_0_010111010110;
      patterns[11959] = 29'b0_010111010110_111_0_010111010110;
      patterns[11960] = 29'b0_010111010111_000_0_010111010111;
      patterns[11961] = 29'b0_010111010111_001_0_010111010111;
      patterns[11962] = 29'b0_010111010111_010_0_101110101110;
      patterns[11963] = 29'b0_010111010111_011_1_011101011100;
      patterns[11964] = 29'b0_010111010111_100_1_001011101011;
      patterns[11965] = 29'b0_010111010111_101_1_100101110101;
      patterns[11966] = 29'b0_010111010111_110_0_010111010111;
      patterns[11967] = 29'b0_010111010111_111_0_010111010111;
      patterns[11968] = 29'b0_010111011000_000_0_010111011000;
      patterns[11969] = 29'b0_010111011000_001_0_011000010111;
      patterns[11970] = 29'b0_010111011000_010_0_101110110000;
      patterns[11971] = 29'b0_010111011000_011_1_011101100000;
      patterns[11972] = 29'b0_010111011000_100_0_001011101100;
      patterns[11973] = 29'b0_010111011000_101_0_000101110110;
      patterns[11974] = 29'b0_010111011000_110_0_010111011000;
      patterns[11975] = 29'b0_010111011000_111_0_010111011000;
      patterns[11976] = 29'b0_010111011001_000_0_010111011001;
      patterns[11977] = 29'b0_010111011001_001_0_011001010111;
      patterns[11978] = 29'b0_010111011001_010_0_101110110010;
      patterns[11979] = 29'b0_010111011001_011_1_011101100100;
      patterns[11980] = 29'b0_010111011001_100_1_001011101100;
      patterns[11981] = 29'b0_010111011001_101_0_100101110110;
      patterns[11982] = 29'b0_010111011001_110_0_010111011001;
      patterns[11983] = 29'b0_010111011001_111_0_010111011001;
      patterns[11984] = 29'b0_010111011010_000_0_010111011010;
      patterns[11985] = 29'b0_010111011010_001_0_011010010111;
      patterns[11986] = 29'b0_010111011010_010_0_101110110100;
      patterns[11987] = 29'b0_010111011010_011_1_011101101000;
      patterns[11988] = 29'b0_010111011010_100_0_001011101101;
      patterns[11989] = 29'b0_010111011010_101_1_000101110110;
      patterns[11990] = 29'b0_010111011010_110_0_010111011010;
      patterns[11991] = 29'b0_010111011010_111_0_010111011010;
      patterns[11992] = 29'b0_010111011011_000_0_010111011011;
      patterns[11993] = 29'b0_010111011011_001_0_011011010111;
      patterns[11994] = 29'b0_010111011011_010_0_101110110110;
      patterns[11995] = 29'b0_010111011011_011_1_011101101100;
      patterns[11996] = 29'b0_010111011011_100_1_001011101101;
      patterns[11997] = 29'b0_010111011011_101_1_100101110110;
      patterns[11998] = 29'b0_010111011011_110_0_010111011011;
      patterns[11999] = 29'b0_010111011011_111_0_010111011011;
      patterns[12000] = 29'b0_010111011100_000_0_010111011100;
      patterns[12001] = 29'b0_010111011100_001_0_011100010111;
      patterns[12002] = 29'b0_010111011100_010_0_101110111000;
      patterns[12003] = 29'b0_010111011100_011_1_011101110000;
      patterns[12004] = 29'b0_010111011100_100_0_001011101110;
      patterns[12005] = 29'b0_010111011100_101_0_000101110111;
      patterns[12006] = 29'b0_010111011100_110_0_010111011100;
      patterns[12007] = 29'b0_010111011100_111_0_010111011100;
      patterns[12008] = 29'b0_010111011101_000_0_010111011101;
      patterns[12009] = 29'b0_010111011101_001_0_011101010111;
      patterns[12010] = 29'b0_010111011101_010_0_101110111010;
      patterns[12011] = 29'b0_010111011101_011_1_011101110100;
      patterns[12012] = 29'b0_010111011101_100_1_001011101110;
      patterns[12013] = 29'b0_010111011101_101_0_100101110111;
      patterns[12014] = 29'b0_010111011101_110_0_010111011101;
      patterns[12015] = 29'b0_010111011101_111_0_010111011101;
      patterns[12016] = 29'b0_010111011110_000_0_010111011110;
      patterns[12017] = 29'b0_010111011110_001_0_011110010111;
      patterns[12018] = 29'b0_010111011110_010_0_101110111100;
      patterns[12019] = 29'b0_010111011110_011_1_011101111000;
      patterns[12020] = 29'b0_010111011110_100_0_001011101111;
      patterns[12021] = 29'b0_010111011110_101_1_000101110111;
      patterns[12022] = 29'b0_010111011110_110_0_010111011110;
      patterns[12023] = 29'b0_010111011110_111_0_010111011110;
      patterns[12024] = 29'b0_010111011111_000_0_010111011111;
      patterns[12025] = 29'b0_010111011111_001_0_011111010111;
      patterns[12026] = 29'b0_010111011111_010_0_101110111110;
      patterns[12027] = 29'b0_010111011111_011_1_011101111100;
      patterns[12028] = 29'b0_010111011111_100_1_001011101111;
      patterns[12029] = 29'b0_010111011111_101_1_100101110111;
      patterns[12030] = 29'b0_010111011111_110_0_010111011111;
      patterns[12031] = 29'b0_010111011111_111_0_010111011111;
      patterns[12032] = 29'b0_010111100000_000_0_010111100000;
      patterns[12033] = 29'b0_010111100000_001_0_100000010111;
      patterns[12034] = 29'b0_010111100000_010_0_101111000000;
      patterns[12035] = 29'b0_010111100000_011_1_011110000000;
      patterns[12036] = 29'b0_010111100000_100_0_001011110000;
      patterns[12037] = 29'b0_010111100000_101_0_000101111000;
      patterns[12038] = 29'b0_010111100000_110_0_010111100000;
      patterns[12039] = 29'b0_010111100000_111_0_010111100000;
      patterns[12040] = 29'b0_010111100001_000_0_010111100001;
      patterns[12041] = 29'b0_010111100001_001_0_100001010111;
      patterns[12042] = 29'b0_010111100001_010_0_101111000010;
      patterns[12043] = 29'b0_010111100001_011_1_011110000100;
      patterns[12044] = 29'b0_010111100001_100_1_001011110000;
      patterns[12045] = 29'b0_010111100001_101_0_100101111000;
      patterns[12046] = 29'b0_010111100001_110_0_010111100001;
      patterns[12047] = 29'b0_010111100001_111_0_010111100001;
      patterns[12048] = 29'b0_010111100010_000_0_010111100010;
      patterns[12049] = 29'b0_010111100010_001_0_100010010111;
      patterns[12050] = 29'b0_010111100010_010_0_101111000100;
      patterns[12051] = 29'b0_010111100010_011_1_011110001000;
      patterns[12052] = 29'b0_010111100010_100_0_001011110001;
      patterns[12053] = 29'b0_010111100010_101_1_000101111000;
      patterns[12054] = 29'b0_010111100010_110_0_010111100010;
      patterns[12055] = 29'b0_010111100010_111_0_010111100010;
      patterns[12056] = 29'b0_010111100011_000_0_010111100011;
      patterns[12057] = 29'b0_010111100011_001_0_100011010111;
      patterns[12058] = 29'b0_010111100011_010_0_101111000110;
      patterns[12059] = 29'b0_010111100011_011_1_011110001100;
      patterns[12060] = 29'b0_010111100011_100_1_001011110001;
      patterns[12061] = 29'b0_010111100011_101_1_100101111000;
      patterns[12062] = 29'b0_010111100011_110_0_010111100011;
      patterns[12063] = 29'b0_010111100011_111_0_010111100011;
      patterns[12064] = 29'b0_010111100100_000_0_010111100100;
      patterns[12065] = 29'b0_010111100100_001_0_100100010111;
      patterns[12066] = 29'b0_010111100100_010_0_101111001000;
      patterns[12067] = 29'b0_010111100100_011_1_011110010000;
      patterns[12068] = 29'b0_010111100100_100_0_001011110010;
      patterns[12069] = 29'b0_010111100100_101_0_000101111001;
      patterns[12070] = 29'b0_010111100100_110_0_010111100100;
      patterns[12071] = 29'b0_010111100100_111_0_010111100100;
      patterns[12072] = 29'b0_010111100101_000_0_010111100101;
      patterns[12073] = 29'b0_010111100101_001_0_100101010111;
      patterns[12074] = 29'b0_010111100101_010_0_101111001010;
      patterns[12075] = 29'b0_010111100101_011_1_011110010100;
      patterns[12076] = 29'b0_010111100101_100_1_001011110010;
      patterns[12077] = 29'b0_010111100101_101_0_100101111001;
      patterns[12078] = 29'b0_010111100101_110_0_010111100101;
      patterns[12079] = 29'b0_010111100101_111_0_010111100101;
      patterns[12080] = 29'b0_010111100110_000_0_010111100110;
      patterns[12081] = 29'b0_010111100110_001_0_100110010111;
      patterns[12082] = 29'b0_010111100110_010_0_101111001100;
      patterns[12083] = 29'b0_010111100110_011_1_011110011000;
      patterns[12084] = 29'b0_010111100110_100_0_001011110011;
      patterns[12085] = 29'b0_010111100110_101_1_000101111001;
      patterns[12086] = 29'b0_010111100110_110_0_010111100110;
      patterns[12087] = 29'b0_010111100110_111_0_010111100110;
      patterns[12088] = 29'b0_010111100111_000_0_010111100111;
      patterns[12089] = 29'b0_010111100111_001_0_100111010111;
      patterns[12090] = 29'b0_010111100111_010_0_101111001110;
      patterns[12091] = 29'b0_010111100111_011_1_011110011100;
      patterns[12092] = 29'b0_010111100111_100_1_001011110011;
      patterns[12093] = 29'b0_010111100111_101_1_100101111001;
      patterns[12094] = 29'b0_010111100111_110_0_010111100111;
      patterns[12095] = 29'b0_010111100111_111_0_010111100111;
      patterns[12096] = 29'b0_010111101000_000_0_010111101000;
      patterns[12097] = 29'b0_010111101000_001_0_101000010111;
      patterns[12098] = 29'b0_010111101000_010_0_101111010000;
      patterns[12099] = 29'b0_010111101000_011_1_011110100000;
      patterns[12100] = 29'b0_010111101000_100_0_001011110100;
      patterns[12101] = 29'b0_010111101000_101_0_000101111010;
      patterns[12102] = 29'b0_010111101000_110_0_010111101000;
      patterns[12103] = 29'b0_010111101000_111_0_010111101000;
      patterns[12104] = 29'b0_010111101001_000_0_010111101001;
      patterns[12105] = 29'b0_010111101001_001_0_101001010111;
      patterns[12106] = 29'b0_010111101001_010_0_101111010010;
      patterns[12107] = 29'b0_010111101001_011_1_011110100100;
      patterns[12108] = 29'b0_010111101001_100_1_001011110100;
      patterns[12109] = 29'b0_010111101001_101_0_100101111010;
      patterns[12110] = 29'b0_010111101001_110_0_010111101001;
      patterns[12111] = 29'b0_010111101001_111_0_010111101001;
      patterns[12112] = 29'b0_010111101010_000_0_010111101010;
      patterns[12113] = 29'b0_010111101010_001_0_101010010111;
      patterns[12114] = 29'b0_010111101010_010_0_101111010100;
      patterns[12115] = 29'b0_010111101010_011_1_011110101000;
      patterns[12116] = 29'b0_010111101010_100_0_001011110101;
      patterns[12117] = 29'b0_010111101010_101_1_000101111010;
      patterns[12118] = 29'b0_010111101010_110_0_010111101010;
      patterns[12119] = 29'b0_010111101010_111_0_010111101010;
      patterns[12120] = 29'b0_010111101011_000_0_010111101011;
      patterns[12121] = 29'b0_010111101011_001_0_101011010111;
      patterns[12122] = 29'b0_010111101011_010_0_101111010110;
      patterns[12123] = 29'b0_010111101011_011_1_011110101100;
      patterns[12124] = 29'b0_010111101011_100_1_001011110101;
      patterns[12125] = 29'b0_010111101011_101_1_100101111010;
      patterns[12126] = 29'b0_010111101011_110_0_010111101011;
      patterns[12127] = 29'b0_010111101011_111_0_010111101011;
      patterns[12128] = 29'b0_010111101100_000_0_010111101100;
      patterns[12129] = 29'b0_010111101100_001_0_101100010111;
      patterns[12130] = 29'b0_010111101100_010_0_101111011000;
      patterns[12131] = 29'b0_010111101100_011_1_011110110000;
      patterns[12132] = 29'b0_010111101100_100_0_001011110110;
      patterns[12133] = 29'b0_010111101100_101_0_000101111011;
      patterns[12134] = 29'b0_010111101100_110_0_010111101100;
      patterns[12135] = 29'b0_010111101100_111_0_010111101100;
      patterns[12136] = 29'b0_010111101101_000_0_010111101101;
      patterns[12137] = 29'b0_010111101101_001_0_101101010111;
      patterns[12138] = 29'b0_010111101101_010_0_101111011010;
      patterns[12139] = 29'b0_010111101101_011_1_011110110100;
      patterns[12140] = 29'b0_010111101101_100_1_001011110110;
      patterns[12141] = 29'b0_010111101101_101_0_100101111011;
      patterns[12142] = 29'b0_010111101101_110_0_010111101101;
      patterns[12143] = 29'b0_010111101101_111_0_010111101101;
      patterns[12144] = 29'b0_010111101110_000_0_010111101110;
      patterns[12145] = 29'b0_010111101110_001_0_101110010111;
      patterns[12146] = 29'b0_010111101110_010_0_101111011100;
      patterns[12147] = 29'b0_010111101110_011_1_011110111000;
      patterns[12148] = 29'b0_010111101110_100_0_001011110111;
      patterns[12149] = 29'b0_010111101110_101_1_000101111011;
      patterns[12150] = 29'b0_010111101110_110_0_010111101110;
      patterns[12151] = 29'b0_010111101110_111_0_010111101110;
      patterns[12152] = 29'b0_010111101111_000_0_010111101111;
      patterns[12153] = 29'b0_010111101111_001_0_101111010111;
      patterns[12154] = 29'b0_010111101111_010_0_101111011110;
      patterns[12155] = 29'b0_010111101111_011_1_011110111100;
      patterns[12156] = 29'b0_010111101111_100_1_001011110111;
      patterns[12157] = 29'b0_010111101111_101_1_100101111011;
      patterns[12158] = 29'b0_010111101111_110_0_010111101111;
      patterns[12159] = 29'b0_010111101111_111_0_010111101111;
      patterns[12160] = 29'b0_010111110000_000_0_010111110000;
      patterns[12161] = 29'b0_010111110000_001_0_110000010111;
      patterns[12162] = 29'b0_010111110000_010_0_101111100000;
      patterns[12163] = 29'b0_010111110000_011_1_011111000000;
      patterns[12164] = 29'b0_010111110000_100_0_001011111000;
      patterns[12165] = 29'b0_010111110000_101_0_000101111100;
      patterns[12166] = 29'b0_010111110000_110_0_010111110000;
      patterns[12167] = 29'b0_010111110000_111_0_010111110000;
      patterns[12168] = 29'b0_010111110001_000_0_010111110001;
      patterns[12169] = 29'b0_010111110001_001_0_110001010111;
      patterns[12170] = 29'b0_010111110001_010_0_101111100010;
      patterns[12171] = 29'b0_010111110001_011_1_011111000100;
      patterns[12172] = 29'b0_010111110001_100_1_001011111000;
      patterns[12173] = 29'b0_010111110001_101_0_100101111100;
      patterns[12174] = 29'b0_010111110001_110_0_010111110001;
      patterns[12175] = 29'b0_010111110001_111_0_010111110001;
      patterns[12176] = 29'b0_010111110010_000_0_010111110010;
      patterns[12177] = 29'b0_010111110010_001_0_110010010111;
      patterns[12178] = 29'b0_010111110010_010_0_101111100100;
      patterns[12179] = 29'b0_010111110010_011_1_011111001000;
      patterns[12180] = 29'b0_010111110010_100_0_001011111001;
      patterns[12181] = 29'b0_010111110010_101_1_000101111100;
      patterns[12182] = 29'b0_010111110010_110_0_010111110010;
      patterns[12183] = 29'b0_010111110010_111_0_010111110010;
      patterns[12184] = 29'b0_010111110011_000_0_010111110011;
      patterns[12185] = 29'b0_010111110011_001_0_110011010111;
      patterns[12186] = 29'b0_010111110011_010_0_101111100110;
      patterns[12187] = 29'b0_010111110011_011_1_011111001100;
      patterns[12188] = 29'b0_010111110011_100_1_001011111001;
      patterns[12189] = 29'b0_010111110011_101_1_100101111100;
      patterns[12190] = 29'b0_010111110011_110_0_010111110011;
      patterns[12191] = 29'b0_010111110011_111_0_010111110011;
      patterns[12192] = 29'b0_010111110100_000_0_010111110100;
      patterns[12193] = 29'b0_010111110100_001_0_110100010111;
      patterns[12194] = 29'b0_010111110100_010_0_101111101000;
      patterns[12195] = 29'b0_010111110100_011_1_011111010000;
      patterns[12196] = 29'b0_010111110100_100_0_001011111010;
      patterns[12197] = 29'b0_010111110100_101_0_000101111101;
      patterns[12198] = 29'b0_010111110100_110_0_010111110100;
      patterns[12199] = 29'b0_010111110100_111_0_010111110100;
      patterns[12200] = 29'b0_010111110101_000_0_010111110101;
      patterns[12201] = 29'b0_010111110101_001_0_110101010111;
      patterns[12202] = 29'b0_010111110101_010_0_101111101010;
      patterns[12203] = 29'b0_010111110101_011_1_011111010100;
      patterns[12204] = 29'b0_010111110101_100_1_001011111010;
      patterns[12205] = 29'b0_010111110101_101_0_100101111101;
      patterns[12206] = 29'b0_010111110101_110_0_010111110101;
      patterns[12207] = 29'b0_010111110101_111_0_010111110101;
      patterns[12208] = 29'b0_010111110110_000_0_010111110110;
      patterns[12209] = 29'b0_010111110110_001_0_110110010111;
      patterns[12210] = 29'b0_010111110110_010_0_101111101100;
      patterns[12211] = 29'b0_010111110110_011_1_011111011000;
      patterns[12212] = 29'b0_010111110110_100_0_001011111011;
      patterns[12213] = 29'b0_010111110110_101_1_000101111101;
      patterns[12214] = 29'b0_010111110110_110_0_010111110110;
      patterns[12215] = 29'b0_010111110110_111_0_010111110110;
      patterns[12216] = 29'b0_010111110111_000_0_010111110111;
      patterns[12217] = 29'b0_010111110111_001_0_110111010111;
      patterns[12218] = 29'b0_010111110111_010_0_101111101110;
      patterns[12219] = 29'b0_010111110111_011_1_011111011100;
      patterns[12220] = 29'b0_010111110111_100_1_001011111011;
      patterns[12221] = 29'b0_010111110111_101_1_100101111101;
      patterns[12222] = 29'b0_010111110111_110_0_010111110111;
      patterns[12223] = 29'b0_010111110111_111_0_010111110111;
      patterns[12224] = 29'b0_010111111000_000_0_010111111000;
      patterns[12225] = 29'b0_010111111000_001_0_111000010111;
      patterns[12226] = 29'b0_010111111000_010_0_101111110000;
      patterns[12227] = 29'b0_010111111000_011_1_011111100000;
      patterns[12228] = 29'b0_010111111000_100_0_001011111100;
      patterns[12229] = 29'b0_010111111000_101_0_000101111110;
      patterns[12230] = 29'b0_010111111000_110_0_010111111000;
      patterns[12231] = 29'b0_010111111000_111_0_010111111000;
      patterns[12232] = 29'b0_010111111001_000_0_010111111001;
      patterns[12233] = 29'b0_010111111001_001_0_111001010111;
      patterns[12234] = 29'b0_010111111001_010_0_101111110010;
      patterns[12235] = 29'b0_010111111001_011_1_011111100100;
      patterns[12236] = 29'b0_010111111001_100_1_001011111100;
      patterns[12237] = 29'b0_010111111001_101_0_100101111110;
      patterns[12238] = 29'b0_010111111001_110_0_010111111001;
      patterns[12239] = 29'b0_010111111001_111_0_010111111001;
      patterns[12240] = 29'b0_010111111010_000_0_010111111010;
      patterns[12241] = 29'b0_010111111010_001_0_111010010111;
      patterns[12242] = 29'b0_010111111010_010_0_101111110100;
      patterns[12243] = 29'b0_010111111010_011_1_011111101000;
      patterns[12244] = 29'b0_010111111010_100_0_001011111101;
      patterns[12245] = 29'b0_010111111010_101_1_000101111110;
      patterns[12246] = 29'b0_010111111010_110_0_010111111010;
      patterns[12247] = 29'b0_010111111010_111_0_010111111010;
      patterns[12248] = 29'b0_010111111011_000_0_010111111011;
      patterns[12249] = 29'b0_010111111011_001_0_111011010111;
      patterns[12250] = 29'b0_010111111011_010_0_101111110110;
      patterns[12251] = 29'b0_010111111011_011_1_011111101100;
      patterns[12252] = 29'b0_010111111011_100_1_001011111101;
      patterns[12253] = 29'b0_010111111011_101_1_100101111110;
      patterns[12254] = 29'b0_010111111011_110_0_010111111011;
      patterns[12255] = 29'b0_010111111011_111_0_010111111011;
      patterns[12256] = 29'b0_010111111100_000_0_010111111100;
      patterns[12257] = 29'b0_010111111100_001_0_111100010111;
      patterns[12258] = 29'b0_010111111100_010_0_101111111000;
      patterns[12259] = 29'b0_010111111100_011_1_011111110000;
      patterns[12260] = 29'b0_010111111100_100_0_001011111110;
      patterns[12261] = 29'b0_010111111100_101_0_000101111111;
      patterns[12262] = 29'b0_010111111100_110_0_010111111100;
      patterns[12263] = 29'b0_010111111100_111_0_010111111100;
      patterns[12264] = 29'b0_010111111101_000_0_010111111101;
      patterns[12265] = 29'b0_010111111101_001_0_111101010111;
      patterns[12266] = 29'b0_010111111101_010_0_101111111010;
      patterns[12267] = 29'b0_010111111101_011_1_011111110100;
      patterns[12268] = 29'b0_010111111101_100_1_001011111110;
      patterns[12269] = 29'b0_010111111101_101_0_100101111111;
      patterns[12270] = 29'b0_010111111101_110_0_010111111101;
      patterns[12271] = 29'b0_010111111101_111_0_010111111101;
      patterns[12272] = 29'b0_010111111110_000_0_010111111110;
      patterns[12273] = 29'b0_010111111110_001_0_111110010111;
      patterns[12274] = 29'b0_010111111110_010_0_101111111100;
      patterns[12275] = 29'b0_010111111110_011_1_011111111000;
      patterns[12276] = 29'b0_010111111110_100_0_001011111111;
      patterns[12277] = 29'b0_010111111110_101_1_000101111111;
      patterns[12278] = 29'b0_010111111110_110_0_010111111110;
      patterns[12279] = 29'b0_010111111110_111_0_010111111110;
      patterns[12280] = 29'b0_010111111111_000_0_010111111111;
      patterns[12281] = 29'b0_010111111111_001_0_111111010111;
      patterns[12282] = 29'b0_010111111111_010_0_101111111110;
      patterns[12283] = 29'b0_010111111111_011_1_011111111100;
      patterns[12284] = 29'b0_010111111111_100_1_001011111111;
      patterns[12285] = 29'b0_010111111111_101_1_100101111111;
      patterns[12286] = 29'b0_010111111111_110_0_010111111111;
      patterns[12287] = 29'b0_010111111111_111_0_010111111111;
      patterns[12288] = 29'b0_011000000000_000_0_011000000000;
      patterns[12289] = 29'b0_011000000000_001_0_000000011000;
      patterns[12290] = 29'b0_011000000000_010_0_110000000000;
      patterns[12291] = 29'b0_011000000000_011_1_100000000000;
      patterns[12292] = 29'b0_011000000000_100_0_001100000000;
      patterns[12293] = 29'b0_011000000000_101_0_000110000000;
      patterns[12294] = 29'b0_011000000000_110_0_011000000000;
      patterns[12295] = 29'b0_011000000000_111_0_011000000000;
      patterns[12296] = 29'b0_011000000001_000_0_011000000001;
      patterns[12297] = 29'b0_011000000001_001_0_000001011000;
      patterns[12298] = 29'b0_011000000001_010_0_110000000010;
      patterns[12299] = 29'b0_011000000001_011_1_100000000100;
      patterns[12300] = 29'b0_011000000001_100_1_001100000000;
      patterns[12301] = 29'b0_011000000001_101_0_100110000000;
      patterns[12302] = 29'b0_011000000001_110_0_011000000001;
      patterns[12303] = 29'b0_011000000001_111_0_011000000001;
      patterns[12304] = 29'b0_011000000010_000_0_011000000010;
      patterns[12305] = 29'b0_011000000010_001_0_000010011000;
      patterns[12306] = 29'b0_011000000010_010_0_110000000100;
      patterns[12307] = 29'b0_011000000010_011_1_100000001000;
      patterns[12308] = 29'b0_011000000010_100_0_001100000001;
      patterns[12309] = 29'b0_011000000010_101_1_000110000000;
      patterns[12310] = 29'b0_011000000010_110_0_011000000010;
      patterns[12311] = 29'b0_011000000010_111_0_011000000010;
      patterns[12312] = 29'b0_011000000011_000_0_011000000011;
      patterns[12313] = 29'b0_011000000011_001_0_000011011000;
      patterns[12314] = 29'b0_011000000011_010_0_110000000110;
      patterns[12315] = 29'b0_011000000011_011_1_100000001100;
      patterns[12316] = 29'b0_011000000011_100_1_001100000001;
      patterns[12317] = 29'b0_011000000011_101_1_100110000000;
      patterns[12318] = 29'b0_011000000011_110_0_011000000011;
      patterns[12319] = 29'b0_011000000011_111_0_011000000011;
      patterns[12320] = 29'b0_011000000100_000_0_011000000100;
      patterns[12321] = 29'b0_011000000100_001_0_000100011000;
      patterns[12322] = 29'b0_011000000100_010_0_110000001000;
      patterns[12323] = 29'b0_011000000100_011_1_100000010000;
      patterns[12324] = 29'b0_011000000100_100_0_001100000010;
      patterns[12325] = 29'b0_011000000100_101_0_000110000001;
      patterns[12326] = 29'b0_011000000100_110_0_011000000100;
      patterns[12327] = 29'b0_011000000100_111_0_011000000100;
      patterns[12328] = 29'b0_011000000101_000_0_011000000101;
      patterns[12329] = 29'b0_011000000101_001_0_000101011000;
      patterns[12330] = 29'b0_011000000101_010_0_110000001010;
      patterns[12331] = 29'b0_011000000101_011_1_100000010100;
      patterns[12332] = 29'b0_011000000101_100_1_001100000010;
      patterns[12333] = 29'b0_011000000101_101_0_100110000001;
      patterns[12334] = 29'b0_011000000101_110_0_011000000101;
      patterns[12335] = 29'b0_011000000101_111_0_011000000101;
      patterns[12336] = 29'b0_011000000110_000_0_011000000110;
      patterns[12337] = 29'b0_011000000110_001_0_000110011000;
      patterns[12338] = 29'b0_011000000110_010_0_110000001100;
      patterns[12339] = 29'b0_011000000110_011_1_100000011000;
      patterns[12340] = 29'b0_011000000110_100_0_001100000011;
      patterns[12341] = 29'b0_011000000110_101_1_000110000001;
      patterns[12342] = 29'b0_011000000110_110_0_011000000110;
      patterns[12343] = 29'b0_011000000110_111_0_011000000110;
      patterns[12344] = 29'b0_011000000111_000_0_011000000111;
      patterns[12345] = 29'b0_011000000111_001_0_000111011000;
      patterns[12346] = 29'b0_011000000111_010_0_110000001110;
      patterns[12347] = 29'b0_011000000111_011_1_100000011100;
      patterns[12348] = 29'b0_011000000111_100_1_001100000011;
      patterns[12349] = 29'b0_011000000111_101_1_100110000001;
      patterns[12350] = 29'b0_011000000111_110_0_011000000111;
      patterns[12351] = 29'b0_011000000111_111_0_011000000111;
      patterns[12352] = 29'b0_011000001000_000_0_011000001000;
      patterns[12353] = 29'b0_011000001000_001_0_001000011000;
      patterns[12354] = 29'b0_011000001000_010_0_110000010000;
      patterns[12355] = 29'b0_011000001000_011_1_100000100000;
      patterns[12356] = 29'b0_011000001000_100_0_001100000100;
      patterns[12357] = 29'b0_011000001000_101_0_000110000010;
      patterns[12358] = 29'b0_011000001000_110_0_011000001000;
      patterns[12359] = 29'b0_011000001000_111_0_011000001000;
      patterns[12360] = 29'b0_011000001001_000_0_011000001001;
      patterns[12361] = 29'b0_011000001001_001_0_001001011000;
      patterns[12362] = 29'b0_011000001001_010_0_110000010010;
      patterns[12363] = 29'b0_011000001001_011_1_100000100100;
      patterns[12364] = 29'b0_011000001001_100_1_001100000100;
      patterns[12365] = 29'b0_011000001001_101_0_100110000010;
      patterns[12366] = 29'b0_011000001001_110_0_011000001001;
      patterns[12367] = 29'b0_011000001001_111_0_011000001001;
      patterns[12368] = 29'b0_011000001010_000_0_011000001010;
      patterns[12369] = 29'b0_011000001010_001_0_001010011000;
      patterns[12370] = 29'b0_011000001010_010_0_110000010100;
      patterns[12371] = 29'b0_011000001010_011_1_100000101000;
      patterns[12372] = 29'b0_011000001010_100_0_001100000101;
      patterns[12373] = 29'b0_011000001010_101_1_000110000010;
      patterns[12374] = 29'b0_011000001010_110_0_011000001010;
      patterns[12375] = 29'b0_011000001010_111_0_011000001010;
      patterns[12376] = 29'b0_011000001011_000_0_011000001011;
      patterns[12377] = 29'b0_011000001011_001_0_001011011000;
      patterns[12378] = 29'b0_011000001011_010_0_110000010110;
      patterns[12379] = 29'b0_011000001011_011_1_100000101100;
      patterns[12380] = 29'b0_011000001011_100_1_001100000101;
      patterns[12381] = 29'b0_011000001011_101_1_100110000010;
      patterns[12382] = 29'b0_011000001011_110_0_011000001011;
      patterns[12383] = 29'b0_011000001011_111_0_011000001011;
      patterns[12384] = 29'b0_011000001100_000_0_011000001100;
      patterns[12385] = 29'b0_011000001100_001_0_001100011000;
      patterns[12386] = 29'b0_011000001100_010_0_110000011000;
      patterns[12387] = 29'b0_011000001100_011_1_100000110000;
      patterns[12388] = 29'b0_011000001100_100_0_001100000110;
      patterns[12389] = 29'b0_011000001100_101_0_000110000011;
      patterns[12390] = 29'b0_011000001100_110_0_011000001100;
      patterns[12391] = 29'b0_011000001100_111_0_011000001100;
      patterns[12392] = 29'b0_011000001101_000_0_011000001101;
      patterns[12393] = 29'b0_011000001101_001_0_001101011000;
      patterns[12394] = 29'b0_011000001101_010_0_110000011010;
      patterns[12395] = 29'b0_011000001101_011_1_100000110100;
      patterns[12396] = 29'b0_011000001101_100_1_001100000110;
      patterns[12397] = 29'b0_011000001101_101_0_100110000011;
      patterns[12398] = 29'b0_011000001101_110_0_011000001101;
      patterns[12399] = 29'b0_011000001101_111_0_011000001101;
      patterns[12400] = 29'b0_011000001110_000_0_011000001110;
      patterns[12401] = 29'b0_011000001110_001_0_001110011000;
      patterns[12402] = 29'b0_011000001110_010_0_110000011100;
      patterns[12403] = 29'b0_011000001110_011_1_100000111000;
      patterns[12404] = 29'b0_011000001110_100_0_001100000111;
      patterns[12405] = 29'b0_011000001110_101_1_000110000011;
      patterns[12406] = 29'b0_011000001110_110_0_011000001110;
      patterns[12407] = 29'b0_011000001110_111_0_011000001110;
      patterns[12408] = 29'b0_011000001111_000_0_011000001111;
      patterns[12409] = 29'b0_011000001111_001_0_001111011000;
      patterns[12410] = 29'b0_011000001111_010_0_110000011110;
      patterns[12411] = 29'b0_011000001111_011_1_100000111100;
      patterns[12412] = 29'b0_011000001111_100_1_001100000111;
      patterns[12413] = 29'b0_011000001111_101_1_100110000011;
      patterns[12414] = 29'b0_011000001111_110_0_011000001111;
      patterns[12415] = 29'b0_011000001111_111_0_011000001111;
      patterns[12416] = 29'b0_011000010000_000_0_011000010000;
      patterns[12417] = 29'b0_011000010000_001_0_010000011000;
      patterns[12418] = 29'b0_011000010000_010_0_110000100000;
      patterns[12419] = 29'b0_011000010000_011_1_100001000000;
      patterns[12420] = 29'b0_011000010000_100_0_001100001000;
      patterns[12421] = 29'b0_011000010000_101_0_000110000100;
      patterns[12422] = 29'b0_011000010000_110_0_011000010000;
      patterns[12423] = 29'b0_011000010000_111_0_011000010000;
      patterns[12424] = 29'b0_011000010001_000_0_011000010001;
      patterns[12425] = 29'b0_011000010001_001_0_010001011000;
      patterns[12426] = 29'b0_011000010001_010_0_110000100010;
      patterns[12427] = 29'b0_011000010001_011_1_100001000100;
      patterns[12428] = 29'b0_011000010001_100_1_001100001000;
      patterns[12429] = 29'b0_011000010001_101_0_100110000100;
      patterns[12430] = 29'b0_011000010001_110_0_011000010001;
      patterns[12431] = 29'b0_011000010001_111_0_011000010001;
      patterns[12432] = 29'b0_011000010010_000_0_011000010010;
      patterns[12433] = 29'b0_011000010010_001_0_010010011000;
      patterns[12434] = 29'b0_011000010010_010_0_110000100100;
      patterns[12435] = 29'b0_011000010010_011_1_100001001000;
      patterns[12436] = 29'b0_011000010010_100_0_001100001001;
      patterns[12437] = 29'b0_011000010010_101_1_000110000100;
      patterns[12438] = 29'b0_011000010010_110_0_011000010010;
      patterns[12439] = 29'b0_011000010010_111_0_011000010010;
      patterns[12440] = 29'b0_011000010011_000_0_011000010011;
      patterns[12441] = 29'b0_011000010011_001_0_010011011000;
      patterns[12442] = 29'b0_011000010011_010_0_110000100110;
      patterns[12443] = 29'b0_011000010011_011_1_100001001100;
      patterns[12444] = 29'b0_011000010011_100_1_001100001001;
      patterns[12445] = 29'b0_011000010011_101_1_100110000100;
      patterns[12446] = 29'b0_011000010011_110_0_011000010011;
      patterns[12447] = 29'b0_011000010011_111_0_011000010011;
      patterns[12448] = 29'b0_011000010100_000_0_011000010100;
      patterns[12449] = 29'b0_011000010100_001_0_010100011000;
      patterns[12450] = 29'b0_011000010100_010_0_110000101000;
      patterns[12451] = 29'b0_011000010100_011_1_100001010000;
      patterns[12452] = 29'b0_011000010100_100_0_001100001010;
      patterns[12453] = 29'b0_011000010100_101_0_000110000101;
      patterns[12454] = 29'b0_011000010100_110_0_011000010100;
      patterns[12455] = 29'b0_011000010100_111_0_011000010100;
      patterns[12456] = 29'b0_011000010101_000_0_011000010101;
      patterns[12457] = 29'b0_011000010101_001_0_010101011000;
      patterns[12458] = 29'b0_011000010101_010_0_110000101010;
      patterns[12459] = 29'b0_011000010101_011_1_100001010100;
      patterns[12460] = 29'b0_011000010101_100_1_001100001010;
      patterns[12461] = 29'b0_011000010101_101_0_100110000101;
      patterns[12462] = 29'b0_011000010101_110_0_011000010101;
      patterns[12463] = 29'b0_011000010101_111_0_011000010101;
      patterns[12464] = 29'b0_011000010110_000_0_011000010110;
      patterns[12465] = 29'b0_011000010110_001_0_010110011000;
      patterns[12466] = 29'b0_011000010110_010_0_110000101100;
      patterns[12467] = 29'b0_011000010110_011_1_100001011000;
      patterns[12468] = 29'b0_011000010110_100_0_001100001011;
      patterns[12469] = 29'b0_011000010110_101_1_000110000101;
      patterns[12470] = 29'b0_011000010110_110_0_011000010110;
      patterns[12471] = 29'b0_011000010110_111_0_011000010110;
      patterns[12472] = 29'b0_011000010111_000_0_011000010111;
      patterns[12473] = 29'b0_011000010111_001_0_010111011000;
      patterns[12474] = 29'b0_011000010111_010_0_110000101110;
      patterns[12475] = 29'b0_011000010111_011_1_100001011100;
      patterns[12476] = 29'b0_011000010111_100_1_001100001011;
      patterns[12477] = 29'b0_011000010111_101_1_100110000101;
      patterns[12478] = 29'b0_011000010111_110_0_011000010111;
      patterns[12479] = 29'b0_011000010111_111_0_011000010111;
      patterns[12480] = 29'b0_011000011000_000_0_011000011000;
      patterns[12481] = 29'b0_011000011000_001_0_011000011000;
      patterns[12482] = 29'b0_011000011000_010_0_110000110000;
      patterns[12483] = 29'b0_011000011000_011_1_100001100000;
      patterns[12484] = 29'b0_011000011000_100_0_001100001100;
      patterns[12485] = 29'b0_011000011000_101_0_000110000110;
      patterns[12486] = 29'b0_011000011000_110_0_011000011000;
      patterns[12487] = 29'b0_011000011000_111_0_011000011000;
      patterns[12488] = 29'b0_011000011001_000_0_011000011001;
      patterns[12489] = 29'b0_011000011001_001_0_011001011000;
      patterns[12490] = 29'b0_011000011001_010_0_110000110010;
      patterns[12491] = 29'b0_011000011001_011_1_100001100100;
      patterns[12492] = 29'b0_011000011001_100_1_001100001100;
      patterns[12493] = 29'b0_011000011001_101_0_100110000110;
      patterns[12494] = 29'b0_011000011001_110_0_011000011001;
      patterns[12495] = 29'b0_011000011001_111_0_011000011001;
      patterns[12496] = 29'b0_011000011010_000_0_011000011010;
      patterns[12497] = 29'b0_011000011010_001_0_011010011000;
      patterns[12498] = 29'b0_011000011010_010_0_110000110100;
      patterns[12499] = 29'b0_011000011010_011_1_100001101000;
      patterns[12500] = 29'b0_011000011010_100_0_001100001101;
      patterns[12501] = 29'b0_011000011010_101_1_000110000110;
      patterns[12502] = 29'b0_011000011010_110_0_011000011010;
      patterns[12503] = 29'b0_011000011010_111_0_011000011010;
      patterns[12504] = 29'b0_011000011011_000_0_011000011011;
      patterns[12505] = 29'b0_011000011011_001_0_011011011000;
      patterns[12506] = 29'b0_011000011011_010_0_110000110110;
      patterns[12507] = 29'b0_011000011011_011_1_100001101100;
      patterns[12508] = 29'b0_011000011011_100_1_001100001101;
      patterns[12509] = 29'b0_011000011011_101_1_100110000110;
      patterns[12510] = 29'b0_011000011011_110_0_011000011011;
      patterns[12511] = 29'b0_011000011011_111_0_011000011011;
      patterns[12512] = 29'b0_011000011100_000_0_011000011100;
      patterns[12513] = 29'b0_011000011100_001_0_011100011000;
      patterns[12514] = 29'b0_011000011100_010_0_110000111000;
      patterns[12515] = 29'b0_011000011100_011_1_100001110000;
      patterns[12516] = 29'b0_011000011100_100_0_001100001110;
      patterns[12517] = 29'b0_011000011100_101_0_000110000111;
      patterns[12518] = 29'b0_011000011100_110_0_011000011100;
      patterns[12519] = 29'b0_011000011100_111_0_011000011100;
      patterns[12520] = 29'b0_011000011101_000_0_011000011101;
      patterns[12521] = 29'b0_011000011101_001_0_011101011000;
      patterns[12522] = 29'b0_011000011101_010_0_110000111010;
      patterns[12523] = 29'b0_011000011101_011_1_100001110100;
      patterns[12524] = 29'b0_011000011101_100_1_001100001110;
      patterns[12525] = 29'b0_011000011101_101_0_100110000111;
      patterns[12526] = 29'b0_011000011101_110_0_011000011101;
      patterns[12527] = 29'b0_011000011101_111_0_011000011101;
      patterns[12528] = 29'b0_011000011110_000_0_011000011110;
      patterns[12529] = 29'b0_011000011110_001_0_011110011000;
      patterns[12530] = 29'b0_011000011110_010_0_110000111100;
      patterns[12531] = 29'b0_011000011110_011_1_100001111000;
      patterns[12532] = 29'b0_011000011110_100_0_001100001111;
      patterns[12533] = 29'b0_011000011110_101_1_000110000111;
      patterns[12534] = 29'b0_011000011110_110_0_011000011110;
      patterns[12535] = 29'b0_011000011110_111_0_011000011110;
      patterns[12536] = 29'b0_011000011111_000_0_011000011111;
      patterns[12537] = 29'b0_011000011111_001_0_011111011000;
      patterns[12538] = 29'b0_011000011111_010_0_110000111110;
      patterns[12539] = 29'b0_011000011111_011_1_100001111100;
      patterns[12540] = 29'b0_011000011111_100_1_001100001111;
      patterns[12541] = 29'b0_011000011111_101_1_100110000111;
      patterns[12542] = 29'b0_011000011111_110_0_011000011111;
      patterns[12543] = 29'b0_011000011111_111_0_011000011111;
      patterns[12544] = 29'b0_011000100000_000_0_011000100000;
      patterns[12545] = 29'b0_011000100000_001_0_100000011000;
      patterns[12546] = 29'b0_011000100000_010_0_110001000000;
      patterns[12547] = 29'b0_011000100000_011_1_100010000000;
      patterns[12548] = 29'b0_011000100000_100_0_001100010000;
      patterns[12549] = 29'b0_011000100000_101_0_000110001000;
      patterns[12550] = 29'b0_011000100000_110_0_011000100000;
      patterns[12551] = 29'b0_011000100000_111_0_011000100000;
      patterns[12552] = 29'b0_011000100001_000_0_011000100001;
      patterns[12553] = 29'b0_011000100001_001_0_100001011000;
      patterns[12554] = 29'b0_011000100001_010_0_110001000010;
      patterns[12555] = 29'b0_011000100001_011_1_100010000100;
      patterns[12556] = 29'b0_011000100001_100_1_001100010000;
      patterns[12557] = 29'b0_011000100001_101_0_100110001000;
      patterns[12558] = 29'b0_011000100001_110_0_011000100001;
      patterns[12559] = 29'b0_011000100001_111_0_011000100001;
      patterns[12560] = 29'b0_011000100010_000_0_011000100010;
      patterns[12561] = 29'b0_011000100010_001_0_100010011000;
      patterns[12562] = 29'b0_011000100010_010_0_110001000100;
      patterns[12563] = 29'b0_011000100010_011_1_100010001000;
      patterns[12564] = 29'b0_011000100010_100_0_001100010001;
      patterns[12565] = 29'b0_011000100010_101_1_000110001000;
      patterns[12566] = 29'b0_011000100010_110_0_011000100010;
      patterns[12567] = 29'b0_011000100010_111_0_011000100010;
      patterns[12568] = 29'b0_011000100011_000_0_011000100011;
      patterns[12569] = 29'b0_011000100011_001_0_100011011000;
      patterns[12570] = 29'b0_011000100011_010_0_110001000110;
      patterns[12571] = 29'b0_011000100011_011_1_100010001100;
      patterns[12572] = 29'b0_011000100011_100_1_001100010001;
      patterns[12573] = 29'b0_011000100011_101_1_100110001000;
      patterns[12574] = 29'b0_011000100011_110_0_011000100011;
      patterns[12575] = 29'b0_011000100011_111_0_011000100011;
      patterns[12576] = 29'b0_011000100100_000_0_011000100100;
      patterns[12577] = 29'b0_011000100100_001_0_100100011000;
      patterns[12578] = 29'b0_011000100100_010_0_110001001000;
      patterns[12579] = 29'b0_011000100100_011_1_100010010000;
      patterns[12580] = 29'b0_011000100100_100_0_001100010010;
      patterns[12581] = 29'b0_011000100100_101_0_000110001001;
      patterns[12582] = 29'b0_011000100100_110_0_011000100100;
      patterns[12583] = 29'b0_011000100100_111_0_011000100100;
      patterns[12584] = 29'b0_011000100101_000_0_011000100101;
      patterns[12585] = 29'b0_011000100101_001_0_100101011000;
      patterns[12586] = 29'b0_011000100101_010_0_110001001010;
      patterns[12587] = 29'b0_011000100101_011_1_100010010100;
      patterns[12588] = 29'b0_011000100101_100_1_001100010010;
      patterns[12589] = 29'b0_011000100101_101_0_100110001001;
      patterns[12590] = 29'b0_011000100101_110_0_011000100101;
      patterns[12591] = 29'b0_011000100101_111_0_011000100101;
      patterns[12592] = 29'b0_011000100110_000_0_011000100110;
      patterns[12593] = 29'b0_011000100110_001_0_100110011000;
      patterns[12594] = 29'b0_011000100110_010_0_110001001100;
      patterns[12595] = 29'b0_011000100110_011_1_100010011000;
      patterns[12596] = 29'b0_011000100110_100_0_001100010011;
      patterns[12597] = 29'b0_011000100110_101_1_000110001001;
      patterns[12598] = 29'b0_011000100110_110_0_011000100110;
      patterns[12599] = 29'b0_011000100110_111_0_011000100110;
      patterns[12600] = 29'b0_011000100111_000_0_011000100111;
      patterns[12601] = 29'b0_011000100111_001_0_100111011000;
      patterns[12602] = 29'b0_011000100111_010_0_110001001110;
      patterns[12603] = 29'b0_011000100111_011_1_100010011100;
      patterns[12604] = 29'b0_011000100111_100_1_001100010011;
      patterns[12605] = 29'b0_011000100111_101_1_100110001001;
      patterns[12606] = 29'b0_011000100111_110_0_011000100111;
      patterns[12607] = 29'b0_011000100111_111_0_011000100111;
      patterns[12608] = 29'b0_011000101000_000_0_011000101000;
      patterns[12609] = 29'b0_011000101000_001_0_101000011000;
      patterns[12610] = 29'b0_011000101000_010_0_110001010000;
      patterns[12611] = 29'b0_011000101000_011_1_100010100000;
      patterns[12612] = 29'b0_011000101000_100_0_001100010100;
      patterns[12613] = 29'b0_011000101000_101_0_000110001010;
      patterns[12614] = 29'b0_011000101000_110_0_011000101000;
      patterns[12615] = 29'b0_011000101000_111_0_011000101000;
      patterns[12616] = 29'b0_011000101001_000_0_011000101001;
      patterns[12617] = 29'b0_011000101001_001_0_101001011000;
      patterns[12618] = 29'b0_011000101001_010_0_110001010010;
      patterns[12619] = 29'b0_011000101001_011_1_100010100100;
      patterns[12620] = 29'b0_011000101001_100_1_001100010100;
      patterns[12621] = 29'b0_011000101001_101_0_100110001010;
      patterns[12622] = 29'b0_011000101001_110_0_011000101001;
      patterns[12623] = 29'b0_011000101001_111_0_011000101001;
      patterns[12624] = 29'b0_011000101010_000_0_011000101010;
      patterns[12625] = 29'b0_011000101010_001_0_101010011000;
      patterns[12626] = 29'b0_011000101010_010_0_110001010100;
      patterns[12627] = 29'b0_011000101010_011_1_100010101000;
      patterns[12628] = 29'b0_011000101010_100_0_001100010101;
      patterns[12629] = 29'b0_011000101010_101_1_000110001010;
      patterns[12630] = 29'b0_011000101010_110_0_011000101010;
      patterns[12631] = 29'b0_011000101010_111_0_011000101010;
      patterns[12632] = 29'b0_011000101011_000_0_011000101011;
      patterns[12633] = 29'b0_011000101011_001_0_101011011000;
      patterns[12634] = 29'b0_011000101011_010_0_110001010110;
      patterns[12635] = 29'b0_011000101011_011_1_100010101100;
      patterns[12636] = 29'b0_011000101011_100_1_001100010101;
      patterns[12637] = 29'b0_011000101011_101_1_100110001010;
      patterns[12638] = 29'b0_011000101011_110_0_011000101011;
      patterns[12639] = 29'b0_011000101011_111_0_011000101011;
      patterns[12640] = 29'b0_011000101100_000_0_011000101100;
      patterns[12641] = 29'b0_011000101100_001_0_101100011000;
      patterns[12642] = 29'b0_011000101100_010_0_110001011000;
      patterns[12643] = 29'b0_011000101100_011_1_100010110000;
      patterns[12644] = 29'b0_011000101100_100_0_001100010110;
      patterns[12645] = 29'b0_011000101100_101_0_000110001011;
      patterns[12646] = 29'b0_011000101100_110_0_011000101100;
      patterns[12647] = 29'b0_011000101100_111_0_011000101100;
      patterns[12648] = 29'b0_011000101101_000_0_011000101101;
      patterns[12649] = 29'b0_011000101101_001_0_101101011000;
      patterns[12650] = 29'b0_011000101101_010_0_110001011010;
      patterns[12651] = 29'b0_011000101101_011_1_100010110100;
      patterns[12652] = 29'b0_011000101101_100_1_001100010110;
      patterns[12653] = 29'b0_011000101101_101_0_100110001011;
      patterns[12654] = 29'b0_011000101101_110_0_011000101101;
      patterns[12655] = 29'b0_011000101101_111_0_011000101101;
      patterns[12656] = 29'b0_011000101110_000_0_011000101110;
      patterns[12657] = 29'b0_011000101110_001_0_101110011000;
      patterns[12658] = 29'b0_011000101110_010_0_110001011100;
      patterns[12659] = 29'b0_011000101110_011_1_100010111000;
      patterns[12660] = 29'b0_011000101110_100_0_001100010111;
      patterns[12661] = 29'b0_011000101110_101_1_000110001011;
      patterns[12662] = 29'b0_011000101110_110_0_011000101110;
      patterns[12663] = 29'b0_011000101110_111_0_011000101110;
      patterns[12664] = 29'b0_011000101111_000_0_011000101111;
      patterns[12665] = 29'b0_011000101111_001_0_101111011000;
      patterns[12666] = 29'b0_011000101111_010_0_110001011110;
      patterns[12667] = 29'b0_011000101111_011_1_100010111100;
      patterns[12668] = 29'b0_011000101111_100_1_001100010111;
      patterns[12669] = 29'b0_011000101111_101_1_100110001011;
      patterns[12670] = 29'b0_011000101111_110_0_011000101111;
      patterns[12671] = 29'b0_011000101111_111_0_011000101111;
      patterns[12672] = 29'b0_011000110000_000_0_011000110000;
      patterns[12673] = 29'b0_011000110000_001_0_110000011000;
      patterns[12674] = 29'b0_011000110000_010_0_110001100000;
      patterns[12675] = 29'b0_011000110000_011_1_100011000000;
      patterns[12676] = 29'b0_011000110000_100_0_001100011000;
      patterns[12677] = 29'b0_011000110000_101_0_000110001100;
      patterns[12678] = 29'b0_011000110000_110_0_011000110000;
      patterns[12679] = 29'b0_011000110000_111_0_011000110000;
      patterns[12680] = 29'b0_011000110001_000_0_011000110001;
      patterns[12681] = 29'b0_011000110001_001_0_110001011000;
      patterns[12682] = 29'b0_011000110001_010_0_110001100010;
      patterns[12683] = 29'b0_011000110001_011_1_100011000100;
      patterns[12684] = 29'b0_011000110001_100_1_001100011000;
      patterns[12685] = 29'b0_011000110001_101_0_100110001100;
      patterns[12686] = 29'b0_011000110001_110_0_011000110001;
      patterns[12687] = 29'b0_011000110001_111_0_011000110001;
      patterns[12688] = 29'b0_011000110010_000_0_011000110010;
      patterns[12689] = 29'b0_011000110010_001_0_110010011000;
      patterns[12690] = 29'b0_011000110010_010_0_110001100100;
      patterns[12691] = 29'b0_011000110010_011_1_100011001000;
      patterns[12692] = 29'b0_011000110010_100_0_001100011001;
      patterns[12693] = 29'b0_011000110010_101_1_000110001100;
      patterns[12694] = 29'b0_011000110010_110_0_011000110010;
      patterns[12695] = 29'b0_011000110010_111_0_011000110010;
      patterns[12696] = 29'b0_011000110011_000_0_011000110011;
      patterns[12697] = 29'b0_011000110011_001_0_110011011000;
      patterns[12698] = 29'b0_011000110011_010_0_110001100110;
      patterns[12699] = 29'b0_011000110011_011_1_100011001100;
      patterns[12700] = 29'b0_011000110011_100_1_001100011001;
      patterns[12701] = 29'b0_011000110011_101_1_100110001100;
      patterns[12702] = 29'b0_011000110011_110_0_011000110011;
      patterns[12703] = 29'b0_011000110011_111_0_011000110011;
      patterns[12704] = 29'b0_011000110100_000_0_011000110100;
      patterns[12705] = 29'b0_011000110100_001_0_110100011000;
      patterns[12706] = 29'b0_011000110100_010_0_110001101000;
      patterns[12707] = 29'b0_011000110100_011_1_100011010000;
      patterns[12708] = 29'b0_011000110100_100_0_001100011010;
      patterns[12709] = 29'b0_011000110100_101_0_000110001101;
      patterns[12710] = 29'b0_011000110100_110_0_011000110100;
      patterns[12711] = 29'b0_011000110100_111_0_011000110100;
      patterns[12712] = 29'b0_011000110101_000_0_011000110101;
      patterns[12713] = 29'b0_011000110101_001_0_110101011000;
      patterns[12714] = 29'b0_011000110101_010_0_110001101010;
      patterns[12715] = 29'b0_011000110101_011_1_100011010100;
      patterns[12716] = 29'b0_011000110101_100_1_001100011010;
      patterns[12717] = 29'b0_011000110101_101_0_100110001101;
      patterns[12718] = 29'b0_011000110101_110_0_011000110101;
      patterns[12719] = 29'b0_011000110101_111_0_011000110101;
      patterns[12720] = 29'b0_011000110110_000_0_011000110110;
      patterns[12721] = 29'b0_011000110110_001_0_110110011000;
      patterns[12722] = 29'b0_011000110110_010_0_110001101100;
      patterns[12723] = 29'b0_011000110110_011_1_100011011000;
      patterns[12724] = 29'b0_011000110110_100_0_001100011011;
      patterns[12725] = 29'b0_011000110110_101_1_000110001101;
      patterns[12726] = 29'b0_011000110110_110_0_011000110110;
      patterns[12727] = 29'b0_011000110110_111_0_011000110110;
      patterns[12728] = 29'b0_011000110111_000_0_011000110111;
      patterns[12729] = 29'b0_011000110111_001_0_110111011000;
      patterns[12730] = 29'b0_011000110111_010_0_110001101110;
      patterns[12731] = 29'b0_011000110111_011_1_100011011100;
      patterns[12732] = 29'b0_011000110111_100_1_001100011011;
      patterns[12733] = 29'b0_011000110111_101_1_100110001101;
      patterns[12734] = 29'b0_011000110111_110_0_011000110111;
      patterns[12735] = 29'b0_011000110111_111_0_011000110111;
      patterns[12736] = 29'b0_011000111000_000_0_011000111000;
      patterns[12737] = 29'b0_011000111000_001_0_111000011000;
      patterns[12738] = 29'b0_011000111000_010_0_110001110000;
      patterns[12739] = 29'b0_011000111000_011_1_100011100000;
      patterns[12740] = 29'b0_011000111000_100_0_001100011100;
      patterns[12741] = 29'b0_011000111000_101_0_000110001110;
      patterns[12742] = 29'b0_011000111000_110_0_011000111000;
      patterns[12743] = 29'b0_011000111000_111_0_011000111000;
      patterns[12744] = 29'b0_011000111001_000_0_011000111001;
      patterns[12745] = 29'b0_011000111001_001_0_111001011000;
      patterns[12746] = 29'b0_011000111001_010_0_110001110010;
      patterns[12747] = 29'b0_011000111001_011_1_100011100100;
      patterns[12748] = 29'b0_011000111001_100_1_001100011100;
      patterns[12749] = 29'b0_011000111001_101_0_100110001110;
      patterns[12750] = 29'b0_011000111001_110_0_011000111001;
      patterns[12751] = 29'b0_011000111001_111_0_011000111001;
      patterns[12752] = 29'b0_011000111010_000_0_011000111010;
      patterns[12753] = 29'b0_011000111010_001_0_111010011000;
      patterns[12754] = 29'b0_011000111010_010_0_110001110100;
      patterns[12755] = 29'b0_011000111010_011_1_100011101000;
      patterns[12756] = 29'b0_011000111010_100_0_001100011101;
      patterns[12757] = 29'b0_011000111010_101_1_000110001110;
      patterns[12758] = 29'b0_011000111010_110_0_011000111010;
      patterns[12759] = 29'b0_011000111010_111_0_011000111010;
      patterns[12760] = 29'b0_011000111011_000_0_011000111011;
      patterns[12761] = 29'b0_011000111011_001_0_111011011000;
      patterns[12762] = 29'b0_011000111011_010_0_110001110110;
      patterns[12763] = 29'b0_011000111011_011_1_100011101100;
      patterns[12764] = 29'b0_011000111011_100_1_001100011101;
      patterns[12765] = 29'b0_011000111011_101_1_100110001110;
      patterns[12766] = 29'b0_011000111011_110_0_011000111011;
      patterns[12767] = 29'b0_011000111011_111_0_011000111011;
      patterns[12768] = 29'b0_011000111100_000_0_011000111100;
      patterns[12769] = 29'b0_011000111100_001_0_111100011000;
      patterns[12770] = 29'b0_011000111100_010_0_110001111000;
      patterns[12771] = 29'b0_011000111100_011_1_100011110000;
      patterns[12772] = 29'b0_011000111100_100_0_001100011110;
      patterns[12773] = 29'b0_011000111100_101_0_000110001111;
      patterns[12774] = 29'b0_011000111100_110_0_011000111100;
      patterns[12775] = 29'b0_011000111100_111_0_011000111100;
      patterns[12776] = 29'b0_011000111101_000_0_011000111101;
      patterns[12777] = 29'b0_011000111101_001_0_111101011000;
      patterns[12778] = 29'b0_011000111101_010_0_110001111010;
      patterns[12779] = 29'b0_011000111101_011_1_100011110100;
      patterns[12780] = 29'b0_011000111101_100_1_001100011110;
      patterns[12781] = 29'b0_011000111101_101_0_100110001111;
      patterns[12782] = 29'b0_011000111101_110_0_011000111101;
      patterns[12783] = 29'b0_011000111101_111_0_011000111101;
      patterns[12784] = 29'b0_011000111110_000_0_011000111110;
      patterns[12785] = 29'b0_011000111110_001_0_111110011000;
      patterns[12786] = 29'b0_011000111110_010_0_110001111100;
      patterns[12787] = 29'b0_011000111110_011_1_100011111000;
      patterns[12788] = 29'b0_011000111110_100_0_001100011111;
      patterns[12789] = 29'b0_011000111110_101_1_000110001111;
      patterns[12790] = 29'b0_011000111110_110_0_011000111110;
      patterns[12791] = 29'b0_011000111110_111_0_011000111110;
      patterns[12792] = 29'b0_011000111111_000_0_011000111111;
      patterns[12793] = 29'b0_011000111111_001_0_111111011000;
      patterns[12794] = 29'b0_011000111111_010_0_110001111110;
      patterns[12795] = 29'b0_011000111111_011_1_100011111100;
      patterns[12796] = 29'b0_011000111111_100_1_001100011111;
      patterns[12797] = 29'b0_011000111111_101_1_100110001111;
      patterns[12798] = 29'b0_011000111111_110_0_011000111111;
      patterns[12799] = 29'b0_011000111111_111_0_011000111111;
      patterns[12800] = 29'b0_011001000000_000_0_011001000000;
      patterns[12801] = 29'b0_011001000000_001_0_000000011001;
      patterns[12802] = 29'b0_011001000000_010_0_110010000000;
      patterns[12803] = 29'b0_011001000000_011_1_100100000000;
      patterns[12804] = 29'b0_011001000000_100_0_001100100000;
      patterns[12805] = 29'b0_011001000000_101_0_000110010000;
      patterns[12806] = 29'b0_011001000000_110_0_011001000000;
      patterns[12807] = 29'b0_011001000000_111_0_011001000000;
      patterns[12808] = 29'b0_011001000001_000_0_011001000001;
      patterns[12809] = 29'b0_011001000001_001_0_000001011001;
      patterns[12810] = 29'b0_011001000001_010_0_110010000010;
      patterns[12811] = 29'b0_011001000001_011_1_100100000100;
      patterns[12812] = 29'b0_011001000001_100_1_001100100000;
      patterns[12813] = 29'b0_011001000001_101_0_100110010000;
      patterns[12814] = 29'b0_011001000001_110_0_011001000001;
      patterns[12815] = 29'b0_011001000001_111_0_011001000001;
      patterns[12816] = 29'b0_011001000010_000_0_011001000010;
      patterns[12817] = 29'b0_011001000010_001_0_000010011001;
      patterns[12818] = 29'b0_011001000010_010_0_110010000100;
      patterns[12819] = 29'b0_011001000010_011_1_100100001000;
      patterns[12820] = 29'b0_011001000010_100_0_001100100001;
      patterns[12821] = 29'b0_011001000010_101_1_000110010000;
      patterns[12822] = 29'b0_011001000010_110_0_011001000010;
      patterns[12823] = 29'b0_011001000010_111_0_011001000010;
      patterns[12824] = 29'b0_011001000011_000_0_011001000011;
      patterns[12825] = 29'b0_011001000011_001_0_000011011001;
      patterns[12826] = 29'b0_011001000011_010_0_110010000110;
      patterns[12827] = 29'b0_011001000011_011_1_100100001100;
      patterns[12828] = 29'b0_011001000011_100_1_001100100001;
      patterns[12829] = 29'b0_011001000011_101_1_100110010000;
      patterns[12830] = 29'b0_011001000011_110_0_011001000011;
      patterns[12831] = 29'b0_011001000011_111_0_011001000011;
      patterns[12832] = 29'b0_011001000100_000_0_011001000100;
      patterns[12833] = 29'b0_011001000100_001_0_000100011001;
      patterns[12834] = 29'b0_011001000100_010_0_110010001000;
      patterns[12835] = 29'b0_011001000100_011_1_100100010000;
      patterns[12836] = 29'b0_011001000100_100_0_001100100010;
      patterns[12837] = 29'b0_011001000100_101_0_000110010001;
      patterns[12838] = 29'b0_011001000100_110_0_011001000100;
      patterns[12839] = 29'b0_011001000100_111_0_011001000100;
      patterns[12840] = 29'b0_011001000101_000_0_011001000101;
      patterns[12841] = 29'b0_011001000101_001_0_000101011001;
      patterns[12842] = 29'b0_011001000101_010_0_110010001010;
      patterns[12843] = 29'b0_011001000101_011_1_100100010100;
      patterns[12844] = 29'b0_011001000101_100_1_001100100010;
      patterns[12845] = 29'b0_011001000101_101_0_100110010001;
      patterns[12846] = 29'b0_011001000101_110_0_011001000101;
      patterns[12847] = 29'b0_011001000101_111_0_011001000101;
      patterns[12848] = 29'b0_011001000110_000_0_011001000110;
      patterns[12849] = 29'b0_011001000110_001_0_000110011001;
      patterns[12850] = 29'b0_011001000110_010_0_110010001100;
      patterns[12851] = 29'b0_011001000110_011_1_100100011000;
      patterns[12852] = 29'b0_011001000110_100_0_001100100011;
      patterns[12853] = 29'b0_011001000110_101_1_000110010001;
      patterns[12854] = 29'b0_011001000110_110_0_011001000110;
      patterns[12855] = 29'b0_011001000110_111_0_011001000110;
      patterns[12856] = 29'b0_011001000111_000_0_011001000111;
      patterns[12857] = 29'b0_011001000111_001_0_000111011001;
      patterns[12858] = 29'b0_011001000111_010_0_110010001110;
      patterns[12859] = 29'b0_011001000111_011_1_100100011100;
      patterns[12860] = 29'b0_011001000111_100_1_001100100011;
      patterns[12861] = 29'b0_011001000111_101_1_100110010001;
      patterns[12862] = 29'b0_011001000111_110_0_011001000111;
      patterns[12863] = 29'b0_011001000111_111_0_011001000111;
      patterns[12864] = 29'b0_011001001000_000_0_011001001000;
      patterns[12865] = 29'b0_011001001000_001_0_001000011001;
      patterns[12866] = 29'b0_011001001000_010_0_110010010000;
      patterns[12867] = 29'b0_011001001000_011_1_100100100000;
      patterns[12868] = 29'b0_011001001000_100_0_001100100100;
      patterns[12869] = 29'b0_011001001000_101_0_000110010010;
      patterns[12870] = 29'b0_011001001000_110_0_011001001000;
      patterns[12871] = 29'b0_011001001000_111_0_011001001000;
      patterns[12872] = 29'b0_011001001001_000_0_011001001001;
      patterns[12873] = 29'b0_011001001001_001_0_001001011001;
      patterns[12874] = 29'b0_011001001001_010_0_110010010010;
      patterns[12875] = 29'b0_011001001001_011_1_100100100100;
      patterns[12876] = 29'b0_011001001001_100_1_001100100100;
      patterns[12877] = 29'b0_011001001001_101_0_100110010010;
      patterns[12878] = 29'b0_011001001001_110_0_011001001001;
      patterns[12879] = 29'b0_011001001001_111_0_011001001001;
      patterns[12880] = 29'b0_011001001010_000_0_011001001010;
      patterns[12881] = 29'b0_011001001010_001_0_001010011001;
      patterns[12882] = 29'b0_011001001010_010_0_110010010100;
      patterns[12883] = 29'b0_011001001010_011_1_100100101000;
      patterns[12884] = 29'b0_011001001010_100_0_001100100101;
      patterns[12885] = 29'b0_011001001010_101_1_000110010010;
      patterns[12886] = 29'b0_011001001010_110_0_011001001010;
      patterns[12887] = 29'b0_011001001010_111_0_011001001010;
      patterns[12888] = 29'b0_011001001011_000_0_011001001011;
      patterns[12889] = 29'b0_011001001011_001_0_001011011001;
      patterns[12890] = 29'b0_011001001011_010_0_110010010110;
      patterns[12891] = 29'b0_011001001011_011_1_100100101100;
      patterns[12892] = 29'b0_011001001011_100_1_001100100101;
      patterns[12893] = 29'b0_011001001011_101_1_100110010010;
      patterns[12894] = 29'b0_011001001011_110_0_011001001011;
      patterns[12895] = 29'b0_011001001011_111_0_011001001011;
      patterns[12896] = 29'b0_011001001100_000_0_011001001100;
      patterns[12897] = 29'b0_011001001100_001_0_001100011001;
      patterns[12898] = 29'b0_011001001100_010_0_110010011000;
      patterns[12899] = 29'b0_011001001100_011_1_100100110000;
      patterns[12900] = 29'b0_011001001100_100_0_001100100110;
      patterns[12901] = 29'b0_011001001100_101_0_000110010011;
      patterns[12902] = 29'b0_011001001100_110_0_011001001100;
      patterns[12903] = 29'b0_011001001100_111_0_011001001100;
      patterns[12904] = 29'b0_011001001101_000_0_011001001101;
      patterns[12905] = 29'b0_011001001101_001_0_001101011001;
      patterns[12906] = 29'b0_011001001101_010_0_110010011010;
      patterns[12907] = 29'b0_011001001101_011_1_100100110100;
      patterns[12908] = 29'b0_011001001101_100_1_001100100110;
      patterns[12909] = 29'b0_011001001101_101_0_100110010011;
      patterns[12910] = 29'b0_011001001101_110_0_011001001101;
      patterns[12911] = 29'b0_011001001101_111_0_011001001101;
      patterns[12912] = 29'b0_011001001110_000_0_011001001110;
      patterns[12913] = 29'b0_011001001110_001_0_001110011001;
      patterns[12914] = 29'b0_011001001110_010_0_110010011100;
      patterns[12915] = 29'b0_011001001110_011_1_100100111000;
      patterns[12916] = 29'b0_011001001110_100_0_001100100111;
      patterns[12917] = 29'b0_011001001110_101_1_000110010011;
      patterns[12918] = 29'b0_011001001110_110_0_011001001110;
      patterns[12919] = 29'b0_011001001110_111_0_011001001110;
      patterns[12920] = 29'b0_011001001111_000_0_011001001111;
      patterns[12921] = 29'b0_011001001111_001_0_001111011001;
      patterns[12922] = 29'b0_011001001111_010_0_110010011110;
      patterns[12923] = 29'b0_011001001111_011_1_100100111100;
      patterns[12924] = 29'b0_011001001111_100_1_001100100111;
      patterns[12925] = 29'b0_011001001111_101_1_100110010011;
      patterns[12926] = 29'b0_011001001111_110_0_011001001111;
      patterns[12927] = 29'b0_011001001111_111_0_011001001111;
      patterns[12928] = 29'b0_011001010000_000_0_011001010000;
      patterns[12929] = 29'b0_011001010000_001_0_010000011001;
      patterns[12930] = 29'b0_011001010000_010_0_110010100000;
      patterns[12931] = 29'b0_011001010000_011_1_100101000000;
      patterns[12932] = 29'b0_011001010000_100_0_001100101000;
      patterns[12933] = 29'b0_011001010000_101_0_000110010100;
      patterns[12934] = 29'b0_011001010000_110_0_011001010000;
      patterns[12935] = 29'b0_011001010000_111_0_011001010000;
      patterns[12936] = 29'b0_011001010001_000_0_011001010001;
      patterns[12937] = 29'b0_011001010001_001_0_010001011001;
      patterns[12938] = 29'b0_011001010001_010_0_110010100010;
      patterns[12939] = 29'b0_011001010001_011_1_100101000100;
      patterns[12940] = 29'b0_011001010001_100_1_001100101000;
      patterns[12941] = 29'b0_011001010001_101_0_100110010100;
      patterns[12942] = 29'b0_011001010001_110_0_011001010001;
      patterns[12943] = 29'b0_011001010001_111_0_011001010001;
      patterns[12944] = 29'b0_011001010010_000_0_011001010010;
      patterns[12945] = 29'b0_011001010010_001_0_010010011001;
      patterns[12946] = 29'b0_011001010010_010_0_110010100100;
      patterns[12947] = 29'b0_011001010010_011_1_100101001000;
      patterns[12948] = 29'b0_011001010010_100_0_001100101001;
      patterns[12949] = 29'b0_011001010010_101_1_000110010100;
      patterns[12950] = 29'b0_011001010010_110_0_011001010010;
      patterns[12951] = 29'b0_011001010010_111_0_011001010010;
      patterns[12952] = 29'b0_011001010011_000_0_011001010011;
      patterns[12953] = 29'b0_011001010011_001_0_010011011001;
      patterns[12954] = 29'b0_011001010011_010_0_110010100110;
      patterns[12955] = 29'b0_011001010011_011_1_100101001100;
      patterns[12956] = 29'b0_011001010011_100_1_001100101001;
      patterns[12957] = 29'b0_011001010011_101_1_100110010100;
      patterns[12958] = 29'b0_011001010011_110_0_011001010011;
      patterns[12959] = 29'b0_011001010011_111_0_011001010011;
      patterns[12960] = 29'b0_011001010100_000_0_011001010100;
      patterns[12961] = 29'b0_011001010100_001_0_010100011001;
      patterns[12962] = 29'b0_011001010100_010_0_110010101000;
      patterns[12963] = 29'b0_011001010100_011_1_100101010000;
      patterns[12964] = 29'b0_011001010100_100_0_001100101010;
      patterns[12965] = 29'b0_011001010100_101_0_000110010101;
      patterns[12966] = 29'b0_011001010100_110_0_011001010100;
      patterns[12967] = 29'b0_011001010100_111_0_011001010100;
      patterns[12968] = 29'b0_011001010101_000_0_011001010101;
      patterns[12969] = 29'b0_011001010101_001_0_010101011001;
      patterns[12970] = 29'b0_011001010101_010_0_110010101010;
      patterns[12971] = 29'b0_011001010101_011_1_100101010100;
      patterns[12972] = 29'b0_011001010101_100_1_001100101010;
      patterns[12973] = 29'b0_011001010101_101_0_100110010101;
      patterns[12974] = 29'b0_011001010101_110_0_011001010101;
      patterns[12975] = 29'b0_011001010101_111_0_011001010101;
      patterns[12976] = 29'b0_011001010110_000_0_011001010110;
      patterns[12977] = 29'b0_011001010110_001_0_010110011001;
      patterns[12978] = 29'b0_011001010110_010_0_110010101100;
      patterns[12979] = 29'b0_011001010110_011_1_100101011000;
      patterns[12980] = 29'b0_011001010110_100_0_001100101011;
      patterns[12981] = 29'b0_011001010110_101_1_000110010101;
      patterns[12982] = 29'b0_011001010110_110_0_011001010110;
      patterns[12983] = 29'b0_011001010110_111_0_011001010110;
      patterns[12984] = 29'b0_011001010111_000_0_011001010111;
      patterns[12985] = 29'b0_011001010111_001_0_010111011001;
      patterns[12986] = 29'b0_011001010111_010_0_110010101110;
      patterns[12987] = 29'b0_011001010111_011_1_100101011100;
      patterns[12988] = 29'b0_011001010111_100_1_001100101011;
      patterns[12989] = 29'b0_011001010111_101_1_100110010101;
      patterns[12990] = 29'b0_011001010111_110_0_011001010111;
      patterns[12991] = 29'b0_011001010111_111_0_011001010111;
      patterns[12992] = 29'b0_011001011000_000_0_011001011000;
      patterns[12993] = 29'b0_011001011000_001_0_011000011001;
      patterns[12994] = 29'b0_011001011000_010_0_110010110000;
      patterns[12995] = 29'b0_011001011000_011_1_100101100000;
      patterns[12996] = 29'b0_011001011000_100_0_001100101100;
      patterns[12997] = 29'b0_011001011000_101_0_000110010110;
      patterns[12998] = 29'b0_011001011000_110_0_011001011000;
      patterns[12999] = 29'b0_011001011000_111_0_011001011000;
      patterns[13000] = 29'b0_011001011001_000_0_011001011001;
      patterns[13001] = 29'b0_011001011001_001_0_011001011001;
      patterns[13002] = 29'b0_011001011001_010_0_110010110010;
      patterns[13003] = 29'b0_011001011001_011_1_100101100100;
      patterns[13004] = 29'b0_011001011001_100_1_001100101100;
      patterns[13005] = 29'b0_011001011001_101_0_100110010110;
      patterns[13006] = 29'b0_011001011001_110_0_011001011001;
      patterns[13007] = 29'b0_011001011001_111_0_011001011001;
      patterns[13008] = 29'b0_011001011010_000_0_011001011010;
      patterns[13009] = 29'b0_011001011010_001_0_011010011001;
      patterns[13010] = 29'b0_011001011010_010_0_110010110100;
      patterns[13011] = 29'b0_011001011010_011_1_100101101000;
      patterns[13012] = 29'b0_011001011010_100_0_001100101101;
      patterns[13013] = 29'b0_011001011010_101_1_000110010110;
      patterns[13014] = 29'b0_011001011010_110_0_011001011010;
      patterns[13015] = 29'b0_011001011010_111_0_011001011010;
      patterns[13016] = 29'b0_011001011011_000_0_011001011011;
      patterns[13017] = 29'b0_011001011011_001_0_011011011001;
      patterns[13018] = 29'b0_011001011011_010_0_110010110110;
      patterns[13019] = 29'b0_011001011011_011_1_100101101100;
      patterns[13020] = 29'b0_011001011011_100_1_001100101101;
      patterns[13021] = 29'b0_011001011011_101_1_100110010110;
      patterns[13022] = 29'b0_011001011011_110_0_011001011011;
      patterns[13023] = 29'b0_011001011011_111_0_011001011011;
      patterns[13024] = 29'b0_011001011100_000_0_011001011100;
      patterns[13025] = 29'b0_011001011100_001_0_011100011001;
      patterns[13026] = 29'b0_011001011100_010_0_110010111000;
      patterns[13027] = 29'b0_011001011100_011_1_100101110000;
      patterns[13028] = 29'b0_011001011100_100_0_001100101110;
      patterns[13029] = 29'b0_011001011100_101_0_000110010111;
      patterns[13030] = 29'b0_011001011100_110_0_011001011100;
      patterns[13031] = 29'b0_011001011100_111_0_011001011100;
      patterns[13032] = 29'b0_011001011101_000_0_011001011101;
      patterns[13033] = 29'b0_011001011101_001_0_011101011001;
      patterns[13034] = 29'b0_011001011101_010_0_110010111010;
      patterns[13035] = 29'b0_011001011101_011_1_100101110100;
      patterns[13036] = 29'b0_011001011101_100_1_001100101110;
      patterns[13037] = 29'b0_011001011101_101_0_100110010111;
      patterns[13038] = 29'b0_011001011101_110_0_011001011101;
      patterns[13039] = 29'b0_011001011101_111_0_011001011101;
      patterns[13040] = 29'b0_011001011110_000_0_011001011110;
      patterns[13041] = 29'b0_011001011110_001_0_011110011001;
      patterns[13042] = 29'b0_011001011110_010_0_110010111100;
      patterns[13043] = 29'b0_011001011110_011_1_100101111000;
      patterns[13044] = 29'b0_011001011110_100_0_001100101111;
      patterns[13045] = 29'b0_011001011110_101_1_000110010111;
      patterns[13046] = 29'b0_011001011110_110_0_011001011110;
      patterns[13047] = 29'b0_011001011110_111_0_011001011110;
      patterns[13048] = 29'b0_011001011111_000_0_011001011111;
      patterns[13049] = 29'b0_011001011111_001_0_011111011001;
      patterns[13050] = 29'b0_011001011111_010_0_110010111110;
      patterns[13051] = 29'b0_011001011111_011_1_100101111100;
      patterns[13052] = 29'b0_011001011111_100_1_001100101111;
      patterns[13053] = 29'b0_011001011111_101_1_100110010111;
      patterns[13054] = 29'b0_011001011111_110_0_011001011111;
      patterns[13055] = 29'b0_011001011111_111_0_011001011111;
      patterns[13056] = 29'b0_011001100000_000_0_011001100000;
      patterns[13057] = 29'b0_011001100000_001_0_100000011001;
      patterns[13058] = 29'b0_011001100000_010_0_110011000000;
      patterns[13059] = 29'b0_011001100000_011_1_100110000000;
      patterns[13060] = 29'b0_011001100000_100_0_001100110000;
      patterns[13061] = 29'b0_011001100000_101_0_000110011000;
      patterns[13062] = 29'b0_011001100000_110_0_011001100000;
      patterns[13063] = 29'b0_011001100000_111_0_011001100000;
      patterns[13064] = 29'b0_011001100001_000_0_011001100001;
      patterns[13065] = 29'b0_011001100001_001_0_100001011001;
      patterns[13066] = 29'b0_011001100001_010_0_110011000010;
      patterns[13067] = 29'b0_011001100001_011_1_100110000100;
      patterns[13068] = 29'b0_011001100001_100_1_001100110000;
      patterns[13069] = 29'b0_011001100001_101_0_100110011000;
      patterns[13070] = 29'b0_011001100001_110_0_011001100001;
      patterns[13071] = 29'b0_011001100001_111_0_011001100001;
      patterns[13072] = 29'b0_011001100010_000_0_011001100010;
      patterns[13073] = 29'b0_011001100010_001_0_100010011001;
      patterns[13074] = 29'b0_011001100010_010_0_110011000100;
      patterns[13075] = 29'b0_011001100010_011_1_100110001000;
      patterns[13076] = 29'b0_011001100010_100_0_001100110001;
      patterns[13077] = 29'b0_011001100010_101_1_000110011000;
      patterns[13078] = 29'b0_011001100010_110_0_011001100010;
      patterns[13079] = 29'b0_011001100010_111_0_011001100010;
      patterns[13080] = 29'b0_011001100011_000_0_011001100011;
      patterns[13081] = 29'b0_011001100011_001_0_100011011001;
      patterns[13082] = 29'b0_011001100011_010_0_110011000110;
      patterns[13083] = 29'b0_011001100011_011_1_100110001100;
      patterns[13084] = 29'b0_011001100011_100_1_001100110001;
      patterns[13085] = 29'b0_011001100011_101_1_100110011000;
      patterns[13086] = 29'b0_011001100011_110_0_011001100011;
      patterns[13087] = 29'b0_011001100011_111_0_011001100011;
      patterns[13088] = 29'b0_011001100100_000_0_011001100100;
      patterns[13089] = 29'b0_011001100100_001_0_100100011001;
      patterns[13090] = 29'b0_011001100100_010_0_110011001000;
      patterns[13091] = 29'b0_011001100100_011_1_100110010000;
      patterns[13092] = 29'b0_011001100100_100_0_001100110010;
      patterns[13093] = 29'b0_011001100100_101_0_000110011001;
      patterns[13094] = 29'b0_011001100100_110_0_011001100100;
      patterns[13095] = 29'b0_011001100100_111_0_011001100100;
      patterns[13096] = 29'b0_011001100101_000_0_011001100101;
      patterns[13097] = 29'b0_011001100101_001_0_100101011001;
      patterns[13098] = 29'b0_011001100101_010_0_110011001010;
      patterns[13099] = 29'b0_011001100101_011_1_100110010100;
      patterns[13100] = 29'b0_011001100101_100_1_001100110010;
      patterns[13101] = 29'b0_011001100101_101_0_100110011001;
      patterns[13102] = 29'b0_011001100101_110_0_011001100101;
      patterns[13103] = 29'b0_011001100101_111_0_011001100101;
      patterns[13104] = 29'b0_011001100110_000_0_011001100110;
      patterns[13105] = 29'b0_011001100110_001_0_100110011001;
      patterns[13106] = 29'b0_011001100110_010_0_110011001100;
      patterns[13107] = 29'b0_011001100110_011_1_100110011000;
      patterns[13108] = 29'b0_011001100110_100_0_001100110011;
      patterns[13109] = 29'b0_011001100110_101_1_000110011001;
      patterns[13110] = 29'b0_011001100110_110_0_011001100110;
      patterns[13111] = 29'b0_011001100110_111_0_011001100110;
      patterns[13112] = 29'b0_011001100111_000_0_011001100111;
      patterns[13113] = 29'b0_011001100111_001_0_100111011001;
      patterns[13114] = 29'b0_011001100111_010_0_110011001110;
      patterns[13115] = 29'b0_011001100111_011_1_100110011100;
      patterns[13116] = 29'b0_011001100111_100_1_001100110011;
      patterns[13117] = 29'b0_011001100111_101_1_100110011001;
      patterns[13118] = 29'b0_011001100111_110_0_011001100111;
      patterns[13119] = 29'b0_011001100111_111_0_011001100111;
      patterns[13120] = 29'b0_011001101000_000_0_011001101000;
      patterns[13121] = 29'b0_011001101000_001_0_101000011001;
      patterns[13122] = 29'b0_011001101000_010_0_110011010000;
      patterns[13123] = 29'b0_011001101000_011_1_100110100000;
      patterns[13124] = 29'b0_011001101000_100_0_001100110100;
      patterns[13125] = 29'b0_011001101000_101_0_000110011010;
      patterns[13126] = 29'b0_011001101000_110_0_011001101000;
      patterns[13127] = 29'b0_011001101000_111_0_011001101000;
      patterns[13128] = 29'b0_011001101001_000_0_011001101001;
      patterns[13129] = 29'b0_011001101001_001_0_101001011001;
      patterns[13130] = 29'b0_011001101001_010_0_110011010010;
      patterns[13131] = 29'b0_011001101001_011_1_100110100100;
      patterns[13132] = 29'b0_011001101001_100_1_001100110100;
      patterns[13133] = 29'b0_011001101001_101_0_100110011010;
      patterns[13134] = 29'b0_011001101001_110_0_011001101001;
      patterns[13135] = 29'b0_011001101001_111_0_011001101001;
      patterns[13136] = 29'b0_011001101010_000_0_011001101010;
      patterns[13137] = 29'b0_011001101010_001_0_101010011001;
      patterns[13138] = 29'b0_011001101010_010_0_110011010100;
      patterns[13139] = 29'b0_011001101010_011_1_100110101000;
      patterns[13140] = 29'b0_011001101010_100_0_001100110101;
      patterns[13141] = 29'b0_011001101010_101_1_000110011010;
      patterns[13142] = 29'b0_011001101010_110_0_011001101010;
      patterns[13143] = 29'b0_011001101010_111_0_011001101010;
      patterns[13144] = 29'b0_011001101011_000_0_011001101011;
      patterns[13145] = 29'b0_011001101011_001_0_101011011001;
      patterns[13146] = 29'b0_011001101011_010_0_110011010110;
      patterns[13147] = 29'b0_011001101011_011_1_100110101100;
      patterns[13148] = 29'b0_011001101011_100_1_001100110101;
      patterns[13149] = 29'b0_011001101011_101_1_100110011010;
      patterns[13150] = 29'b0_011001101011_110_0_011001101011;
      patterns[13151] = 29'b0_011001101011_111_0_011001101011;
      patterns[13152] = 29'b0_011001101100_000_0_011001101100;
      patterns[13153] = 29'b0_011001101100_001_0_101100011001;
      patterns[13154] = 29'b0_011001101100_010_0_110011011000;
      patterns[13155] = 29'b0_011001101100_011_1_100110110000;
      patterns[13156] = 29'b0_011001101100_100_0_001100110110;
      patterns[13157] = 29'b0_011001101100_101_0_000110011011;
      patterns[13158] = 29'b0_011001101100_110_0_011001101100;
      patterns[13159] = 29'b0_011001101100_111_0_011001101100;
      patterns[13160] = 29'b0_011001101101_000_0_011001101101;
      patterns[13161] = 29'b0_011001101101_001_0_101101011001;
      patterns[13162] = 29'b0_011001101101_010_0_110011011010;
      patterns[13163] = 29'b0_011001101101_011_1_100110110100;
      patterns[13164] = 29'b0_011001101101_100_1_001100110110;
      patterns[13165] = 29'b0_011001101101_101_0_100110011011;
      patterns[13166] = 29'b0_011001101101_110_0_011001101101;
      patterns[13167] = 29'b0_011001101101_111_0_011001101101;
      patterns[13168] = 29'b0_011001101110_000_0_011001101110;
      patterns[13169] = 29'b0_011001101110_001_0_101110011001;
      patterns[13170] = 29'b0_011001101110_010_0_110011011100;
      patterns[13171] = 29'b0_011001101110_011_1_100110111000;
      patterns[13172] = 29'b0_011001101110_100_0_001100110111;
      patterns[13173] = 29'b0_011001101110_101_1_000110011011;
      patterns[13174] = 29'b0_011001101110_110_0_011001101110;
      patterns[13175] = 29'b0_011001101110_111_0_011001101110;
      patterns[13176] = 29'b0_011001101111_000_0_011001101111;
      patterns[13177] = 29'b0_011001101111_001_0_101111011001;
      patterns[13178] = 29'b0_011001101111_010_0_110011011110;
      patterns[13179] = 29'b0_011001101111_011_1_100110111100;
      patterns[13180] = 29'b0_011001101111_100_1_001100110111;
      patterns[13181] = 29'b0_011001101111_101_1_100110011011;
      patterns[13182] = 29'b0_011001101111_110_0_011001101111;
      patterns[13183] = 29'b0_011001101111_111_0_011001101111;
      patterns[13184] = 29'b0_011001110000_000_0_011001110000;
      patterns[13185] = 29'b0_011001110000_001_0_110000011001;
      patterns[13186] = 29'b0_011001110000_010_0_110011100000;
      patterns[13187] = 29'b0_011001110000_011_1_100111000000;
      patterns[13188] = 29'b0_011001110000_100_0_001100111000;
      patterns[13189] = 29'b0_011001110000_101_0_000110011100;
      patterns[13190] = 29'b0_011001110000_110_0_011001110000;
      patterns[13191] = 29'b0_011001110000_111_0_011001110000;
      patterns[13192] = 29'b0_011001110001_000_0_011001110001;
      patterns[13193] = 29'b0_011001110001_001_0_110001011001;
      patterns[13194] = 29'b0_011001110001_010_0_110011100010;
      patterns[13195] = 29'b0_011001110001_011_1_100111000100;
      patterns[13196] = 29'b0_011001110001_100_1_001100111000;
      patterns[13197] = 29'b0_011001110001_101_0_100110011100;
      patterns[13198] = 29'b0_011001110001_110_0_011001110001;
      patterns[13199] = 29'b0_011001110001_111_0_011001110001;
      patterns[13200] = 29'b0_011001110010_000_0_011001110010;
      patterns[13201] = 29'b0_011001110010_001_0_110010011001;
      patterns[13202] = 29'b0_011001110010_010_0_110011100100;
      patterns[13203] = 29'b0_011001110010_011_1_100111001000;
      patterns[13204] = 29'b0_011001110010_100_0_001100111001;
      patterns[13205] = 29'b0_011001110010_101_1_000110011100;
      patterns[13206] = 29'b0_011001110010_110_0_011001110010;
      patterns[13207] = 29'b0_011001110010_111_0_011001110010;
      patterns[13208] = 29'b0_011001110011_000_0_011001110011;
      patterns[13209] = 29'b0_011001110011_001_0_110011011001;
      patterns[13210] = 29'b0_011001110011_010_0_110011100110;
      patterns[13211] = 29'b0_011001110011_011_1_100111001100;
      patterns[13212] = 29'b0_011001110011_100_1_001100111001;
      patterns[13213] = 29'b0_011001110011_101_1_100110011100;
      patterns[13214] = 29'b0_011001110011_110_0_011001110011;
      patterns[13215] = 29'b0_011001110011_111_0_011001110011;
      patterns[13216] = 29'b0_011001110100_000_0_011001110100;
      patterns[13217] = 29'b0_011001110100_001_0_110100011001;
      patterns[13218] = 29'b0_011001110100_010_0_110011101000;
      patterns[13219] = 29'b0_011001110100_011_1_100111010000;
      patterns[13220] = 29'b0_011001110100_100_0_001100111010;
      patterns[13221] = 29'b0_011001110100_101_0_000110011101;
      patterns[13222] = 29'b0_011001110100_110_0_011001110100;
      patterns[13223] = 29'b0_011001110100_111_0_011001110100;
      patterns[13224] = 29'b0_011001110101_000_0_011001110101;
      patterns[13225] = 29'b0_011001110101_001_0_110101011001;
      patterns[13226] = 29'b0_011001110101_010_0_110011101010;
      patterns[13227] = 29'b0_011001110101_011_1_100111010100;
      patterns[13228] = 29'b0_011001110101_100_1_001100111010;
      patterns[13229] = 29'b0_011001110101_101_0_100110011101;
      patterns[13230] = 29'b0_011001110101_110_0_011001110101;
      patterns[13231] = 29'b0_011001110101_111_0_011001110101;
      patterns[13232] = 29'b0_011001110110_000_0_011001110110;
      patterns[13233] = 29'b0_011001110110_001_0_110110011001;
      patterns[13234] = 29'b0_011001110110_010_0_110011101100;
      patterns[13235] = 29'b0_011001110110_011_1_100111011000;
      patterns[13236] = 29'b0_011001110110_100_0_001100111011;
      patterns[13237] = 29'b0_011001110110_101_1_000110011101;
      patterns[13238] = 29'b0_011001110110_110_0_011001110110;
      patterns[13239] = 29'b0_011001110110_111_0_011001110110;
      patterns[13240] = 29'b0_011001110111_000_0_011001110111;
      patterns[13241] = 29'b0_011001110111_001_0_110111011001;
      patterns[13242] = 29'b0_011001110111_010_0_110011101110;
      patterns[13243] = 29'b0_011001110111_011_1_100111011100;
      patterns[13244] = 29'b0_011001110111_100_1_001100111011;
      patterns[13245] = 29'b0_011001110111_101_1_100110011101;
      patterns[13246] = 29'b0_011001110111_110_0_011001110111;
      patterns[13247] = 29'b0_011001110111_111_0_011001110111;
      patterns[13248] = 29'b0_011001111000_000_0_011001111000;
      patterns[13249] = 29'b0_011001111000_001_0_111000011001;
      patterns[13250] = 29'b0_011001111000_010_0_110011110000;
      patterns[13251] = 29'b0_011001111000_011_1_100111100000;
      patterns[13252] = 29'b0_011001111000_100_0_001100111100;
      patterns[13253] = 29'b0_011001111000_101_0_000110011110;
      patterns[13254] = 29'b0_011001111000_110_0_011001111000;
      patterns[13255] = 29'b0_011001111000_111_0_011001111000;
      patterns[13256] = 29'b0_011001111001_000_0_011001111001;
      patterns[13257] = 29'b0_011001111001_001_0_111001011001;
      patterns[13258] = 29'b0_011001111001_010_0_110011110010;
      patterns[13259] = 29'b0_011001111001_011_1_100111100100;
      patterns[13260] = 29'b0_011001111001_100_1_001100111100;
      patterns[13261] = 29'b0_011001111001_101_0_100110011110;
      patterns[13262] = 29'b0_011001111001_110_0_011001111001;
      patterns[13263] = 29'b0_011001111001_111_0_011001111001;
      patterns[13264] = 29'b0_011001111010_000_0_011001111010;
      patterns[13265] = 29'b0_011001111010_001_0_111010011001;
      patterns[13266] = 29'b0_011001111010_010_0_110011110100;
      patterns[13267] = 29'b0_011001111010_011_1_100111101000;
      patterns[13268] = 29'b0_011001111010_100_0_001100111101;
      patterns[13269] = 29'b0_011001111010_101_1_000110011110;
      patterns[13270] = 29'b0_011001111010_110_0_011001111010;
      patterns[13271] = 29'b0_011001111010_111_0_011001111010;
      patterns[13272] = 29'b0_011001111011_000_0_011001111011;
      patterns[13273] = 29'b0_011001111011_001_0_111011011001;
      patterns[13274] = 29'b0_011001111011_010_0_110011110110;
      patterns[13275] = 29'b0_011001111011_011_1_100111101100;
      patterns[13276] = 29'b0_011001111011_100_1_001100111101;
      patterns[13277] = 29'b0_011001111011_101_1_100110011110;
      patterns[13278] = 29'b0_011001111011_110_0_011001111011;
      patterns[13279] = 29'b0_011001111011_111_0_011001111011;
      patterns[13280] = 29'b0_011001111100_000_0_011001111100;
      patterns[13281] = 29'b0_011001111100_001_0_111100011001;
      patterns[13282] = 29'b0_011001111100_010_0_110011111000;
      patterns[13283] = 29'b0_011001111100_011_1_100111110000;
      patterns[13284] = 29'b0_011001111100_100_0_001100111110;
      patterns[13285] = 29'b0_011001111100_101_0_000110011111;
      patterns[13286] = 29'b0_011001111100_110_0_011001111100;
      patterns[13287] = 29'b0_011001111100_111_0_011001111100;
      patterns[13288] = 29'b0_011001111101_000_0_011001111101;
      patterns[13289] = 29'b0_011001111101_001_0_111101011001;
      patterns[13290] = 29'b0_011001111101_010_0_110011111010;
      patterns[13291] = 29'b0_011001111101_011_1_100111110100;
      patterns[13292] = 29'b0_011001111101_100_1_001100111110;
      patterns[13293] = 29'b0_011001111101_101_0_100110011111;
      patterns[13294] = 29'b0_011001111101_110_0_011001111101;
      patterns[13295] = 29'b0_011001111101_111_0_011001111101;
      patterns[13296] = 29'b0_011001111110_000_0_011001111110;
      patterns[13297] = 29'b0_011001111110_001_0_111110011001;
      patterns[13298] = 29'b0_011001111110_010_0_110011111100;
      patterns[13299] = 29'b0_011001111110_011_1_100111111000;
      patterns[13300] = 29'b0_011001111110_100_0_001100111111;
      patterns[13301] = 29'b0_011001111110_101_1_000110011111;
      patterns[13302] = 29'b0_011001111110_110_0_011001111110;
      patterns[13303] = 29'b0_011001111110_111_0_011001111110;
      patterns[13304] = 29'b0_011001111111_000_0_011001111111;
      patterns[13305] = 29'b0_011001111111_001_0_111111011001;
      patterns[13306] = 29'b0_011001111111_010_0_110011111110;
      patterns[13307] = 29'b0_011001111111_011_1_100111111100;
      patterns[13308] = 29'b0_011001111111_100_1_001100111111;
      patterns[13309] = 29'b0_011001111111_101_1_100110011111;
      patterns[13310] = 29'b0_011001111111_110_0_011001111111;
      patterns[13311] = 29'b0_011001111111_111_0_011001111111;
      patterns[13312] = 29'b0_011010000000_000_0_011010000000;
      patterns[13313] = 29'b0_011010000000_001_0_000000011010;
      patterns[13314] = 29'b0_011010000000_010_0_110100000000;
      patterns[13315] = 29'b0_011010000000_011_1_101000000000;
      patterns[13316] = 29'b0_011010000000_100_0_001101000000;
      patterns[13317] = 29'b0_011010000000_101_0_000110100000;
      patterns[13318] = 29'b0_011010000000_110_0_011010000000;
      patterns[13319] = 29'b0_011010000000_111_0_011010000000;
      patterns[13320] = 29'b0_011010000001_000_0_011010000001;
      patterns[13321] = 29'b0_011010000001_001_0_000001011010;
      patterns[13322] = 29'b0_011010000001_010_0_110100000010;
      patterns[13323] = 29'b0_011010000001_011_1_101000000100;
      patterns[13324] = 29'b0_011010000001_100_1_001101000000;
      patterns[13325] = 29'b0_011010000001_101_0_100110100000;
      patterns[13326] = 29'b0_011010000001_110_0_011010000001;
      patterns[13327] = 29'b0_011010000001_111_0_011010000001;
      patterns[13328] = 29'b0_011010000010_000_0_011010000010;
      patterns[13329] = 29'b0_011010000010_001_0_000010011010;
      patterns[13330] = 29'b0_011010000010_010_0_110100000100;
      patterns[13331] = 29'b0_011010000010_011_1_101000001000;
      patterns[13332] = 29'b0_011010000010_100_0_001101000001;
      patterns[13333] = 29'b0_011010000010_101_1_000110100000;
      patterns[13334] = 29'b0_011010000010_110_0_011010000010;
      patterns[13335] = 29'b0_011010000010_111_0_011010000010;
      patterns[13336] = 29'b0_011010000011_000_0_011010000011;
      patterns[13337] = 29'b0_011010000011_001_0_000011011010;
      patterns[13338] = 29'b0_011010000011_010_0_110100000110;
      patterns[13339] = 29'b0_011010000011_011_1_101000001100;
      patterns[13340] = 29'b0_011010000011_100_1_001101000001;
      patterns[13341] = 29'b0_011010000011_101_1_100110100000;
      patterns[13342] = 29'b0_011010000011_110_0_011010000011;
      patterns[13343] = 29'b0_011010000011_111_0_011010000011;
      patterns[13344] = 29'b0_011010000100_000_0_011010000100;
      patterns[13345] = 29'b0_011010000100_001_0_000100011010;
      patterns[13346] = 29'b0_011010000100_010_0_110100001000;
      patterns[13347] = 29'b0_011010000100_011_1_101000010000;
      patterns[13348] = 29'b0_011010000100_100_0_001101000010;
      patterns[13349] = 29'b0_011010000100_101_0_000110100001;
      patterns[13350] = 29'b0_011010000100_110_0_011010000100;
      patterns[13351] = 29'b0_011010000100_111_0_011010000100;
      patterns[13352] = 29'b0_011010000101_000_0_011010000101;
      patterns[13353] = 29'b0_011010000101_001_0_000101011010;
      patterns[13354] = 29'b0_011010000101_010_0_110100001010;
      patterns[13355] = 29'b0_011010000101_011_1_101000010100;
      patterns[13356] = 29'b0_011010000101_100_1_001101000010;
      patterns[13357] = 29'b0_011010000101_101_0_100110100001;
      patterns[13358] = 29'b0_011010000101_110_0_011010000101;
      patterns[13359] = 29'b0_011010000101_111_0_011010000101;
      patterns[13360] = 29'b0_011010000110_000_0_011010000110;
      patterns[13361] = 29'b0_011010000110_001_0_000110011010;
      patterns[13362] = 29'b0_011010000110_010_0_110100001100;
      patterns[13363] = 29'b0_011010000110_011_1_101000011000;
      patterns[13364] = 29'b0_011010000110_100_0_001101000011;
      patterns[13365] = 29'b0_011010000110_101_1_000110100001;
      patterns[13366] = 29'b0_011010000110_110_0_011010000110;
      patterns[13367] = 29'b0_011010000110_111_0_011010000110;
      patterns[13368] = 29'b0_011010000111_000_0_011010000111;
      patterns[13369] = 29'b0_011010000111_001_0_000111011010;
      patterns[13370] = 29'b0_011010000111_010_0_110100001110;
      patterns[13371] = 29'b0_011010000111_011_1_101000011100;
      patterns[13372] = 29'b0_011010000111_100_1_001101000011;
      patterns[13373] = 29'b0_011010000111_101_1_100110100001;
      patterns[13374] = 29'b0_011010000111_110_0_011010000111;
      patterns[13375] = 29'b0_011010000111_111_0_011010000111;
      patterns[13376] = 29'b0_011010001000_000_0_011010001000;
      patterns[13377] = 29'b0_011010001000_001_0_001000011010;
      patterns[13378] = 29'b0_011010001000_010_0_110100010000;
      patterns[13379] = 29'b0_011010001000_011_1_101000100000;
      patterns[13380] = 29'b0_011010001000_100_0_001101000100;
      patterns[13381] = 29'b0_011010001000_101_0_000110100010;
      patterns[13382] = 29'b0_011010001000_110_0_011010001000;
      patterns[13383] = 29'b0_011010001000_111_0_011010001000;
      patterns[13384] = 29'b0_011010001001_000_0_011010001001;
      patterns[13385] = 29'b0_011010001001_001_0_001001011010;
      patterns[13386] = 29'b0_011010001001_010_0_110100010010;
      patterns[13387] = 29'b0_011010001001_011_1_101000100100;
      patterns[13388] = 29'b0_011010001001_100_1_001101000100;
      patterns[13389] = 29'b0_011010001001_101_0_100110100010;
      patterns[13390] = 29'b0_011010001001_110_0_011010001001;
      patterns[13391] = 29'b0_011010001001_111_0_011010001001;
      patterns[13392] = 29'b0_011010001010_000_0_011010001010;
      patterns[13393] = 29'b0_011010001010_001_0_001010011010;
      patterns[13394] = 29'b0_011010001010_010_0_110100010100;
      patterns[13395] = 29'b0_011010001010_011_1_101000101000;
      patterns[13396] = 29'b0_011010001010_100_0_001101000101;
      patterns[13397] = 29'b0_011010001010_101_1_000110100010;
      patterns[13398] = 29'b0_011010001010_110_0_011010001010;
      patterns[13399] = 29'b0_011010001010_111_0_011010001010;
      patterns[13400] = 29'b0_011010001011_000_0_011010001011;
      patterns[13401] = 29'b0_011010001011_001_0_001011011010;
      patterns[13402] = 29'b0_011010001011_010_0_110100010110;
      patterns[13403] = 29'b0_011010001011_011_1_101000101100;
      patterns[13404] = 29'b0_011010001011_100_1_001101000101;
      patterns[13405] = 29'b0_011010001011_101_1_100110100010;
      patterns[13406] = 29'b0_011010001011_110_0_011010001011;
      patterns[13407] = 29'b0_011010001011_111_0_011010001011;
      patterns[13408] = 29'b0_011010001100_000_0_011010001100;
      patterns[13409] = 29'b0_011010001100_001_0_001100011010;
      patterns[13410] = 29'b0_011010001100_010_0_110100011000;
      patterns[13411] = 29'b0_011010001100_011_1_101000110000;
      patterns[13412] = 29'b0_011010001100_100_0_001101000110;
      patterns[13413] = 29'b0_011010001100_101_0_000110100011;
      patterns[13414] = 29'b0_011010001100_110_0_011010001100;
      patterns[13415] = 29'b0_011010001100_111_0_011010001100;
      patterns[13416] = 29'b0_011010001101_000_0_011010001101;
      patterns[13417] = 29'b0_011010001101_001_0_001101011010;
      patterns[13418] = 29'b0_011010001101_010_0_110100011010;
      patterns[13419] = 29'b0_011010001101_011_1_101000110100;
      patterns[13420] = 29'b0_011010001101_100_1_001101000110;
      patterns[13421] = 29'b0_011010001101_101_0_100110100011;
      patterns[13422] = 29'b0_011010001101_110_0_011010001101;
      patterns[13423] = 29'b0_011010001101_111_0_011010001101;
      patterns[13424] = 29'b0_011010001110_000_0_011010001110;
      patterns[13425] = 29'b0_011010001110_001_0_001110011010;
      patterns[13426] = 29'b0_011010001110_010_0_110100011100;
      patterns[13427] = 29'b0_011010001110_011_1_101000111000;
      patterns[13428] = 29'b0_011010001110_100_0_001101000111;
      patterns[13429] = 29'b0_011010001110_101_1_000110100011;
      patterns[13430] = 29'b0_011010001110_110_0_011010001110;
      patterns[13431] = 29'b0_011010001110_111_0_011010001110;
      patterns[13432] = 29'b0_011010001111_000_0_011010001111;
      patterns[13433] = 29'b0_011010001111_001_0_001111011010;
      patterns[13434] = 29'b0_011010001111_010_0_110100011110;
      patterns[13435] = 29'b0_011010001111_011_1_101000111100;
      patterns[13436] = 29'b0_011010001111_100_1_001101000111;
      patterns[13437] = 29'b0_011010001111_101_1_100110100011;
      patterns[13438] = 29'b0_011010001111_110_0_011010001111;
      patterns[13439] = 29'b0_011010001111_111_0_011010001111;
      patterns[13440] = 29'b0_011010010000_000_0_011010010000;
      patterns[13441] = 29'b0_011010010000_001_0_010000011010;
      patterns[13442] = 29'b0_011010010000_010_0_110100100000;
      patterns[13443] = 29'b0_011010010000_011_1_101001000000;
      patterns[13444] = 29'b0_011010010000_100_0_001101001000;
      patterns[13445] = 29'b0_011010010000_101_0_000110100100;
      patterns[13446] = 29'b0_011010010000_110_0_011010010000;
      patterns[13447] = 29'b0_011010010000_111_0_011010010000;
      patterns[13448] = 29'b0_011010010001_000_0_011010010001;
      patterns[13449] = 29'b0_011010010001_001_0_010001011010;
      patterns[13450] = 29'b0_011010010001_010_0_110100100010;
      patterns[13451] = 29'b0_011010010001_011_1_101001000100;
      patterns[13452] = 29'b0_011010010001_100_1_001101001000;
      patterns[13453] = 29'b0_011010010001_101_0_100110100100;
      patterns[13454] = 29'b0_011010010001_110_0_011010010001;
      patterns[13455] = 29'b0_011010010001_111_0_011010010001;
      patterns[13456] = 29'b0_011010010010_000_0_011010010010;
      patterns[13457] = 29'b0_011010010010_001_0_010010011010;
      patterns[13458] = 29'b0_011010010010_010_0_110100100100;
      patterns[13459] = 29'b0_011010010010_011_1_101001001000;
      patterns[13460] = 29'b0_011010010010_100_0_001101001001;
      patterns[13461] = 29'b0_011010010010_101_1_000110100100;
      patterns[13462] = 29'b0_011010010010_110_0_011010010010;
      patterns[13463] = 29'b0_011010010010_111_0_011010010010;
      patterns[13464] = 29'b0_011010010011_000_0_011010010011;
      patterns[13465] = 29'b0_011010010011_001_0_010011011010;
      patterns[13466] = 29'b0_011010010011_010_0_110100100110;
      patterns[13467] = 29'b0_011010010011_011_1_101001001100;
      patterns[13468] = 29'b0_011010010011_100_1_001101001001;
      patterns[13469] = 29'b0_011010010011_101_1_100110100100;
      patterns[13470] = 29'b0_011010010011_110_0_011010010011;
      patterns[13471] = 29'b0_011010010011_111_0_011010010011;
      patterns[13472] = 29'b0_011010010100_000_0_011010010100;
      patterns[13473] = 29'b0_011010010100_001_0_010100011010;
      patterns[13474] = 29'b0_011010010100_010_0_110100101000;
      patterns[13475] = 29'b0_011010010100_011_1_101001010000;
      patterns[13476] = 29'b0_011010010100_100_0_001101001010;
      patterns[13477] = 29'b0_011010010100_101_0_000110100101;
      patterns[13478] = 29'b0_011010010100_110_0_011010010100;
      patterns[13479] = 29'b0_011010010100_111_0_011010010100;
      patterns[13480] = 29'b0_011010010101_000_0_011010010101;
      patterns[13481] = 29'b0_011010010101_001_0_010101011010;
      patterns[13482] = 29'b0_011010010101_010_0_110100101010;
      patterns[13483] = 29'b0_011010010101_011_1_101001010100;
      patterns[13484] = 29'b0_011010010101_100_1_001101001010;
      patterns[13485] = 29'b0_011010010101_101_0_100110100101;
      patterns[13486] = 29'b0_011010010101_110_0_011010010101;
      patterns[13487] = 29'b0_011010010101_111_0_011010010101;
      patterns[13488] = 29'b0_011010010110_000_0_011010010110;
      patterns[13489] = 29'b0_011010010110_001_0_010110011010;
      patterns[13490] = 29'b0_011010010110_010_0_110100101100;
      patterns[13491] = 29'b0_011010010110_011_1_101001011000;
      patterns[13492] = 29'b0_011010010110_100_0_001101001011;
      patterns[13493] = 29'b0_011010010110_101_1_000110100101;
      patterns[13494] = 29'b0_011010010110_110_0_011010010110;
      patterns[13495] = 29'b0_011010010110_111_0_011010010110;
      patterns[13496] = 29'b0_011010010111_000_0_011010010111;
      patterns[13497] = 29'b0_011010010111_001_0_010111011010;
      patterns[13498] = 29'b0_011010010111_010_0_110100101110;
      patterns[13499] = 29'b0_011010010111_011_1_101001011100;
      patterns[13500] = 29'b0_011010010111_100_1_001101001011;
      patterns[13501] = 29'b0_011010010111_101_1_100110100101;
      patterns[13502] = 29'b0_011010010111_110_0_011010010111;
      patterns[13503] = 29'b0_011010010111_111_0_011010010111;
      patterns[13504] = 29'b0_011010011000_000_0_011010011000;
      patterns[13505] = 29'b0_011010011000_001_0_011000011010;
      patterns[13506] = 29'b0_011010011000_010_0_110100110000;
      patterns[13507] = 29'b0_011010011000_011_1_101001100000;
      patterns[13508] = 29'b0_011010011000_100_0_001101001100;
      patterns[13509] = 29'b0_011010011000_101_0_000110100110;
      patterns[13510] = 29'b0_011010011000_110_0_011010011000;
      patterns[13511] = 29'b0_011010011000_111_0_011010011000;
      patterns[13512] = 29'b0_011010011001_000_0_011010011001;
      patterns[13513] = 29'b0_011010011001_001_0_011001011010;
      patterns[13514] = 29'b0_011010011001_010_0_110100110010;
      patterns[13515] = 29'b0_011010011001_011_1_101001100100;
      patterns[13516] = 29'b0_011010011001_100_1_001101001100;
      patterns[13517] = 29'b0_011010011001_101_0_100110100110;
      patterns[13518] = 29'b0_011010011001_110_0_011010011001;
      patterns[13519] = 29'b0_011010011001_111_0_011010011001;
      patterns[13520] = 29'b0_011010011010_000_0_011010011010;
      patterns[13521] = 29'b0_011010011010_001_0_011010011010;
      patterns[13522] = 29'b0_011010011010_010_0_110100110100;
      patterns[13523] = 29'b0_011010011010_011_1_101001101000;
      patterns[13524] = 29'b0_011010011010_100_0_001101001101;
      patterns[13525] = 29'b0_011010011010_101_1_000110100110;
      patterns[13526] = 29'b0_011010011010_110_0_011010011010;
      patterns[13527] = 29'b0_011010011010_111_0_011010011010;
      patterns[13528] = 29'b0_011010011011_000_0_011010011011;
      patterns[13529] = 29'b0_011010011011_001_0_011011011010;
      patterns[13530] = 29'b0_011010011011_010_0_110100110110;
      patterns[13531] = 29'b0_011010011011_011_1_101001101100;
      patterns[13532] = 29'b0_011010011011_100_1_001101001101;
      patterns[13533] = 29'b0_011010011011_101_1_100110100110;
      patterns[13534] = 29'b0_011010011011_110_0_011010011011;
      patterns[13535] = 29'b0_011010011011_111_0_011010011011;
      patterns[13536] = 29'b0_011010011100_000_0_011010011100;
      patterns[13537] = 29'b0_011010011100_001_0_011100011010;
      patterns[13538] = 29'b0_011010011100_010_0_110100111000;
      patterns[13539] = 29'b0_011010011100_011_1_101001110000;
      patterns[13540] = 29'b0_011010011100_100_0_001101001110;
      patterns[13541] = 29'b0_011010011100_101_0_000110100111;
      patterns[13542] = 29'b0_011010011100_110_0_011010011100;
      patterns[13543] = 29'b0_011010011100_111_0_011010011100;
      patterns[13544] = 29'b0_011010011101_000_0_011010011101;
      patterns[13545] = 29'b0_011010011101_001_0_011101011010;
      patterns[13546] = 29'b0_011010011101_010_0_110100111010;
      patterns[13547] = 29'b0_011010011101_011_1_101001110100;
      patterns[13548] = 29'b0_011010011101_100_1_001101001110;
      patterns[13549] = 29'b0_011010011101_101_0_100110100111;
      patterns[13550] = 29'b0_011010011101_110_0_011010011101;
      patterns[13551] = 29'b0_011010011101_111_0_011010011101;
      patterns[13552] = 29'b0_011010011110_000_0_011010011110;
      patterns[13553] = 29'b0_011010011110_001_0_011110011010;
      patterns[13554] = 29'b0_011010011110_010_0_110100111100;
      patterns[13555] = 29'b0_011010011110_011_1_101001111000;
      patterns[13556] = 29'b0_011010011110_100_0_001101001111;
      patterns[13557] = 29'b0_011010011110_101_1_000110100111;
      patterns[13558] = 29'b0_011010011110_110_0_011010011110;
      patterns[13559] = 29'b0_011010011110_111_0_011010011110;
      patterns[13560] = 29'b0_011010011111_000_0_011010011111;
      patterns[13561] = 29'b0_011010011111_001_0_011111011010;
      patterns[13562] = 29'b0_011010011111_010_0_110100111110;
      patterns[13563] = 29'b0_011010011111_011_1_101001111100;
      patterns[13564] = 29'b0_011010011111_100_1_001101001111;
      patterns[13565] = 29'b0_011010011111_101_1_100110100111;
      patterns[13566] = 29'b0_011010011111_110_0_011010011111;
      patterns[13567] = 29'b0_011010011111_111_0_011010011111;
      patterns[13568] = 29'b0_011010100000_000_0_011010100000;
      patterns[13569] = 29'b0_011010100000_001_0_100000011010;
      patterns[13570] = 29'b0_011010100000_010_0_110101000000;
      patterns[13571] = 29'b0_011010100000_011_1_101010000000;
      patterns[13572] = 29'b0_011010100000_100_0_001101010000;
      patterns[13573] = 29'b0_011010100000_101_0_000110101000;
      patterns[13574] = 29'b0_011010100000_110_0_011010100000;
      patterns[13575] = 29'b0_011010100000_111_0_011010100000;
      patterns[13576] = 29'b0_011010100001_000_0_011010100001;
      patterns[13577] = 29'b0_011010100001_001_0_100001011010;
      patterns[13578] = 29'b0_011010100001_010_0_110101000010;
      patterns[13579] = 29'b0_011010100001_011_1_101010000100;
      patterns[13580] = 29'b0_011010100001_100_1_001101010000;
      patterns[13581] = 29'b0_011010100001_101_0_100110101000;
      patterns[13582] = 29'b0_011010100001_110_0_011010100001;
      patterns[13583] = 29'b0_011010100001_111_0_011010100001;
      patterns[13584] = 29'b0_011010100010_000_0_011010100010;
      patterns[13585] = 29'b0_011010100010_001_0_100010011010;
      patterns[13586] = 29'b0_011010100010_010_0_110101000100;
      patterns[13587] = 29'b0_011010100010_011_1_101010001000;
      patterns[13588] = 29'b0_011010100010_100_0_001101010001;
      patterns[13589] = 29'b0_011010100010_101_1_000110101000;
      patterns[13590] = 29'b0_011010100010_110_0_011010100010;
      patterns[13591] = 29'b0_011010100010_111_0_011010100010;
      patterns[13592] = 29'b0_011010100011_000_0_011010100011;
      patterns[13593] = 29'b0_011010100011_001_0_100011011010;
      patterns[13594] = 29'b0_011010100011_010_0_110101000110;
      patterns[13595] = 29'b0_011010100011_011_1_101010001100;
      patterns[13596] = 29'b0_011010100011_100_1_001101010001;
      patterns[13597] = 29'b0_011010100011_101_1_100110101000;
      patterns[13598] = 29'b0_011010100011_110_0_011010100011;
      patterns[13599] = 29'b0_011010100011_111_0_011010100011;
      patterns[13600] = 29'b0_011010100100_000_0_011010100100;
      patterns[13601] = 29'b0_011010100100_001_0_100100011010;
      patterns[13602] = 29'b0_011010100100_010_0_110101001000;
      patterns[13603] = 29'b0_011010100100_011_1_101010010000;
      patterns[13604] = 29'b0_011010100100_100_0_001101010010;
      patterns[13605] = 29'b0_011010100100_101_0_000110101001;
      patterns[13606] = 29'b0_011010100100_110_0_011010100100;
      patterns[13607] = 29'b0_011010100100_111_0_011010100100;
      patterns[13608] = 29'b0_011010100101_000_0_011010100101;
      patterns[13609] = 29'b0_011010100101_001_0_100101011010;
      patterns[13610] = 29'b0_011010100101_010_0_110101001010;
      patterns[13611] = 29'b0_011010100101_011_1_101010010100;
      patterns[13612] = 29'b0_011010100101_100_1_001101010010;
      patterns[13613] = 29'b0_011010100101_101_0_100110101001;
      patterns[13614] = 29'b0_011010100101_110_0_011010100101;
      patterns[13615] = 29'b0_011010100101_111_0_011010100101;
      patterns[13616] = 29'b0_011010100110_000_0_011010100110;
      patterns[13617] = 29'b0_011010100110_001_0_100110011010;
      patterns[13618] = 29'b0_011010100110_010_0_110101001100;
      patterns[13619] = 29'b0_011010100110_011_1_101010011000;
      patterns[13620] = 29'b0_011010100110_100_0_001101010011;
      patterns[13621] = 29'b0_011010100110_101_1_000110101001;
      patterns[13622] = 29'b0_011010100110_110_0_011010100110;
      patterns[13623] = 29'b0_011010100110_111_0_011010100110;
      patterns[13624] = 29'b0_011010100111_000_0_011010100111;
      patterns[13625] = 29'b0_011010100111_001_0_100111011010;
      patterns[13626] = 29'b0_011010100111_010_0_110101001110;
      patterns[13627] = 29'b0_011010100111_011_1_101010011100;
      patterns[13628] = 29'b0_011010100111_100_1_001101010011;
      patterns[13629] = 29'b0_011010100111_101_1_100110101001;
      patterns[13630] = 29'b0_011010100111_110_0_011010100111;
      patterns[13631] = 29'b0_011010100111_111_0_011010100111;
      patterns[13632] = 29'b0_011010101000_000_0_011010101000;
      patterns[13633] = 29'b0_011010101000_001_0_101000011010;
      patterns[13634] = 29'b0_011010101000_010_0_110101010000;
      patterns[13635] = 29'b0_011010101000_011_1_101010100000;
      patterns[13636] = 29'b0_011010101000_100_0_001101010100;
      patterns[13637] = 29'b0_011010101000_101_0_000110101010;
      patterns[13638] = 29'b0_011010101000_110_0_011010101000;
      patterns[13639] = 29'b0_011010101000_111_0_011010101000;
      patterns[13640] = 29'b0_011010101001_000_0_011010101001;
      patterns[13641] = 29'b0_011010101001_001_0_101001011010;
      patterns[13642] = 29'b0_011010101001_010_0_110101010010;
      patterns[13643] = 29'b0_011010101001_011_1_101010100100;
      patterns[13644] = 29'b0_011010101001_100_1_001101010100;
      patterns[13645] = 29'b0_011010101001_101_0_100110101010;
      patterns[13646] = 29'b0_011010101001_110_0_011010101001;
      patterns[13647] = 29'b0_011010101001_111_0_011010101001;
      patterns[13648] = 29'b0_011010101010_000_0_011010101010;
      patterns[13649] = 29'b0_011010101010_001_0_101010011010;
      patterns[13650] = 29'b0_011010101010_010_0_110101010100;
      patterns[13651] = 29'b0_011010101010_011_1_101010101000;
      patterns[13652] = 29'b0_011010101010_100_0_001101010101;
      patterns[13653] = 29'b0_011010101010_101_1_000110101010;
      patterns[13654] = 29'b0_011010101010_110_0_011010101010;
      patterns[13655] = 29'b0_011010101010_111_0_011010101010;
      patterns[13656] = 29'b0_011010101011_000_0_011010101011;
      patterns[13657] = 29'b0_011010101011_001_0_101011011010;
      patterns[13658] = 29'b0_011010101011_010_0_110101010110;
      patterns[13659] = 29'b0_011010101011_011_1_101010101100;
      patterns[13660] = 29'b0_011010101011_100_1_001101010101;
      patterns[13661] = 29'b0_011010101011_101_1_100110101010;
      patterns[13662] = 29'b0_011010101011_110_0_011010101011;
      patterns[13663] = 29'b0_011010101011_111_0_011010101011;
      patterns[13664] = 29'b0_011010101100_000_0_011010101100;
      patterns[13665] = 29'b0_011010101100_001_0_101100011010;
      patterns[13666] = 29'b0_011010101100_010_0_110101011000;
      patterns[13667] = 29'b0_011010101100_011_1_101010110000;
      patterns[13668] = 29'b0_011010101100_100_0_001101010110;
      patterns[13669] = 29'b0_011010101100_101_0_000110101011;
      patterns[13670] = 29'b0_011010101100_110_0_011010101100;
      patterns[13671] = 29'b0_011010101100_111_0_011010101100;
      patterns[13672] = 29'b0_011010101101_000_0_011010101101;
      patterns[13673] = 29'b0_011010101101_001_0_101101011010;
      patterns[13674] = 29'b0_011010101101_010_0_110101011010;
      patterns[13675] = 29'b0_011010101101_011_1_101010110100;
      patterns[13676] = 29'b0_011010101101_100_1_001101010110;
      patterns[13677] = 29'b0_011010101101_101_0_100110101011;
      patterns[13678] = 29'b0_011010101101_110_0_011010101101;
      patterns[13679] = 29'b0_011010101101_111_0_011010101101;
      patterns[13680] = 29'b0_011010101110_000_0_011010101110;
      patterns[13681] = 29'b0_011010101110_001_0_101110011010;
      patterns[13682] = 29'b0_011010101110_010_0_110101011100;
      patterns[13683] = 29'b0_011010101110_011_1_101010111000;
      patterns[13684] = 29'b0_011010101110_100_0_001101010111;
      patterns[13685] = 29'b0_011010101110_101_1_000110101011;
      patterns[13686] = 29'b0_011010101110_110_0_011010101110;
      patterns[13687] = 29'b0_011010101110_111_0_011010101110;
      patterns[13688] = 29'b0_011010101111_000_0_011010101111;
      patterns[13689] = 29'b0_011010101111_001_0_101111011010;
      patterns[13690] = 29'b0_011010101111_010_0_110101011110;
      patterns[13691] = 29'b0_011010101111_011_1_101010111100;
      patterns[13692] = 29'b0_011010101111_100_1_001101010111;
      patterns[13693] = 29'b0_011010101111_101_1_100110101011;
      patterns[13694] = 29'b0_011010101111_110_0_011010101111;
      patterns[13695] = 29'b0_011010101111_111_0_011010101111;
      patterns[13696] = 29'b0_011010110000_000_0_011010110000;
      patterns[13697] = 29'b0_011010110000_001_0_110000011010;
      patterns[13698] = 29'b0_011010110000_010_0_110101100000;
      patterns[13699] = 29'b0_011010110000_011_1_101011000000;
      patterns[13700] = 29'b0_011010110000_100_0_001101011000;
      patterns[13701] = 29'b0_011010110000_101_0_000110101100;
      patterns[13702] = 29'b0_011010110000_110_0_011010110000;
      patterns[13703] = 29'b0_011010110000_111_0_011010110000;
      patterns[13704] = 29'b0_011010110001_000_0_011010110001;
      patterns[13705] = 29'b0_011010110001_001_0_110001011010;
      patterns[13706] = 29'b0_011010110001_010_0_110101100010;
      patterns[13707] = 29'b0_011010110001_011_1_101011000100;
      patterns[13708] = 29'b0_011010110001_100_1_001101011000;
      patterns[13709] = 29'b0_011010110001_101_0_100110101100;
      patterns[13710] = 29'b0_011010110001_110_0_011010110001;
      patterns[13711] = 29'b0_011010110001_111_0_011010110001;
      patterns[13712] = 29'b0_011010110010_000_0_011010110010;
      patterns[13713] = 29'b0_011010110010_001_0_110010011010;
      patterns[13714] = 29'b0_011010110010_010_0_110101100100;
      patterns[13715] = 29'b0_011010110010_011_1_101011001000;
      patterns[13716] = 29'b0_011010110010_100_0_001101011001;
      patterns[13717] = 29'b0_011010110010_101_1_000110101100;
      patterns[13718] = 29'b0_011010110010_110_0_011010110010;
      patterns[13719] = 29'b0_011010110010_111_0_011010110010;
      patterns[13720] = 29'b0_011010110011_000_0_011010110011;
      patterns[13721] = 29'b0_011010110011_001_0_110011011010;
      patterns[13722] = 29'b0_011010110011_010_0_110101100110;
      patterns[13723] = 29'b0_011010110011_011_1_101011001100;
      patterns[13724] = 29'b0_011010110011_100_1_001101011001;
      patterns[13725] = 29'b0_011010110011_101_1_100110101100;
      patterns[13726] = 29'b0_011010110011_110_0_011010110011;
      patterns[13727] = 29'b0_011010110011_111_0_011010110011;
      patterns[13728] = 29'b0_011010110100_000_0_011010110100;
      patterns[13729] = 29'b0_011010110100_001_0_110100011010;
      patterns[13730] = 29'b0_011010110100_010_0_110101101000;
      patterns[13731] = 29'b0_011010110100_011_1_101011010000;
      patterns[13732] = 29'b0_011010110100_100_0_001101011010;
      patterns[13733] = 29'b0_011010110100_101_0_000110101101;
      patterns[13734] = 29'b0_011010110100_110_0_011010110100;
      patterns[13735] = 29'b0_011010110100_111_0_011010110100;
      patterns[13736] = 29'b0_011010110101_000_0_011010110101;
      patterns[13737] = 29'b0_011010110101_001_0_110101011010;
      patterns[13738] = 29'b0_011010110101_010_0_110101101010;
      patterns[13739] = 29'b0_011010110101_011_1_101011010100;
      patterns[13740] = 29'b0_011010110101_100_1_001101011010;
      patterns[13741] = 29'b0_011010110101_101_0_100110101101;
      patterns[13742] = 29'b0_011010110101_110_0_011010110101;
      patterns[13743] = 29'b0_011010110101_111_0_011010110101;
      patterns[13744] = 29'b0_011010110110_000_0_011010110110;
      patterns[13745] = 29'b0_011010110110_001_0_110110011010;
      patterns[13746] = 29'b0_011010110110_010_0_110101101100;
      patterns[13747] = 29'b0_011010110110_011_1_101011011000;
      patterns[13748] = 29'b0_011010110110_100_0_001101011011;
      patterns[13749] = 29'b0_011010110110_101_1_000110101101;
      patterns[13750] = 29'b0_011010110110_110_0_011010110110;
      patterns[13751] = 29'b0_011010110110_111_0_011010110110;
      patterns[13752] = 29'b0_011010110111_000_0_011010110111;
      patterns[13753] = 29'b0_011010110111_001_0_110111011010;
      patterns[13754] = 29'b0_011010110111_010_0_110101101110;
      patterns[13755] = 29'b0_011010110111_011_1_101011011100;
      patterns[13756] = 29'b0_011010110111_100_1_001101011011;
      patterns[13757] = 29'b0_011010110111_101_1_100110101101;
      patterns[13758] = 29'b0_011010110111_110_0_011010110111;
      patterns[13759] = 29'b0_011010110111_111_0_011010110111;
      patterns[13760] = 29'b0_011010111000_000_0_011010111000;
      patterns[13761] = 29'b0_011010111000_001_0_111000011010;
      patterns[13762] = 29'b0_011010111000_010_0_110101110000;
      patterns[13763] = 29'b0_011010111000_011_1_101011100000;
      patterns[13764] = 29'b0_011010111000_100_0_001101011100;
      patterns[13765] = 29'b0_011010111000_101_0_000110101110;
      patterns[13766] = 29'b0_011010111000_110_0_011010111000;
      patterns[13767] = 29'b0_011010111000_111_0_011010111000;
      patterns[13768] = 29'b0_011010111001_000_0_011010111001;
      patterns[13769] = 29'b0_011010111001_001_0_111001011010;
      patterns[13770] = 29'b0_011010111001_010_0_110101110010;
      patterns[13771] = 29'b0_011010111001_011_1_101011100100;
      patterns[13772] = 29'b0_011010111001_100_1_001101011100;
      patterns[13773] = 29'b0_011010111001_101_0_100110101110;
      patterns[13774] = 29'b0_011010111001_110_0_011010111001;
      patterns[13775] = 29'b0_011010111001_111_0_011010111001;
      patterns[13776] = 29'b0_011010111010_000_0_011010111010;
      patterns[13777] = 29'b0_011010111010_001_0_111010011010;
      patterns[13778] = 29'b0_011010111010_010_0_110101110100;
      patterns[13779] = 29'b0_011010111010_011_1_101011101000;
      patterns[13780] = 29'b0_011010111010_100_0_001101011101;
      patterns[13781] = 29'b0_011010111010_101_1_000110101110;
      patterns[13782] = 29'b0_011010111010_110_0_011010111010;
      patterns[13783] = 29'b0_011010111010_111_0_011010111010;
      patterns[13784] = 29'b0_011010111011_000_0_011010111011;
      patterns[13785] = 29'b0_011010111011_001_0_111011011010;
      patterns[13786] = 29'b0_011010111011_010_0_110101110110;
      patterns[13787] = 29'b0_011010111011_011_1_101011101100;
      patterns[13788] = 29'b0_011010111011_100_1_001101011101;
      patterns[13789] = 29'b0_011010111011_101_1_100110101110;
      patterns[13790] = 29'b0_011010111011_110_0_011010111011;
      patterns[13791] = 29'b0_011010111011_111_0_011010111011;
      patterns[13792] = 29'b0_011010111100_000_0_011010111100;
      patterns[13793] = 29'b0_011010111100_001_0_111100011010;
      patterns[13794] = 29'b0_011010111100_010_0_110101111000;
      patterns[13795] = 29'b0_011010111100_011_1_101011110000;
      patterns[13796] = 29'b0_011010111100_100_0_001101011110;
      patterns[13797] = 29'b0_011010111100_101_0_000110101111;
      patterns[13798] = 29'b0_011010111100_110_0_011010111100;
      patterns[13799] = 29'b0_011010111100_111_0_011010111100;
      patterns[13800] = 29'b0_011010111101_000_0_011010111101;
      patterns[13801] = 29'b0_011010111101_001_0_111101011010;
      patterns[13802] = 29'b0_011010111101_010_0_110101111010;
      patterns[13803] = 29'b0_011010111101_011_1_101011110100;
      patterns[13804] = 29'b0_011010111101_100_1_001101011110;
      patterns[13805] = 29'b0_011010111101_101_0_100110101111;
      patterns[13806] = 29'b0_011010111101_110_0_011010111101;
      patterns[13807] = 29'b0_011010111101_111_0_011010111101;
      patterns[13808] = 29'b0_011010111110_000_0_011010111110;
      patterns[13809] = 29'b0_011010111110_001_0_111110011010;
      patterns[13810] = 29'b0_011010111110_010_0_110101111100;
      patterns[13811] = 29'b0_011010111110_011_1_101011111000;
      patterns[13812] = 29'b0_011010111110_100_0_001101011111;
      patterns[13813] = 29'b0_011010111110_101_1_000110101111;
      patterns[13814] = 29'b0_011010111110_110_0_011010111110;
      patterns[13815] = 29'b0_011010111110_111_0_011010111110;
      patterns[13816] = 29'b0_011010111111_000_0_011010111111;
      patterns[13817] = 29'b0_011010111111_001_0_111111011010;
      patterns[13818] = 29'b0_011010111111_010_0_110101111110;
      patterns[13819] = 29'b0_011010111111_011_1_101011111100;
      patterns[13820] = 29'b0_011010111111_100_1_001101011111;
      patterns[13821] = 29'b0_011010111111_101_1_100110101111;
      patterns[13822] = 29'b0_011010111111_110_0_011010111111;
      patterns[13823] = 29'b0_011010111111_111_0_011010111111;
      patterns[13824] = 29'b0_011011000000_000_0_011011000000;
      patterns[13825] = 29'b0_011011000000_001_0_000000011011;
      patterns[13826] = 29'b0_011011000000_010_0_110110000000;
      patterns[13827] = 29'b0_011011000000_011_1_101100000000;
      patterns[13828] = 29'b0_011011000000_100_0_001101100000;
      patterns[13829] = 29'b0_011011000000_101_0_000110110000;
      patterns[13830] = 29'b0_011011000000_110_0_011011000000;
      patterns[13831] = 29'b0_011011000000_111_0_011011000000;
      patterns[13832] = 29'b0_011011000001_000_0_011011000001;
      patterns[13833] = 29'b0_011011000001_001_0_000001011011;
      patterns[13834] = 29'b0_011011000001_010_0_110110000010;
      patterns[13835] = 29'b0_011011000001_011_1_101100000100;
      patterns[13836] = 29'b0_011011000001_100_1_001101100000;
      patterns[13837] = 29'b0_011011000001_101_0_100110110000;
      patterns[13838] = 29'b0_011011000001_110_0_011011000001;
      patterns[13839] = 29'b0_011011000001_111_0_011011000001;
      patterns[13840] = 29'b0_011011000010_000_0_011011000010;
      patterns[13841] = 29'b0_011011000010_001_0_000010011011;
      patterns[13842] = 29'b0_011011000010_010_0_110110000100;
      patterns[13843] = 29'b0_011011000010_011_1_101100001000;
      patterns[13844] = 29'b0_011011000010_100_0_001101100001;
      patterns[13845] = 29'b0_011011000010_101_1_000110110000;
      patterns[13846] = 29'b0_011011000010_110_0_011011000010;
      patterns[13847] = 29'b0_011011000010_111_0_011011000010;
      patterns[13848] = 29'b0_011011000011_000_0_011011000011;
      patterns[13849] = 29'b0_011011000011_001_0_000011011011;
      patterns[13850] = 29'b0_011011000011_010_0_110110000110;
      patterns[13851] = 29'b0_011011000011_011_1_101100001100;
      patterns[13852] = 29'b0_011011000011_100_1_001101100001;
      patterns[13853] = 29'b0_011011000011_101_1_100110110000;
      patterns[13854] = 29'b0_011011000011_110_0_011011000011;
      patterns[13855] = 29'b0_011011000011_111_0_011011000011;
      patterns[13856] = 29'b0_011011000100_000_0_011011000100;
      patterns[13857] = 29'b0_011011000100_001_0_000100011011;
      patterns[13858] = 29'b0_011011000100_010_0_110110001000;
      patterns[13859] = 29'b0_011011000100_011_1_101100010000;
      patterns[13860] = 29'b0_011011000100_100_0_001101100010;
      patterns[13861] = 29'b0_011011000100_101_0_000110110001;
      patterns[13862] = 29'b0_011011000100_110_0_011011000100;
      patterns[13863] = 29'b0_011011000100_111_0_011011000100;
      patterns[13864] = 29'b0_011011000101_000_0_011011000101;
      patterns[13865] = 29'b0_011011000101_001_0_000101011011;
      patterns[13866] = 29'b0_011011000101_010_0_110110001010;
      patterns[13867] = 29'b0_011011000101_011_1_101100010100;
      patterns[13868] = 29'b0_011011000101_100_1_001101100010;
      patterns[13869] = 29'b0_011011000101_101_0_100110110001;
      patterns[13870] = 29'b0_011011000101_110_0_011011000101;
      patterns[13871] = 29'b0_011011000101_111_0_011011000101;
      patterns[13872] = 29'b0_011011000110_000_0_011011000110;
      patterns[13873] = 29'b0_011011000110_001_0_000110011011;
      patterns[13874] = 29'b0_011011000110_010_0_110110001100;
      patterns[13875] = 29'b0_011011000110_011_1_101100011000;
      patterns[13876] = 29'b0_011011000110_100_0_001101100011;
      patterns[13877] = 29'b0_011011000110_101_1_000110110001;
      patterns[13878] = 29'b0_011011000110_110_0_011011000110;
      patterns[13879] = 29'b0_011011000110_111_0_011011000110;
      patterns[13880] = 29'b0_011011000111_000_0_011011000111;
      patterns[13881] = 29'b0_011011000111_001_0_000111011011;
      patterns[13882] = 29'b0_011011000111_010_0_110110001110;
      patterns[13883] = 29'b0_011011000111_011_1_101100011100;
      patterns[13884] = 29'b0_011011000111_100_1_001101100011;
      patterns[13885] = 29'b0_011011000111_101_1_100110110001;
      patterns[13886] = 29'b0_011011000111_110_0_011011000111;
      patterns[13887] = 29'b0_011011000111_111_0_011011000111;
      patterns[13888] = 29'b0_011011001000_000_0_011011001000;
      patterns[13889] = 29'b0_011011001000_001_0_001000011011;
      patterns[13890] = 29'b0_011011001000_010_0_110110010000;
      patterns[13891] = 29'b0_011011001000_011_1_101100100000;
      patterns[13892] = 29'b0_011011001000_100_0_001101100100;
      patterns[13893] = 29'b0_011011001000_101_0_000110110010;
      patterns[13894] = 29'b0_011011001000_110_0_011011001000;
      patterns[13895] = 29'b0_011011001000_111_0_011011001000;
      patterns[13896] = 29'b0_011011001001_000_0_011011001001;
      patterns[13897] = 29'b0_011011001001_001_0_001001011011;
      patterns[13898] = 29'b0_011011001001_010_0_110110010010;
      patterns[13899] = 29'b0_011011001001_011_1_101100100100;
      patterns[13900] = 29'b0_011011001001_100_1_001101100100;
      patterns[13901] = 29'b0_011011001001_101_0_100110110010;
      patterns[13902] = 29'b0_011011001001_110_0_011011001001;
      patterns[13903] = 29'b0_011011001001_111_0_011011001001;
      patterns[13904] = 29'b0_011011001010_000_0_011011001010;
      patterns[13905] = 29'b0_011011001010_001_0_001010011011;
      patterns[13906] = 29'b0_011011001010_010_0_110110010100;
      patterns[13907] = 29'b0_011011001010_011_1_101100101000;
      patterns[13908] = 29'b0_011011001010_100_0_001101100101;
      patterns[13909] = 29'b0_011011001010_101_1_000110110010;
      patterns[13910] = 29'b0_011011001010_110_0_011011001010;
      patterns[13911] = 29'b0_011011001010_111_0_011011001010;
      patterns[13912] = 29'b0_011011001011_000_0_011011001011;
      patterns[13913] = 29'b0_011011001011_001_0_001011011011;
      patterns[13914] = 29'b0_011011001011_010_0_110110010110;
      patterns[13915] = 29'b0_011011001011_011_1_101100101100;
      patterns[13916] = 29'b0_011011001011_100_1_001101100101;
      patterns[13917] = 29'b0_011011001011_101_1_100110110010;
      patterns[13918] = 29'b0_011011001011_110_0_011011001011;
      patterns[13919] = 29'b0_011011001011_111_0_011011001011;
      patterns[13920] = 29'b0_011011001100_000_0_011011001100;
      patterns[13921] = 29'b0_011011001100_001_0_001100011011;
      patterns[13922] = 29'b0_011011001100_010_0_110110011000;
      patterns[13923] = 29'b0_011011001100_011_1_101100110000;
      patterns[13924] = 29'b0_011011001100_100_0_001101100110;
      patterns[13925] = 29'b0_011011001100_101_0_000110110011;
      patterns[13926] = 29'b0_011011001100_110_0_011011001100;
      patterns[13927] = 29'b0_011011001100_111_0_011011001100;
      patterns[13928] = 29'b0_011011001101_000_0_011011001101;
      patterns[13929] = 29'b0_011011001101_001_0_001101011011;
      patterns[13930] = 29'b0_011011001101_010_0_110110011010;
      patterns[13931] = 29'b0_011011001101_011_1_101100110100;
      patterns[13932] = 29'b0_011011001101_100_1_001101100110;
      patterns[13933] = 29'b0_011011001101_101_0_100110110011;
      patterns[13934] = 29'b0_011011001101_110_0_011011001101;
      patterns[13935] = 29'b0_011011001101_111_0_011011001101;
      patterns[13936] = 29'b0_011011001110_000_0_011011001110;
      patterns[13937] = 29'b0_011011001110_001_0_001110011011;
      patterns[13938] = 29'b0_011011001110_010_0_110110011100;
      patterns[13939] = 29'b0_011011001110_011_1_101100111000;
      patterns[13940] = 29'b0_011011001110_100_0_001101100111;
      patterns[13941] = 29'b0_011011001110_101_1_000110110011;
      patterns[13942] = 29'b0_011011001110_110_0_011011001110;
      patterns[13943] = 29'b0_011011001110_111_0_011011001110;
      patterns[13944] = 29'b0_011011001111_000_0_011011001111;
      patterns[13945] = 29'b0_011011001111_001_0_001111011011;
      patterns[13946] = 29'b0_011011001111_010_0_110110011110;
      patterns[13947] = 29'b0_011011001111_011_1_101100111100;
      patterns[13948] = 29'b0_011011001111_100_1_001101100111;
      patterns[13949] = 29'b0_011011001111_101_1_100110110011;
      patterns[13950] = 29'b0_011011001111_110_0_011011001111;
      patterns[13951] = 29'b0_011011001111_111_0_011011001111;
      patterns[13952] = 29'b0_011011010000_000_0_011011010000;
      patterns[13953] = 29'b0_011011010000_001_0_010000011011;
      patterns[13954] = 29'b0_011011010000_010_0_110110100000;
      patterns[13955] = 29'b0_011011010000_011_1_101101000000;
      patterns[13956] = 29'b0_011011010000_100_0_001101101000;
      patterns[13957] = 29'b0_011011010000_101_0_000110110100;
      patterns[13958] = 29'b0_011011010000_110_0_011011010000;
      patterns[13959] = 29'b0_011011010000_111_0_011011010000;
      patterns[13960] = 29'b0_011011010001_000_0_011011010001;
      patterns[13961] = 29'b0_011011010001_001_0_010001011011;
      patterns[13962] = 29'b0_011011010001_010_0_110110100010;
      patterns[13963] = 29'b0_011011010001_011_1_101101000100;
      patterns[13964] = 29'b0_011011010001_100_1_001101101000;
      patterns[13965] = 29'b0_011011010001_101_0_100110110100;
      patterns[13966] = 29'b0_011011010001_110_0_011011010001;
      patterns[13967] = 29'b0_011011010001_111_0_011011010001;
      patterns[13968] = 29'b0_011011010010_000_0_011011010010;
      patterns[13969] = 29'b0_011011010010_001_0_010010011011;
      patterns[13970] = 29'b0_011011010010_010_0_110110100100;
      patterns[13971] = 29'b0_011011010010_011_1_101101001000;
      patterns[13972] = 29'b0_011011010010_100_0_001101101001;
      patterns[13973] = 29'b0_011011010010_101_1_000110110100;
      patterns[13974] = 29'b0_011011010010_110_0_011011010010;
      patterns[13975] = 29'b0_011011010010_111_0_011011010010;
      patterns[13976] = 29'b0_011011010011_000_0_011011010011;
      patterns[13977] = 29'b0_011011010011_001_0_010011011011;
      patterns[13978] = 29'b0_011011010011_010_0_110110100110;
      patterns[13979] = 29'b0_011011010011_011_1_101101001100;
      patterns[13980] = 29'b0_011011010011_100_1_001101101001;
      patterns[13981] = 29'b0_011011010011_101_1_100110110100;
      patterns[13982] = 29'b0_011011010011_110_0_011011010011;
      patterns[13983] = 29'b0_011011010011_111_0_011011010011;
      patterns[13984] = 29'b0_011011010100_000_0_011011010100;
      patterns[13985] = 29'b0_011011010100_001_0_010100011011;
      patterns[13986] = 29'b0_011011010100_010_0_110110101000;
      patterns[13987] = 29'b0_011011010100_011_1_101101010000;
      patterns[13988] = 29'b0_011011010100_100_0_001101101010;
      patterns[13989] = 29'b0_011011010100_101_0_000110110101;
      patterns[13990] = 29'b0_011011010100_110_0_011011010100;
      patterns[13991] = 29'b0_011011010100_111_0_011011010100;
      patterns[13992] = 29'b0_011011010101_000_0_011011010101;
      patterns[13993] = 29'b0_011011010101_001_0_010101011011;
      patterns[13994] = 29'b0_011011010101_010_0_110110101010;
      patterns[13995] = 29'b0_011011010101_011_1_101101010100;
      patterns[13996] = 29'b0_011011010101_100_1_001101101010;
      patterns[13997] = 29'b0_011011010101_101_0_100110110101;
      patterns[13998] = 29'b0_011011010101_110_0_011011010101;
      patterns[13999] = 29'b0_011011010101_111_0_011011010101;
      patterns[14000] = 29'b0_011011010110_000_0_011011010110;
      patterns[14001] = 29'b0_011011010110_001_0_010110011011;
      patterns[14002] = 29'b0_011011010110_010_0_110110101100;
      patterns[14003] = 29'b0_011011010110_011_1_101101011000;
      patterns[14004] = 29'b0_011011010110_100_0_001101101011;
      patterns[14005] = 29'b0_011011010110_101_1_000110110101;
      patterns[14006] = 29'b0_011011010110_110_0_011011010110;
      patterns[14007] = 29'b0_011011010110_111_0_011011010110;
      patterns[14008] = 29'b0_011011010111_000_0_011011010111;
      patterns[14009] = 29'b0_011011010111_001_0_010111011011;
      patterns[14010] = 29'b0_011011010111_010_0_110110101110;
      patterns[14011] = 29'b0_011011010111_011_1_101101011100;
      patterns[14012] = 29'b0_011011010111_100_1_001101101011;
      patterns[14013] = 29'b0_011011010111_101_1_100110110101;
      patterns[14014] = 29'b0_011011010111_110_0_011011010111;
      patterns[14015] = 29'b0_011011010111_111_0_011011010111;
      patterns[14016] = 29'b0_011011011000_000_0_011011011000;
      patterns[14017] = 29'b0_011011011000_001_0_011000011011;
      patterns[14018] = 29'b0_011011011000_010_0_110110110000;
      patterns[14019] = 29'b0_011011011000_011_1_101101100000;
      patterns[14020] = 29'b0_011011011000_100_0_001101101100;
      patterns[14021] = 29'b0_011011011000_101_0_000110110110;
      patterns[14022] = 29'b0_011011011000_110_0_011011011000;
      patterns[14023] = 29'b0_011011011000_111_0_011011011000;
      patterns[14024] = 29'b0_011011011001_000_0_011011011001;
      patterns[14025] = 29'b0_011011011001_001_0_011001011011;
      patterns[14026] = 29'b0_011011011001_010_0_110110110010;
      patterns[14027] = 29'b0_011011011001_011_1_101101100100;
      patterns[14028] = 29'b0_011011011001_100_1_001101101100;
      patterns[14029] = 29'b0_011011011001_101_0_100110110110;
      patterns[14030] = 29'b0_011011011001_110_0_011011011001;
      patterns[14031] = 29'b0_011011011001_111_0_011011011001;
      patterns[14032] = 29'b0_011011011010_000_0_011011011010;
      patterns[14033] = 29'b0_011011011010_001_0_011010011011;
      patterns[14034] = 29'b0_011011011010_010_0_110110110100;
      patterns[14035] = 29'b0_011011011010_011_1_101101101000;
      patterns[14036] = 29'b0_011011011010_100_0_001101101101;
      patterns[14037] = 29'b0_011011011010_101_1_000110110110;
      patterns[14038] = 29'b0_011011011010_110_0_011011011010;
      patterns[14039] = 29'b0_011011011010_111_0_011011011010;
      patterns[14040] = 29'b0_011011011011_000_0_011011011011;
      patterns[14041] = 29'b0_011011011011_001_0_011011011011;
      patterns[14042] = 29'b0_011011011011_010_0_110110110110;
      patterns[14043] = 29'b0_011011011011_011_1_101101101100;
      patterns[14044] = 29'b0_011011011011_100_1_001101101101;
      patterns[14045] = 29'b0_011011011011_101_1_100110110110;
      patterns[14046] = 29'b0_011011011011_110_0_011011011011;
      patterns[14047] = 29'b0_011011011011_111_0_011011011011;
      patterns[14048] = 29'b0_011011011100_000_0_011011011100;
      patterns[14049] = 29'b0_011011011100_001_0_011100011011;
      patterns[14050] = 29'b0_011011011100_010_0_110110111000;
      patterns[14051] = 29'b0_011011011100_011_1_101101110000;
      patterns[14052] = 29'b0_011011011100_100_0_001101101110;
      patterns[14053] = 29'b0_011011011100_101_0_000110110111;
      patterns[14054] = 29'b0_011011011100_110_0_011011011100;
      patterns[14055] = 29'b0_011011011100_111_0_011011011100;
      patterns[14056] = 29'b0_011011011101_000_0_011011011101;
      patterns[14057] = 29'b0_011011011101_001_0_011101011011;
      patterns[14058] = 29'b0_011011011101_010_0_110110111010;
      patterns[14059] = 29'b0_011011011101_011_1_101101110100;
      patterns[14060] = 29'b0_011011011101_100_1_001101101110;
      patterns[14061] = 29'b0_011011011101_101_0_100110110111;
      patterns[14062] = 29'b0_011011011101_110_0_011011011101;
      patterns[14063] = 29'b0_011011011101_111_0_011011011101;
      patterns[14064] = 29'b0_011011011110_000_0_011011011110;
      patterns[14065] = 29'b0_011011011110_001_0_011110011011;
      patterns[14066] = 29'b0_011011011110_010_0_110110111100;
      patterns[14067] = 29'b0_011011011110_011_1_101101111000;
      patterns[14068] = 29'b0_011011011110_100_0_001101101111;
      patterns[14069] = 29'b0_011011011110_101_1_000110110111;
      patterns[14070] = 29'b0_011011011110_110_0_011011011110;
      patterns[14071] = 29'b0_011011011110_111_0_011011011110;
      patterns[14072] = 29'b0_011011011111_000_0_011011011111;
      patterns[14073] = 29'b0_011011011111_001_0_011111011011;
      patterns[14074] = 29'b0_011011011111_010_0_110110111110;
      patterns[14075] = 29'b0_011011011111_011_1_101101111100;
      patterns[14076] = 29'b0_011011011111_100_1_001101101111;
      patterns[14077] = 29'b0_011011011111_101_1_100110110111;
      patterns[14078] = 29'b0_011011011111_110_0_011011011111;
      patterns[14079] = 29'b0_011011011111_111_0_011011011111;
      patterns[14080] = 29'b0_011011100000_000_0_011011100000;
      patterns[14081] = 29'b0_011011100000_001_0_100000011011;
      patterns[14082] = 29'b0_011011100000_010_0_110111000000;
      patterns[14083] = 29'b0_011011100000_011_1_101110000000;
      patterns[14084] = 29'b0_011011100000_100_0_001101110000;
      patterns[14085] = 29'b0_011011100000_101_0_000110111000;
      patterns[14086] = 29'b0_011011100000_110_0_011011100000;
      patterns[14087] = 29'b0_011011100000_111_0_011011100000;
      patterns[14088] = 29'b0_011011100001_000_0_011011100001;
      patterns[14089] = 29'b0_011011100001_001_0_100001011011;
      patterns[14090] = 29'b0_011011100001_010_0_110111000010;
      patterns[14091] = 29'b0_011011100001_011_1_101110000100;
      patterns[14092] = 29'b0_011011100001_100_1_001101110000;
      patterns[14093] = 29'b0_011011100001_101_0_100110111000;
      patterns[14094] = 29'b0_011011100001_110_0_011011100001;
      patterns[14095] = 29'b0_011011100001_111_0_011011100001;
      patterns[14096] = 29'b0_011011100010_000_0_011011100010;
      patterns[14097] = 29'b0_011011100010_001_0_100010011011;
      patterns[14098] = 29'b0_011011100010_010_0_110111000100;
      patterns[14099] = 29'b0_011011100010_011_1_101110001000;
      patterns[14100] = 29'b0_011011100010_100_0_001101110001;
      patterns[14101] = 29'b0_011011100010_101_1_000110111000;
      patterns[14102] = 29'b0_011011100010_110_0_011011100010;
      patterns[14103] = 29'b0_011011100010_111_0_011011100010;
      patterns[14104] = 29'b0_011011100011_000_0_011011100011;
      patterns[14105] = 29'b0_011011100011_001_0_100011011011;
      patterns[14106] = 29'b0_011011100011_010_0_110111000110;
      patterns[14107] = 29'b0_011011100011_011_1_101110001100;
      patterns[14108] = 29'b0_011011100011_100_1_001101110001;
      patterns[14109] = 29'b0_011011100011_101_1_100110111000;
      patterns[14110] = 29'b0_011011100011_110_0_011011100011;
      patterns[14111] = 29'b0_011011100011_111_0_011011100011;
      patterns[14112] = 29'b0_011011100100_000_0_011011100100;
      patterns[14113] = 29'b0_011011100100_001_0_100100011011;
      patterns[14114] = 29'b0_011011100100_010_0_110111001000;
      patterns[14115] = 29'b0_011011100100_011_1_101110010000;
      patterns[14116] = 29'b0_011011100100_100_0_001101110010;
      patterns[14117] = 29'b0_011011100100_101_0_000110111001;
      patterns[14118] = 29'b0_011011100100_110_0_011011100100;
      patterns[14119] = 29'b0_011011100100_111_0_011011100100;
      patterns[14120] = 29'b0_011011100101_000_0_011011100101;
      patterns[14121] = 29'b0_011011100101_001_0_100101011011;
      patterns[14122] = 29'b0_011011100101_010_0_110111001010;
      patterns[14123] = 29'b0_011011100101_011_1_101110010100;
      patterns[14124] = 29'b0_011011100101_100_1_001101110010;
      patterns[14125] = 29'b0_011011100101_101_0_100110111001;
      patterns[14126] = 29'b0_011011100101_110_0_011011100101;
      patterns[14127] = 29'b0_011011100101_111_0_011011100101;
      patterns[14128] = 29'b0_011011100110_000_0_011011100110;
      patterns[14129] = 29'b0_011011100110_001_0_100110011011;
      patterns[14130] = 29'b0_011011100110_010_0_110111001100;
      patterns[14131] = 29'b0_011011100110_011_1_101110011000;
      patterns[14132] = 29'b0_011011100110_100_0_001101110011;
      patterns[14133] = 29'b0_011011100110_101_1_000110111001;
      patterns[14134] = 29'b0_011011100110_110_0_011011100110;
      patterns[14135] = 29'b0_011011100110_111_0_011011100110;
      patterns[14136] = 29'b0_011011100111_000_0_011011100111;
      patterns[14137] = 29'b0_011011100111_001_0_100111011011;
      patterns[14138] = 29'b0_011011100111_010_0_110111001110;
      patterns[14139] = 29'b0_011011100111_011_1_101110011100;
      patterns[14140] = 29'b0_011011100111_100_1_001101110011;
      patterns[14141] = 29'b0_011011100111_101_1_100110111001;
      patterns[14142] = 29'b0_011011100111_110_0_011011100111;
      patterns[14143] = 29'b0_011011100111_111_0_011011100111;
      patterns[14144] = 29'b0_011011101000_000_0_011011101000;
      patterns[14145] = 29'b0_011011101000_001_0_101000011011;
      patterns[14146] = 29'b0_011011101000_010_0_110111010000;
      patterns[14147] = 29'b0_011011101000_011_1_101110100000;
      patterns[14148] = 29'b0_011011101000_100_0_001101110100;
      patterns[14149] = 29'b0_011011101000_101_0_000110111010;
      patterns[14150] = 29'b0_011011101000_110_0_011011101000;
      patterns[14151] = 29'b0_011011101000_111_0_011011101000;
      patterns[14152] = 29'b0_011011101001_000_0_011011101001;
      patterns[14153] = 29'b0_011011101001_001_0_101001011011;
      patterns[14154] = 29'b0_011011101001_010_0_110111010010;
      patterns[14155] = 29'b0_011011101001_011_1_101110100100;
      patterns[14156] = 29'b0_011011101001_100_1_001101110100;
      patterns[14157] = 29'b0_011011101001_101_0_100110111010;
      patterns[14158] = 29'b0_011011101001_110_0_011011101001;
      patterns[14159] = 29'b0_011011101001_111_0_011011101001;
      patterns[14160] = 29'b0_011011101010_000_0_011011101010;
      patterns[14161] = 29'b0_011011101010_001_0_101010011011;
      patterns[14162] = 29'b0_011011101010_010_0_110111010100;
      patterns[14163] = 29'b0_011011101010_011_1_101110101000;
      patterns[14164] = 29'b0_011011101010_100_0_001101110101;
      patterns[14165] = 29'b0_011011101010_101_1_000110111010;
      patterns[14166] = 29'b0_011011101010_110_0_011011101010;
      patterns[14167] = 29'b0_011011101010_111_0_011011101010;
      patterns[14168] = 29'b0_011011101011_000_0_011011101011;
      patterns[14169] = 29'b0_011011101011_001_0_101011011011;
      patterns[14170] = 29'b0_011011101011_010_0_110111010110;
      patterns[14171] = 29'b0_011011101011_011_1_101110101100;
      patterns[14172] = 29'b0_011011101011_100_1_001101110101;
      patterns[14173] = 29'b0_011011101011_101_1_100110111010;
      patterns[14174] = 29'b0_011011101011_110_0_011011101011;
      patterns[14175] = 29'b0_011011101011_111_0_011011101011;
      patterns[14176] = 29'b0_011011101100_000_0_011011101100;
      patterns[14177] = 29'b0_011011101100_001_0_101100011011;
      patterns[14178] = 29'b0_011011101100_010_0_110111011000;
      patterns[14179] = 29'b0_011011101100_011_1_101110110000;
      patterns[14180] = 29'b0_011011101100_100_0_001101110110;
      patterns[14181] = 29'b0_011011101100_101_0_000110111011;
      patterns[14182] = 29'b0_011011101100_110_0_011011101100;
      patterns[14183] = 29'b0_011011101100_111_0_011011101100;
      patterns[14184] = 29'b0_011011101101_000_0_011011101101;
      patterns[14185] = 29'b0_011011101101_001_0_101101011011;
      patterns[14186] = 29'b0_011011101101_010_0_110111011010;
      patterns[14187] = 29'b0_011011101101_011_1_101110110100;
      patterns[14188] = 29'b0_011011101101_100_1_001101110110;
      patterns[14189] = 29'b0_011011101101_101_0_100110111011;
      patterns[14190] = 29'b0_011011101101_110_0_011011101101;
      patterns[14191] = 29'b0_011011101101_111_0_011011101101;
      patterns[14192] = 29'b0_011011101110_000_0_011011101110;
      patterns[14193] = 29'b0_011011101110_001_0_101110011011;
      patterns[14194] = 29'b0_011011101110_010_0_110111011100;
      patterns[14195] = 29'b0_011011101110_011_1_101110111000;
      patterns[14196] = 29'b0_011011101110_100_0_001101110111;
      patterns[14197] = 29'b0_011011101110_101_1_000110111011;
      patterns[14198] = 29'b0_011011101110_110_0_011011101110;
      patterns[14199] = 29'b0_011011101110_111_0_011011101110;
      patterns[14200] = 29'b0_011011101111_000_0_011011101111;
      patterns[14201] = 29'b0_011011101111_001_0_101111011011;
      patterns[14202] = 29'b0_011011101111_010_0_110111011110;
      patterns[14203] = 29'b0_011011101111_011_1_101110111100;
      patterns[14204] = 29'b0_011011101111_100_1_001101110111;
      patterns[14205] = 29'b0_011011101111_101_1_100110111011;
      patterns[14206] = 29'b0_011011101111_110_0_011011101111;
      patterns[14207] = 29'b0_011011101111_111_0_011011101111;
      patterns[14208] = 29'b0_011011110000_000_0_011011110000;
      patterns[14209] = 29'b0_011011110000_001_0_110000011011;
      patterns[14210] = 29'b0_011011110000_010_0_110111100000;
      patterns[14211] = 29'b0_011011110000_011_1_101111000000;
      patterns[14212] = 29'b0_011011110000_100_0_001101111000;
      patterns[14213] = 29'b0_011011110000_101_0_000110111100;
      patterns[14214] = 29'b0_011011110000_110_0_011011110000;
      patterns[14215] = 29'b0_011011110000_111_0_011011110000;
      patterns[14216] = 29'b0_011011110001_000_0_011011110001;
      patterns[14217] = 29'b0_011011110001_001_0_110001011011;
      patterns[14218] = 29'b0_011011110001_010_0_110111100010;
      patterns[14219] = 29'b0_011011110001_011_1_101111000100;
      patterns[14220] = 29'b0_011011110001_100_1_001101111000;
      patterns[14221] = 29'b0_011011110001_101_0_100110111100;
      patterns[14222] = 29'b0_011011110001_110_0_011011110001;
      patterns[14223] = 29'b0_011011110001_111_0_011011110001;
      patterns[14224] = 29'b0_011011110010_000_0_011011110010;
      patterns[14225] = 29'b0_011011110010_001_0_110010011011;
      patterns[14226] = 29'b0_011011110010_010_0_110111100100;
      patterns[14227] = 29'b0_011011110010_011_1_101111001000;
      patterns[14228] = 29'b0_011011110010_100_0_001101111001;
      patterns[14229] = 29'b0_011011110010_101_1_000110111100;
      patterns[14230] = 29'b0_011011110010_110_0_011011110010;
      patterns[14231] = 29'b0_011011110010_111_0_011011110010;
      patterns[14232] = 29'b0_011011110011_000_0_011011110011;
      patterns[14233] = 29'b0_011011110011_001_0_110011011011;
      patterns[14234] = 29'b0_011011110011_010_0_110111100110;
      patterns[14235] = 29'b0_011011110011_011_1_101111001100;
      patterns[14236] = 29'b0_011011110011_100_1_001101111001;
      patterns[14237] = 29'b0_011011110011_101_1_100110111100;
      patterns[14238] = 29'b0_011011110011_110_0_011011110011;
      patterns[14239] = 29'b0_011011110011_111_0_011011110011;
      patterns[14240] = 29'b0_011011110100_000_0_011011110100;
      patterns[14241] = 29'b0_011011110100_001_0_110100011011;
      patterns[14242] = 29'b0_011011110100_010_0_110111101000;
      patterns[14243] = 29'b0_011011110100_011_1_101111010000;
      patterns[14244] = 29'b0_011011110100_100_0_001101111010;
      patterns[14245] = 29'b0_011011110100_101_0_000110111101;
      patterns[14246] = 29'b0_011011110100_110_0_011011110100;
      patterns[14247] = 29'b0_011011110100_111_0_011011110100;
      patterns[14248] = 29'b0_011011110101_000_0_011011110101;
      patterns[14249] = 29'b0_011011110101_001_0_110101011011;
      patterns[14250] = 29'b0_011011110101_010_0_110111101010;
      patterns[14251] = 29'b0_011011110101_011_1_101111010100;
      patterns[14252] = 29'b0_011011110101_100_1_001101111010;
      patterns[14253] = 29'b0_011011110101_101_0_100110111101;
      patterns[14254] = 29'b0_011011110101_110_0_011011110101;
      patterns[14255] = 29'b0_011011110101_111_0_011011110101;
      patterns[14256] = 29'b0_011011110110_000_0_011011110110;
      patterns[14257] = 29'b0_011011110110_001_0_110110011011;
      patterns[14258] = 29'b0_011011110110_010_0_110111101100;
      patterns[14259] = 29'b0_011011110110_011_1_101111011000;
      patterns[14260] = 29'b0_011011110110_100_0_001101111011;
      patterns[14261] = 29'b0_011011110110_101_1_000110111101;
      patterns[14262] = 29'b0_011011110110_110_0_011011110110;
      patterns[14263] = 29'b0_011011110110_111_0_011011110110;
      patterns[14264] = 29'b0_011011110111_000_0_011011110111;
      patterns[14265] = 29'b0_011011110111_001_0_110111011011;
      patterns[14266] = 29'b0_011011110111_010_0_110111101110;
      patterns[14267] = 29'b0_011011110111_011_1_101111011100;
      patterns[14268] = 29'b0_011011110111_100_1_001101111011;
      patterns[14269] = 29'b0_011011110111_101_1_100110111101;
      patterns[14270] = 29'b0_011011110111_110_0_011011110111;
      patterns[14271] = 29'b0_011011110111_111_0_011011110111;
      patterns[14272] = 29'b0_011011111000_000_0_011011111000;
      patterns[14273] = 29'b0_011011111000_001_0_111000011011;
      patterns[14274] = 29'b0_011011111000_010_0_110111110000;
      patterns[14275] = 29'b0_011011111000_011_1_101111100000;
      patterns[14276] = 29'b0_011011111000_100_0_001101111100;
      patterns[14277] = 29'b0_011011111000_101_0_000110111110;
      patterns[14278] = 29'b0_011011111000_110_0_011011111000;
      patterns[14279] = 29'b0_011011111000_111_0_011011111000;
      patterns[14280] = 29'b0_011011111001_000_0_011011111001;
      patterns[14281] = 29'b0_011011111001_001_0_111001011011;
      patterns[14282] = 29'b0_011011111001_010_0_110111110010;
      patterns[14283] = 29'b0_011011111001_011_1_101111100100;
      patterns[14284] = 29'b0_011011111001_100_1_001101111100;
      patterns[14285] = 29'b0_011011111001_101_0_100110111110;
      patterns[14286] = 29'b0_011011111001_110_0_011011111001;
      patterns[14287] = 29'b0_011011111001_111_0_011011111001;
      patterns[14288] = 29'b0_011011111010_000_0_011011111010;
      patterns[14289] = 29'b0_011011111010_001_0_111010011011;
      patterns[14290] = 29'b0_011011111010_010_0_110111110100;
      patterns[14291] = 29'b0_011011111010_011_1_101111101000;
      patterns[14292] = 29'b0_011011111010_100_0_001101111101;
      patterns[14293] = 29'b0_011011111010_101_1_000110111110;
      patterns[14294] = 29'b0_011011111010_110_0_011011111010;
      patterns[14295] = 29'b0_011011111010_111_0_011011111010;
      patterns[14296] = 29'b0_011011111011_000_0_011011111011;
      patterns[14297] = 29'b0_011011111011_001_0_111011011011;
      patterns[14298] = 29'b0_011011111011_010_0_110111110110;
      patterns[14299] = 29'b0_011011111011_011_1_101111101100;
      patterns[14300] = 29'b0_011011111011_100_1_001101111101;
      patterns[14301] = 29'b0_011011111011_101_1_100110111110;
      patterns[14302] = 29'b0_011011111011_110_0_011011111011;
      patterns[14303] = 29'b0_011011111011_111_0_011011111011;
      patterns[14304] = 29'b0_011011111100_000_0_011011111100;
      patterns[14305] = 29'b0_011011111100_001_0_111100011011;
      patterns[14306] = 29'b0_011011111100_010_0_110111111000;
      patterns[14307] = 29'b0_011011111100_011_1_101111110000;
      patterns[14308] = 29'b0_011011111100_100_0_001101111110;
      patterns[14309] = 29'b0_011011111100_101_0_000110111111;
      patterns[14310] = 29'b0_011011111100_110_0_011011111100;
      patterns[14311] = 29'b0_011011111100_111_0_011011111100;
      patterns[14312] = 29'b0_011011111101_000_0_011011111101;
      patterns[14313] = 29'b0_011011111101_001_0_111101011011;
      patterns[14314] = 29'b0_011011111101_010_0_110111111010;
      patterns[14315] = 29'b0_011011111101_011_1_101111110100;
      patterns[14316] = 29'b0_011011111101_100_1_001101111110;
      patterns[14317] = 29'b0_011011111101_101_0_100110111111;
      patterns[14318] = 29'b0_011011111101_110_0_011011111101;
      patterns[14319] = 29'b0_011011111101_111_0_011011111101;
      patterns[14320] = 29'b0_011011111110_000_0_011011111110;
      patterns[14321] = 29'b0_011011111110_001_0_111110011011;
      patterns[14322] = 29'b0_011011111110_010_0_110111111100;
      patterns[14323] = 29'b0_011011111110_011_1_101111111000;
      patterns[14324] = 29'b0_011011111110_100_0_001101111111;
      patterns[14325] = 29'b0_011011111110_101_1_000110111111;
      patterns[14326] = 29'b0_011011111110_110_0_011011111110;
      patterns[14327] = 29'b0_011011111110_111_0_011011111110;
      patterns[14328] = 29'b0_011011111111_000_0_011011111111;
      patterns[14329] = 29'b0_011011111111_001_0_111111011011;
      patterns[14330] = 29'b0_011011111111_010_0_110111111110;
      patterns[14331] = 29'b0_011011111111_011_1_101111111100;
      patterns[14332] = 29'b0_011011111111_100_1_001101111111;
      patterns[14333] = 29'b0_011011111111_101_1_100110111111;
      patterns[14334] = 29'b0_011011111111_110_0_011011111111;
      patterns[14335] = 29'b0_011011111111_111_0_011011111111;
      patterns[14336] = 29'b0_011100000000_000_0_011100000000;
      patterns[14337] = 29'b0_011100000000_001_0_000000011100;
      patterns[14338] = 29'b0_011100000000_010_0_111000000000;
      patterns[14339] = 29'b0_011100000000_011_1_110000000000;
      patterns[14340] = 29'b0_011100000000_100_0_001110000000;
      patterns[14341] = 29'b0_011100000000_101_0_000111000000;
      patterns[14342] = 29'b0_011100000000_110_0_011100000000;
      patterns[14343] = 29'b0_011100000000_111_0_011100000000;
      patterns[14344] = 29'b0_011100000001_000_0_011100000001;
      patterns[14345] = 29'b0_011100000001_001_0_000001011100;
      patterns[14346] = 29'b0_011100000001_010_0_111000000010;
      patterns[14347] = 29'b0_011100000001_011_1_110000000100;
      patterns[14348] = 29'b0_011100000001_100_1_001110000000;
      patterns[14349] = 29'b0_011100000001_101_0_100111000000;
      patterns[14350] = 29'b0_011100000001_110_0_011100000001;
      patterns[14351] = 29'b0_011100000001_111_0_011100000001;
      patterns[14352] = 29'b0_011100000010_000_0_011100000010;
      patterns[14353] = 29'b0_011100000010_001_0_000010011100;
      patterns[14354] = 29'b0_011100000010_010_0_111000000100;
      patterns[14355] = 29'b0_011100000010_011_1_110000001000;
      patterns[14356] = 29'b0_011100000010_100_0_001110000001;
      patterns[14357] = 29'b0_011100000010_101_1_000111000000;
      patterns[14358] = 29'b0_011100000010_110_0_011100000010;
      patterns[14359] = 29'b0_011100000010_111_0_011100000010;
      patterns[14360] = 29'b0_011100000011_000_0_011100000011;
      patterns[14361] = 29'b0_011100000011_001_0_000011011100;
      patterns[14362] = 29'b0_011100000011_010_0_111000000110;
      patterns[14363] = 29'b0_011100000011_011_1_110000001100;
      patterns[14364] = 29'b0_011100000011_100_1_001110000001;
      patterns[14365] = 29'b0_011100000011_101_1_100111000000;
      patterns[14366] = 29'b0_011100000011_110_0_011100000011;
      patterns[14367] = 29'b0_011100000011_111_0_011100000011;
      patterns[14368] = 29'b0_011100000100_000_0_011100000100;
      patterns[14369] = 29'b0_011100000100_001_0_000100011100;
      patterns[14370] = 29'b0_011100000100_010_0_111000001000;
      patterns[14371] = 29'b0_011100000100_011_1_110000010000;
      patterns[14372] = 29'b0_011100000100_100_0_001110000010;
      patterns[14373] = 29'b0_011100000100_101_0_000111000001;
      patterns[14374] = 29'b0_011100000100_110_0_011100000100;
      patterns[14375] = 29'b0_011100000100_111_0_011100000100;
      patterns[14376] = 29'b0_011100000101_000_0_011100000101;
      patterns[14377] = 29'b0_011100000101_001_0_000101011100;
      patterns[14378] = 29'b0_011100000101_010_0_111000001010;
      patterns[14379] = 29'b0_011100000101_011_1_110000010100;
      patterns[14380] = 29'b0_011100000101_100_1_001110000010;
      patterns[14381] = 29'b0_011100000101_101_0_100111000001;
      patterns[14382] = 29'b0_011100000101_110_0_011100000101;
      patterns[14383] = 29'b0_011100000101_111_0_011100000101;
      patterns[14384] = 29'b0_011100000110_000_0_011100000110;
      patterns[14385] = 29'b0_011100000110_001_0_000110011100;
      patterns[14386] = 29'b0_011100000110_010_0_111000001100;
      patterns[14387] = 29'b0_011100000110_011_1_110000011000;
      patterns[14388] = 29'b0_011100000110_100_0_001110000011;
      patterns[14389] = 29'b0_011100000110_101_1_000111000001;
      patterns[14390] = 29'b0_011100000110_110_0_011100000110;
      patterns[14391] = 29'b0_011100000110_111_0_011100000110;
      patterns[14392] = 29'b0_011100000111_000_0_011100000111;
      patterns[14393] = 29'b0_011100000111_001_0_000111011100;
      patterns[14394] = 29'b0_011100000111_010_0_111000001110;
      patterns[14395] = 29'b0_011100000111_011_1_110000011100;
      patterns[14396] = 29'b0_011100000111_100_1_001110000011;
      patterns[14397] = 29'b0_011100000111_101_1_100111000001;
      patterns[14398] = 29'b0_011100000111_110_0_011100000111;
      patterns[14399] = 29'b0_011100000111_111_0_011100000111;
      patterns[14400] = 29'b0_011100001000_000_0_011100001000;
      patterns[14401] = 29'b0_011100001000_001_0_001000011100;
      patterns[14402] = 29'b0_011100001000_010_0_111000010000;
      patterns[14403] = 29'b0_011100001000_011_1_110000100000;
      patterns[14404] = 29'b0_011100001000_100_0_001110000100;
      patterns[14405] = 29'b0_011100001000_101_0_000111000010;
      patterns[14406] = 29'b0_011100001000_110_0_011100001000;
      patterns[14407] = 29'b0_011100001000_111_0_011100001000;
      patterns[14408] = 29'b0_011100001001_000_0_011100001001;
      patterns[14409] = 29'b0_011100001001_001_0_001001011100;
      patterns[14410] = 29'b0_011100001001_010_0_111000010010;
      patterns[14411] = 29'b0_011100001001_011_1_110000100100;
      patterns[14412] = 29'b0_011100001001_100_1_001110000100;
      patterns[14413] = 29'b0_011100001001_101_0_100111000010;
      patterns[14414] = 29'b0_011100001001_110_0_011100001001;
      patterns[14415] = 29'b0_011100001001_111_0_011100001001;
      patterns[14416] = 29'b0_011100001010_000_0_011100001010;
      patterns[14417] = 29'b0_011100001010_001_0_001010011100;
      patterns[14418] = 29'b0_011100001010_010_0_111000010100;
      patterns[14419] = 29'b0_011100001010_011_1_110000101000;
      patterns[14420] = 29'b0_011100001010_100_0_001110000101;
      patterns[14421] = 29'b0_011100001010_101_1_000111000010;
      patterns[14422] = 29'b0_011100001010_110_0_011100001010;
      patterns[14423] = 29'b0_011100001010_111_0_011100001010;
      patterns[14424] = 29'b0_011100001011_000_0_011100001011;
      patterns[14425] = 29'b0_011100001011_001_0_001011011100;
      patterns[14426] = 29'b0_011100001011_010_0_111000010110;
      patterns[14427] = 29'b0_011100001011_011_1_110000101100;
      patterns[14428] = 29'b0_011100001011_100_1_001110000101;
      patterns[14429] = 29'b0_011100001011_101_1_100111000010;
      patterns[14430] = 29'b0_011100001011_110_0_011100001011;
      patterns[14431] = 29'b0_011100001011_111_0_011100001011;
      patterns[14432] = 29'b0_011100001100_000_0_011100001100;
      patterns[14433] = 29'b0_011100001100_001_0_001100011100;
      patterns[14434] = 29'b0_011100001100_010_0_111000011000;
      patterns[14435] = 29'b0_011100001100_011_1_110000110000;
      patterns[14436] = 29'b0_011100001100_100_0_001110000110;
      patterns[14437] = 29'b0_011100001100_101_0_000111000011;
      patterns[14438] = 29'b0_011100001100_110_0_011100001100;
      patterns[14439] = 29'b0_011100001100_111_0_011100001100;
      patterns[14440] = 29'b0_011100001101_000_0_011100001101;
      patterns[14441] = 29'b0_011100001101_001_0_001101011100;
      patterns[14442] = 29'b0_011100001101_010_0_111000011010;
      patterns[14443] = 29'b0_011100001101_011_1_110000110100;
      patterns[14444] = 29'b0_011100001101_100_1_001110000110;
      patterns[14445] = 29'b0_011100001101_101_0_100111000011;
      patterns[14446] = 29'b0_011100001101_110_0_011100001101;
      patterns[14447] = 29'b0_011100001101_111_0_011100001101;
      patterns[14448] = 29'b0_011100001110_000_0_011100001110;
      patterns[14449] = 29'b0_011100001110_001_0_001110011100;
      patterns[14450] = 29'b0_011100001110_010_0_111000011100;
      patterns[14451] = 29'b0_011100001110_011_1_110000111000;
      patterns[14452] = 29'b0_011100001110_100_0_001110000111;
      patterns[14453] = 29'b0_011100001110_101_1_000111000011;
      patterns[14454] = 29'b0_011100001110_110_0_011100001110;
      patterns[14455] = 29'b0_011100001110_111_0_011100001110;
      patterns[14456] = 29'b0_011100001111_000_0_011100001111;
      patterns[14457] = 29'b0_011100001111_001_0_001111011100;
      patterns[14458] = 29'b0_011100001111_010_0_111000011110;
      patterns[14459] = 29'b0_011100001111_011_1_110000111100;
      patterns[14460] = 29'b0_011100001111_100_1_001110000111;
      patterns[14461] = 29'b0_011100001111_101_1_100111000011;
      patterns[14462] = 29'b0_011100001111_110_0_011100001111;
      patterns[14463] = 29'b0_011100001111_111_0_011100001111;
      patterns[14464] = 29'b0_011100010000_000_0_011100010000;
      patterns[14465] = 29'b0_011100010000_001_0_010000011100;
      patterns[14466] = 29'b0_011100010000_010_0_111000100000;
      patterns[14467] = 29'b0_011100010000_011_1_110001000000;
      patterns[14468] = 29'b0_011100010000_100_0_001110001000;
      patterns[14469] = 29'b0_011100010000_101_0_000111000100;
      patterns[14470] = 29'b0_011100010000_110_0_011100010000;
      patterns[14471] = 29'b0_011100010000_111_0_011100010000;
      patterns[14472] = 29'b0_011100010001_000_0_011100010001;
      patterns[14473] = 29'b0_011100010001_001_0_010001011100;
      patterns[14474] = 29'b0_011100010001_010_0_111000100010;
      patterns[14475] = 29'b0_011100010001_011_1_110001000100;
      patterns[14476] = 29'b0_011100010001_100_1_001110001000;
      patterns[14477] = 29'b0_011100010001_101_0_100111000100;
      patterns[14478] = 29'b0_011100010001_110_0_011100010001;
      patterns[14479] = 29'b0_011100010001_111_0_011100010001;
      patterns[14480] = 29'b0_011100010010_000_0_011100010010;
      patterns[14481] = 29'b0_011100010010_001_0_010010011100;
      patterns[14482] = 29'b0_011100010010_010_0_111000100100;
      patterns[14483] = 29'b0_011100010010_011_1_110001001000;
      patterns[14484] = 29'b0_011100010010_100_0_001110001001;
      patterns[14485] = 29'b0_011100010010_101_1_000111000100;
      patterns[14486] = 29'b0_011100010010_110_0_011100010010;
      patterns[14487] = 29'b0_011100010010_111_0_011100010010;
      patterns[14488] = 29'b0_011100010011_000_0_011100010011;
      patterns[14489] = 29'b0_011100010011_001_0_010011011100;
      patterns[14490] = 29'b0_011100010011_010_0_111000100110;
      patterns[14491] = 29'b0_011100010011_011_1_110001001100;
      patterns[14492] = 29'b0_011100010011_100_1_001110001001;
      patterns[14493] = 29'b0_011100010011_101_1_100111000100;
      patterns[14494] = 29'b0_011100010011_110_0_011100010011;
      patterns[14495] = 29'b0_011100010011_111_0_011100010011;
      patterns[14496] = 29'b0_011100010100_000_0_011100010100;
      patterns[14497] = 29'b0_011100010100_001_0_010100011100;
      patterns[14498] = 29'b0_011100010100_010_0_111000101000;
      patterns[14499] = 29'b0_011100010100_011_1_110001010000;
      patterns[14500] = 29'b0_011100010100_100_0_001110001010;
      patterns[14501] = 29'b0_011100010100_101_0_000111000101;
      patterns[14502] = 29'b0_011100010100_110_0_011100010100;
      patterns[14503] = 29'b0_011100010100_111_0_011100010100;
      patterns[14504] = 29'b0_011100010101_000_0_011100010101;
      patterns[14505] = 29'b0_011100010101_001_0_010101011100;
      patterns[14506] = 29'b0_011100010101_010_0_111000101010;
      patterns[14507] = 29'b0_011100010101_011_1_110001010100;
      patterns[14508] = 29'b0_011100010101_100_1_001110001010;
      patterns[14509] = 29'b0_011100010101_101_0_100111000101;
      patterns[14510] = 29'b0_011100010101_110_0_011100010101;
      patterns[14511] = 29'b0_011100010101_111_0_011100010101;
      patterns[14512] = 29'b0_011100010110_000_0_011100010110;
      patterns[14513] = 29'b0_011100010110_001_0_010110011100;
      patterns[14514] = 29'b0_011100010110_010_0_111000101100;
      patterns[14515] = 29'b0_011100010110_011_1_110001011000;
      patterns[14516] = 29'b0_011100010110_100_0_001110001011;
      patterns[14517] = 29'b0_011100010110_101_1_000111000101;
      patterns[14518] = 29'b0_011100010110_110_0_011100010110;
      patterns[14519] = 29'b0_011100010110_111_0_011100010110;
      patterns[14520] = 29'b0_011100010111_000_0_011100010111;
      patterns[14521] = 29'b0_011100010111_001_0_010111011100;
      patterns[14522] = 29'b0_011100010111_010_0_111000101110;
      patterns[14523] = 29'b0_011100010111_011_1_110001011100;
      patterns[14524] = 29'b0_011100010111_100_1_001110001011;
      patterns[14525] = 29'b0_011100010111_101_1_100111000101;
      patterns[14526] = 29'b0_011100010111_110_0_011100010111;
      patterns[14527] = 29'b0_011100010111_111_0_011100010111;
      patterns[14528] = 29'b0_011100011000_000_0_011100011000;
      patterns[14529] = 29'b0_011100011000_001_0_011000011100;
      patterns[14530] = 29'b0_011100011000_010_0_111000110000;
      patterns[14531] = 29'b0_011100011000_011_1_110001100000;
      patterns[14532] = 29'b0_011100011000_100_0_001110001100;
      patterns[14533] = 29'b0_011100011000_101_0_000111000110;
      patterns[14534] = 29'b0_011100011000_110_0_011100011000;
      patterns[14535] = 29'b0_011100011000_111_0_011100011000;
      patterns[14536] = 29'b0_011100011001_000_0_011100011001;
      patterns[14537] = 29'b0_011100011001_001_0_011001011100;
      patterns[14538] = 29'b0_011100011001_010_0_111000110010;
      patterns[14539] = 29'b0_011100011001_011_1_110001100100;
      patterns[14540] = 29'b0_011100011001_100_1_001110001100;
      patterns[14541] = 29'b0_011100011001_101_0_100111000110;
      patterns[14542] = 29'b0_011100011001_110_0_011100011001;
      patterns[14543] = 29'b0_011100011001_111_0_011100011001;
      patterns[14544] = 29'b0_011100011010_000_0_011100011010;
      patterns[14545] = 29'b0_011100011010_001_0_011010011100;
      patterns[14546] = 29'b0_011100011010_010_0_111000110100;
      patterns[14547] = 29'b0_011100011010_011_1_110001101000;
      patterns[14548] = 29'b0_011100011010_100_0_001110001101;
      patterns[14549] = 29'b0_011100011010_101_1_000111000110;
      patterns[14550] = 29'b0_011100011010_110_0_011100011010;
      patterns[14551] = 29'b0_011100011010_111_0_011100011010;
      patterns[14552] = 29'b0_011100011011_000_0_011100011011;
      patterns[14553] = 29'b0_011100011011_001_0_011011011100;
      patterns[14554] = 29'b0_011100011011_010_0_111000110110;
      patterns[14555] = 29'b0_011100011011_011_1_110001101100;
      patterns[14556] = 29'b0_011100011011_100_1_001110001101;
      patterns[14557] = 29'b0_011100011011_101_1_100111000110;
      patterns[14558] = 29'b0_011100011011_110_0_011100011011;
      patterns[14559] = 29'b0_011100011011_111_0_011100011011;
      patterns[14560] = 29'b0_011100011100_000_0_011100011100;
      patterns[14561] = 29'b0_011100011100_001_0_011100011100;
      patterns[14562] = 29'b0_011100011100_010_0_111000111000;
      patterns[14563] = 29'b0_011100011100_011_1_110001110000;
      patterns[14564] = 29'b0_011100011100_100_0_001110001110;
      patterns[14565] = 29'b0_011100011100_101_0_000111000111;
      patterns[14566] = 29'b0_011100011100_110_0_011100011100;
      patterns[14567] = 29'b0_011100011100_111_0_011100011100;
      patterns[14568] = 29'b0_011100011101_000_0_011100011101;
      patterns[14569] = 29'b0_011100011101_001_0_011101011100;
      patterns[14570] = 29'b0_011100011101_010_0_111000111010;
      patterns[14571] = 29'b0_011100011101_011_1_110001110100;
      patterns[14572] = 29'b0_011100011101_100_1_001110001110;
      patterns[14573] = 29'b0_011100011101_101_0_100111000111;
      patterns[14574] = 29'b0_011100011101_110_0_011100011101;
      patterns[14575] = 29'b0_011100011101_111_0_011100011101;
      patterns[14576] = 29'b0_011100011110_000_0_011100011110;
      patterns[14577] = 29'b0_011100011110_001_0_011110011100;
      patterns[14578] = 29'b0_011100011110_010_0_111000111100;
      patterns[14579] = 29'b0_011100011110_011_1_110001111000;
      patterns[14580] = 29'b0_011100011110_100_0_001110001111;
      patterns[14581] = 29'b0_011100011110_101_1_000111000111;
      patterns[14582] = 29'b0_011100011110_110_0_011100011110;
      patterns[14583] = 29'b0_011100011110_111_0_011100011110;
      patterns[14584] = 29'b0_011100011111_000_0_011100011111;
      patterns[14585] = 29'b0_011100011111_001_0_011111011100;
      patterns[14586] = 29'b0_011100011111_010_0_111000111110;
      patterns[14587] = 29'b0_011100011111_011_1_110001111100;
      patterns[14588] = 29'b0_011100011111_100_1_001110001111;
      patterns[14589] = 29'b0_011100011111_101_1_100111000111;
      patterns[14590] = 29'b0_011100011111_110_0_011100011111;
      patterns[14591] = 29'b0_011100011111_111_0_011100011111;
      patterns[14592] = 29'b0_011100100000_000_0_011100100000;
      patterns[14593] = 29'b0_011100100000_001_0_100000011100;
      patterns[14594] = 29'b0_011100100000_010_0_111001000000;
      patterns[14595] = 29'b0_011100100000_011_1_110010000000;
      patterns[14596] = 29'b0_011100100000_100_0_001110010000;
      patterns[14597] = 29'b0_011100100000_101_0_000111001000;
      patterns[14598] = 29'b0_011100100000_110_0_011100100000;
      patterns[14599] = 29'b0_011100100000_111_0_011100100000;
      patterns[14600] = 29'b0_011100100001_000_0_011100100001;
      patterns[14601] = 29'b0_011100100001_001_0_100001011100;
      patterns[14602] = 29'b0_011100100001_010_0_111001000010;
      patterns[14603] = 29'b0_011100100001_011_1_110010000100;
      patterns[14604] = 29'b0_011100100001_100_1_001110010000;
      patterns[14605] = 29'b0_011100100001_101_0_100111001000;
      patterns[14606] = 29'b0_011100100001_110_0_011100100001;
      patterns[14607] = 29'b0_011100100001_111_0_011100100001;
      patterns[14608] = 29'b0_011100100010_000_0_011100100010;
      patterns[14609] = 29'b0_011100100010_001_0_100010011100;
      patterns[14610] = 29'b0_011100100010_010_0_111001000100;
      patterns[14611] = 29'b0_011100100010_011_1_110010001000;
      patterns[14612] = 29'b0_011100100010_100_0_001110010001;
      patterns[14613] = 29'b0_011100100010_101_1_000111001000;
      patterns[14614] = 29'b0_011100100010_110_0_011100100010;
      patterns[14615] = 29'b0_011100100010_111_0_011100100010;
      patterns[14616] = 29'b0_011100100011_000_0_011100100011;
      patterns[14617] = 29'b0_011100100011_001_0_100011011100;
      patterns[14618] = 29'b0_011100100011_010_0_111001000110;
      patterns[14619] = 29'b0_011100100011_011_1_110010001100;
      patterns[14620] = 29'b0_011100100011_100_1_001110010001;
      patterns[14621] = 29'b0_011100100011_101_1_100111001000;
      patterns[14622] = 29'b0_011100100011_110_0_011100100011;
      patterns[14623] = 29'b0_011100100011_111_0_011100100011;
      patterns[14624] = 29'b0_011100100100_000_0_011100100100;
      patterns[14625] = 29'b0_011100100100_001_0_100100011100;
      patterns[14626] = 29'b0_011100100100_010_0_111001001000;
      patterns[14627] = 29'b0_011100100100_011_1_110010010000;
      patterns[14628] = 29'b0_011100100100_100_0_001110010010;
      patterns[14629] = 29'b0_011100100100_101_0_000111001001;
      patterns[14630] = 29'b0_011100100100_110_0_011100100100;
      patterns[14631] = 29'b0_011100100100_111_0_011100100100;
      patterns[14632] = 29'b0_011100100101_000_0_011100100101;
      patterns[14633] = 29'b0_011100100101_001_0_100101011100;
      patterns[14634] = 29'b0_011100100101_010_0_111001001010;
      patterns[14635] = 29'b0_011100100101_011_1_110010010100;
      patterns[14636] = 29'b0_011100100101_100_1_001110010010;
      patterns[14637] = 29'b0_011100100101_101_0_100111001001;
      patterns[14638] = 29'b0_011100100101_110_0_011100100101;
      patterns[14639] = 29'b0_011100100101_111_0_011100100101;
      patterns[14640] = 29'b0_011100100110_000_0_011100100110;
      patterns[14641] = 29'b0_011100100110_001_0_100110011100;
      patterns[14642] = 29'b0_011100100110_010_0_111001001100;
      patterns[14643] = 29'b0_011100100110_011_1_110010011000;
      patterns[14644] = 29'b0_011100100110_100_0_001110010011;
      patterns[14645] = 29'b0_011100100110_101_1_000111001001;
      patterns[14646] = 29'b0_011100100110_110_0_011100100110;
      patterns[14647] = 29'b0_011100100110_111_0_011100100110;
      patterns[14648] = 29'b0_011100100111_000_0_011100100111;
      patterns[14649] = 29'b0_011100100111_001_0_100111011100;
      patterns[14650] = 29'b0_011100100111_010_0_111001001110;
      patterns[14651] = 29'b0_011100100111_011_1_110010011100;
      patterns[14652] = 29'b0_011100100111_100_1_001110010011;
      patterns[14653] = 29'b0_011100100111_101_1_100111001001;
      patterns[14654] = 29'b0_011100100111_110_0_011100100111;
      patterns[14655] = 29'b0_011100100111_111_0_011100100111;
      patterns[14656] = 29'b0_011100101000_000_0_011100101000;
      patterns[14657] = 29'b0_011100101000_001_0_101000011100;
      patterns[14658] = 29'b0_011100101000_010_0_111001010000;
      patterns[14659] = 29'b0_011100101000_011_1_110010100000;
      patterns[14660] = 29'b0_011100101000_100_0_001110010100;
      patterns[14661] = 29'b0_011100101000_101_0_000111001010;
      patterns[14662] = 29'b0_011100101000_110_0_011100101000;
      patterns[14663] = 29'b0_011100101000_111_0_011100101000;
      patterns[14664] = 29'b0_011100101001_000_0_011100101001;
      patterns[14665] = 29'b0_011100101001_001_0_101001011100;
      patterns[14666] = 29'b0_011100101001_010_0_111001010010;
      patterns[14667] = 29'b0_011100101001_011_1_110010100100;
      patterns[14668] = 29'b0_011100101001_100_1_001110010100;
      patterns[14669] = 29'b0_011100101001_101_0_100111001010;
      patterns[14670] = 29'b0_011100101001_110_0_011100101001;
      patterns[14671] = 29'b0_011100101001_111_0_011100101001;
      patterns[14672] = 29'b0_011100101010_000_0_011100101010;
      patterns[14673] = 29'b0_011100101010_001_0_101010011100;
      patterns[14674] = 29'b0_011100101010_010_0_111001010100;
      patterns[14675] = 29'b0_011100101010_011_1_110010101000;
      patterns[14676] = 29'b0_011100101010_100_0_001110010101;
      patterns[14677] = 29'b0_011100101010_101_1_000111001010;
      patterns[14678] = 29'b0_011100101010_110_0_011100101010;
      patterns[14679] = 29'b0_011100101010_111_0_011100101010;
      patterns[14680] = 29'b0_011100101011_000_0_011100101011;
      patterns[14681] = 29'b0_011100101011_001_0_101011011100;
      patterns[14682] = 29'b0_011100101011_010_0_111001010110;
      patterns[14683] = 29'b0_011100101011_011_1_110010101100;
      patterns[14684] = 29'b0_011100101011_100_1_001110010101;
      patterns[14685] = 29'b0_011100101011_101_1_100111001010;
      patterns[14686] = 29'b0_011100101011_110_0_011100101011;
      patterns[14687] = 29'b0_011100101011_111_0_011100101011;
      patterns[14688] = 29'b0_011100101100_000_0_011100101100;
      patterns[14689] = 29'b0_011100101100_001_0_101100011100;
      patterns[14690] = 29'b0_011100101100_010_0_111001011000;
      patterns[14691] = 29'b0_011100101100_011_1_110010110000;
      patterns[14692] = 29'b0_011100101100_100_0_001110010110;
      patterns[14693] = 29'b0_011100101100_101_0_000111001011;
      patterns[14694] = 29'b0_011100101100_110_0_011100101100;
      patterns[14695] = 29'b0_011100101100_111_0_011100101100;
      patterns[14696] = 29'b0_011100101101_000_0_011100101101;
      patterns[14697] = 29'b0_011100101101_001_0_101101011100;
      patterns[14698] = 29'b0_011100101101_010_0_111001011010;
      patterns[14699] = 29'b0_011100101101_011_1_110010110100;
      patterns[14700] = 29'b0_011100101101_100_1_001110010110;
      patterns[14701] = 29'b0_011100101101_101_0_100111001011;
      patterns[14702] = 29'b0_011100101101_110_0_011100101101;
      patterns[14703] = 29'b0_011100101101_111_0_011100101101;
      patterns[14704] = 29'b0_011100101110_000_0_011100101110;
      patterns[14705] = 29'b0_011100101110_001_0_101110011100;
      patterns[14706] = 29'b0_011100101110_010_0_111001011100;
      patterns[14707] = 29'b0_011100101110_011_1_110010111000;
      patterns[14708] = 29'b0_011100101110_100_0_001110010111;
      patterns[14709] = 29'b0_011100101110_101_1_000111001011;
      patterns[14710] = 29'b0_011100101110_110_0_011100101110;
      patterns[14711] = 29'b0_011100101110_111_0_011100101110;
      patterns[14712] = 29'b0_011100101111_000_0_011100101111;
      patterns[14713] = 29'b0_011100101111_001_0_101111011100;
      patterns[14714] = 29'b0_011100101111_010_0_111001011110;
      patterns[14715] = 29'b0_011100101111_011_1_110010111100;
      patterns[14716] = 29'b0_011100101111_100_1_001110010111;
      patterns[14717] = 29'b0_011100101111_101_1_100111001011;
      patterns[14718] = 29'b0_011100101111_110_0_011100101111;
      patterns[14719] = 29'b0_011100101111_111_0_011100101111;
      patterns[14720] = 29'b0_011100110000_000_0_011100110000;
      patterns[14721] = 29'b0_011100110000_001_0_110000011100;
      patterns[14722] = 29'b0_011100110000_010_0_111001100000;
      patterns[14723] = 29'b0_011100110000_011_1_110011000000;
      patterns[14724] = 29'b0_011100110000_100_0_001110011000;
      patterns[14725] = 29'b0_011100110000_101_0_000111001100;
      patterns[14726] = 29'b0_011100110000_110_0_011100110000;
      patterns[14727] = 29'b0_011100110000_111_0_011100110000;
      patterns[14728] = 29'b0_011100110001_000_0_011100110001;
      patterns[14729] = 29'b0_011100110001_001_0_110001011100;
      patterns[14730] = 29'b0_011100110001_010_0_111001100010;
      patterns[14731] = 29'b0_011100110001_011_1_110011000100;
      patterns[14732] = 29'b0_011100110001_100_1_001110011000;
      patterns[14733] = 29'b0_011100110001_101_0_100111001100;
      patterns[14734] = 29'b0_011100110001_110_0_011100110001;
      patterns[14735] = 29'b0_011100110001_111_0_011100110001;
      patterns[14736] = 29'b0_011100110010_000_0_011100110010;
      patterns[14737] = 29'b0_011100110010_001_0_110010011100;
      patterns[14738] = 29'b0_011100110010_010_0_111001100100;
      patterns[14739] = 29'b0_011100110010_011_1_110011001000;
      patterns[14740] = 29'b0_011100110010_100_0_001110011001;
      patterns[14741] = 29'b0_011100110010_101_1_000111001100;
      patterns[14742] = 29'b0_011100110010_110_0_011100110010;
      patterns[14743] = 29'b0_011100110010_111_0_011100110010;
      patterns[14744] = 29'b0_011100110011_000_0_011100110011;
      patterns[14745] = 29'b0_011100110011_001_0_110011011100;
      patterns[14746] = 29'b0_011100110011_010_0_111001100110;
      patterns[14747] = 29'b0_011100110011_011_1_110011001100;
      patterns[14748] = 29'b0_011100110011_100_1_001110011001;
      patterns[14749] = 29'b0_011100110011_101_1_100111001100;
      patterns[14750] = 29'b0_011100110011_110_0_011100110011;
      patterns[14751] = 29'b0_011100110011_111_0_011100110011;
      patterns[14752] = 29'b0_011100110100_000_0_011100110100;
      patterns[14753] = 29'b0_011100110100_001_0_110100011100;
      patterns[14754] = 29'b0_011100110100_010_0_111001101000;
      patterns[14755] = 29'b0_011100110100_011_1_110011010000;
      patterns[14756] = 29'b0_011100110100_100_0_001110011010;
      patterns[14757] = 29'b0_011100110100_101_0_000111001101;
      patterns[14758] = 29'b0_011100110100_110_0_011100110100;
      patterns[14759] = 29'b0_011100110100_111_0_011100110100;
      patterns[14760] = 29'b0_011100110101_000_0_011100110101;
      patterns[14761] = 29'b0_011100110101_001_0_110101011100;
      patterns[14762] = 29'b0_011100110101_010_0_111001101010;
      patterns[14763] = 29'b0_011100110101_011_1_110011010100;
      patterns[14764] = 29'b0_011100110101_100_1_001110011010;
      patterns[14765] = 29'b0_011100110101_101_0_100111001101;
      patterns[14766] = 29'b0_011100110101_110_0_011100110101;
      patterns[14767] = 29'b0_011100110101_111_0_011100110101;
      patterns[14768] = 29'b0_011100110110_000_0_011100110110;
      patterns[14769] = 29'b0_011100110110_001_0_110110011100;
      patterns[14770] = 29'b0_011100110110_010_0_111001101100;
      patterns[14771] = 29'b0_011100110110_011_1_110011011000;
      patterns[14772] = 29'b0_011100110110_100_0_001110011011;
      patterns[14773] = 29'b0_011100110110_101_1_000111001101;
      patterns[14774] = 29'b0_011100110110_110_0_011100110110;
      patterns[14775] = 29'b0_011100110110_111_0_011100110110;
      patterns[14776] = 29'b0_011100110111_000_0_011100110111;
      patterns[14777] = 29'b0_011100110111_001_0_110111011100;
      patterns[14778] = 29'b0_011100110111_010_0_111001101110;
      patterns[14779] = 29'b0_011100110111_011_1_110011011100;
      patterns[14780] = 29'b0_011100110111_100_1_001110011011;
      patterns[14781] = 29'b0_011100110111_101_1_100111001101;
      patterns[14782] = 29'b0_011100110111_110_0_011100110111;
      patterns[14783] = 29'b0_011100110111_111_0_011100110111;
      patterns[14784] = 29'b0_011100111000_000_0_011100111000;
      patterns[14785] = 29'b0_011100111000_001_0_111000011100;
      patterns[14786] = 29'b0_011100111000_010_0_111001110000;
      patterns[14787] = 29'b0_011100111000_011_1_110011100000;
      patterns[14788] = 29'b0_011100111000_100_0_001110011100;
      patterns[14789] = 29'b0_011100111000_101_0_000111001110;
      patterns[14790] = 29'b0_011100111000_110_0_011100111000;
      patterns[14791] = 29'b0_011100111000_111_0_011100111000;
      patterns[14792] = 29'b0_011100111001_000_0_011100111001;
      patterns[14793] = 29'b0_011100111001_001_0_111001011100;
      patterns[14794] = 29'b0_011100111001_010_0_111001110010;
      patterns[14795] = 29'b0_011100111001_011_1_110011100100;
      patterns[14796] = 29'b0_011100111001_100_1_001110011100;
      patterns[14797] = 29'b0_011100111001_101_0_100111001110;
      patterns[14798] = 29'b0_011100111001_110_0_011100111001;
      patterns[14799] = 29'b0_011100111001_111_0_011100111001;
      patterns[14800] = 29'b0_011100111010_000_0_011100111010;
      patterns[14801] = 29'b0_011100111010_001_0_111010011100;
      patterns[14802] = 29'b0_011100111010_010_0_111001110100;
      patterns[14803] = 29'b0_011100111010_011_1_110011101000;
      patterns[14804] = 29'b0_011100111010_100_0_001110011101;
      patterns[14805] = 29'b0_011100111010_101_1_000111001110;
      patterns[14806] = 29'b0_011100111010_110_0_011100111010;
      patterns[14807] = 29'b0_011100111010_111_0_011100111010;
      patterns[14808] = 29'b0_011100111011_000_0_011100111011;
      patterns[14809] = 29'b0_011100111011_001_0_111011011100;
      patterns[14810] = 29'b0_011100111011_010_0_111001110110;
      patterns[14811] = 29'b0_011100111011_011_1_110011101100;
      patterns[14812] = 29'b0_011100111011_100_1_001110011101;
      patterns[14813] = 29'b0_011100111011_101_1_100111001110;
      patterns[14814] = 29'b0_011100111011_110_0_011100111011;
      patterns[14815] = 29'b0_011100111011_111_0_011100111011;
      patterns[14816] = 29'b0_011100111100_000_0_011100111100;
      patterns[14817] = 29'b0_011100111100_001_0_111100011100;
      patterns[14818] = 29'b0_011100111100_010_0_111001111000;
      patterns[14819] = 29'b0_011100111100_011_1_110011110000;
      patterns[14820] = 29'b0_011100111100_100_0_001110011110;
      patterns[14821] = 29'b0_011100111100_101_0_000111001111;
      patterns[14822] = 29'b0_011100111100_110_0_011100111100;
      patterns[14823] = 29'b0_011100111100_111_0_011100111100;
      patterns[14824] = 29'b0_011100111101_000_0_011100111101;
      patterns[14825] = 29'b0_011100111101_001_0_111101011100;
      patterns[14826] = 29'b0_011100111101_010_0_111001111010;
      patterns[14827] = 29'b0_011100111101_011_1_110011110100;
      patterns[14828] = 29'b0_011100111101_100_1_001110011110;
      patterns[14829] = 29'b0_011100111101_101_0_100111001111;
      patterns[14830] = 29'b0_011100111101_110_0_011100111101;
      patterns[14831] = 29'b0_011100111101_111_0_011100111101;
      patterns[14832] = 29'b0_011100111110_000_0_011100111110;
      patterns[14833] = 29'b0_011100111110_001_0_111110011100;
      patterns[14834] = 29'b0_011100111110_010_0_111001111100;
      patterns[14835] = 29'b0_011100111110_011_1_110011111000;
      patterns[14836] = 29'b0_011100111110_100_0_001110011111;
      patterns[14837] = 29'b0_011100111110_101_1_000111001111;
      patterns[14838] = 29'b0_011100111110_110_0_011100111110;
      patterns[14839] = 29'b0_011100111110_111_0_011100111110;
      patterns[14840] = 29'b0_011100111111_000_0_011100111111;
      patterns[14841] = 29'b0_011100111111_001_0_111111011100;
      patterns[14842] = 29'b0_011100111111_010_0_111001111110;
      patterns[14843] = 29'b0_011100111111_011_1_110011111100;
      patterns[14844] = 29'b0_011100111111_100_1_001110011111;
      patterns[14845] = 29'b0_011100111111_101_1_100111001111;
      patterns[14846] = 29'b0_011100111111_110_0_011100111111;
      patterns[14847] = 29'b0_011100111111_111_0_011100111111;
      patterns[14848] = 29'b0_011101000000_000_0_011101000000;
      patterns[14849] = 29'b0_011101000000_001_0_000000011101;
      patterns[14850] = 29'b0_011101000000_010_0_111010000000;
      patterns[14851] = 29'b0_011101000000_011_1_110100000000;
      patterns[14852] = 29'b0_011101000000_100_0_001110100000;
      patterns[14853] = 29'b0_011101000000_101_0_000111010000;
      patterns[14854] = 29'b0_011101000000_110_0_011101000000;
      patterns[14855] = 29'b0_011101000000_111_0_011101000000;
      patterns[14856] = 29'b0_011101000001_000_0_011101000001;
      patterns[14857] = 29'b0_011101000001_001_0_000001011101;
      patterns[14858] = 29'b0_011101000001_010_0_111010000010;
      patterns[14859] = 29'b0_011101000001_011_1_110100000100;
      patterns[14860] = 29'b0_011101000001_100_1_001110100000;
      patterns[14861] = 29'b0_011101000001_101_0_100111010000;
      patterns[14862] = 29'b0_011101000001_110_0_011101000001;
      patterns[14863] = 29'b0_011101000001_111_0_011101000001;
      patterns[14864] = 29'b0_011101000010_000_0_011101000010;
      patterns[14865] = 29'b0_011101000010_001_0_000010011101;
      patterns[14866] = 29'b0_011101000010_010_0_111010000100;
      patterns[14867] = 29'b0_011101000010_011_1_110100001000;
      patterns[14868] = 29'b0_011101000010_100_0_001110100001;
      patterns[14869] = 29'b0_011101000010_101_1_000111010000;
      patterns[14870] = 29'b0_011101000010_110_0_011101000010;
      patterns[14871] = 29'b0_011101000010_111_0_011101000010;
      patterns[14872] = 29'b0_011101000011_000_0_011101000011;
      patterns[14873] = 29'b0_011101000011_001_0_000011011101;
      patterns[14874] = 29'b0_011101000011_010_0_111010000110;
      patterns[14875] = 29'b0_011101000011_011_1_110100001100;
      patterns[14876] = 29'b0_011101000011_100_1_001110100001;
      patterns[14877] = 29'b0_011101000011_101_1_100111010000;
      patterns[14878] = 29'b0_011101000011_110_0_011101000011;
      patterns[14879] = 29'b0_011101000011_111_0_011101000011;
      patterns[14880] = 29'b0_011101000100_000_0_011101000100;
      patterns[14881] = 29'b0_011101000100_001_0_000100011101;
      patterns[14882] = 29'b0_011101000100_010_0_111010001000;
      patterns[14883] = 29'b0_011101000100_011_1_110100010000;
      patterns[14884] = 29'b0_011101000100_100_0_001110100010;
      patterns[14885] = 29'b0_011101000100_101_0_000111010001;
      patterns[14886] = 29'b0_011101000100_110_0_011101000100;
      patterns[14887] = 29'b0_011101000100_111_0_011101000100;
      patterns[14888] = 29'b0_011101000101_000_0_011101000101;
      patterns[14889] = 29'b0_011101000101_001_0_000101011101;
      patterns[14890] = 29'b0_011101000101_010_0_111010001010;
      patterns[14891] = 29'b0_011101000101_011_1_110100010100;
      patterns[14892] = 29'b0_011101000101_100_1_001110100010;
      patterns[14893] = 29'b0_011101000101_101_0_100111010001;
      patterns[14894] = 29'b0_011101000101_110_0_011101000101;
      patterns[14895] = 29'b0_011101000101_111_0_011101000101;
      patterns[14896] = 29'b0_011101000110_000_0_011101000110;
      patterns[14897] = 29'b0_011101000110_001_0_000110011101;
      patterns[14898] = 29'b0_011101000110_010_0_111010001100;
      patterns[14899] = 29'b0_011101000110_011_1_110100011000;
      patterns[14900] = 29'b0_011101000110_100_0_001110100011;
      patterns[14901] = 29'b0_011101000110_101_1_000111010001;
      patterns[14902] = 29'b0_011101000110_110_0_011101000110;
      patterns[14903] = 29'b0_011101000110_111_0_011101000110;
      patterns[14904] = 29'b0_011101000111_000_0_011101000111;
      patterns[14905] = 29'b0_011101000111_001_0_000111011101;
      patterns[14906] = 29'b0_011101000111_010_0_111010001110;
      patterns[14907] = 29'b0_011101000111_011_1_110100011100;
      patterns[14908] = 29'b0_011101000111_100_1_001110100011;
      patterns[14909] = 29'b0_011101000111_101_1_100111010001;
      patterns[14910] = 29'b0_011101000111_110_0_011101000111;
      patterns[14911] = 29'b0_011101000111_111_0_011101000111;
      patterns[14912] = 29'b0_011101001000_000_0_011101001000;
      patterns[14913] = 29'b0_011101001000_001_0_001000011101;
      patterns[14914] = 29'b0_011101001000_010_0_111010010000;
      patterns[14915] = 29'b0_011101001000_011_1_110100100000;
      patterns[14916] = 29'b0_011101001000_100_0_001110100100;
      patterns[14917] = 29'b0_011101001000_101_0_000111010010;
      patterns[14918] = 29'b0_011101001000_110_0_011101001000;
      patterns[14919] = 29'b0_011101001000_111_0_011101001000;
      patterns[14920] = 29'b0_011101001001_000_0_011101001001;
      patterns[14921] = 29'b0_011101001001_001_0_001001011101;
      patterns[14922] = 29'b0_011101001001_010_0_111010010010;
      patterns[14923] = 29'b0_011101001001_011_1_110100100100;
      patterns[14924] = 29'b0_011101001001_100_1_001110100100;
      patterns[14925] = 29'b0_011101001001_101_0_100111010010;
      patterns[14926] = 29'b0_011101001001_110_0_011101001001;
      patterns[14927] = 29'b0_011101001001_111_0_011101001001;
      patterns[14928] = 29'b0_011101001010_000_0_011101001010;
      patterns[14929] = 29'b0_011101001010_001_0_001010011101;
      patterns[14930] = 29'b0_011101001010_010_0_111010010100;
      patterns[14931] = 29'b0_011101001010_011_1_110100101000;
      patterns[14932] = 29'b0_011101001010_100_0_001110100101;
      patterns[14933] = 29'b0_011101001010_101_1_000111010010;
      patterns[14934] = 29'b0_011101001010_110_0_011101001010;
      patterns[14935] = 29'b0_011101001010_111_0_011101001010;
      patterns[14936] = 29'b0_011101001011_000_0_011101001011;
      patterns[14937] = 29'b0_011101001011_001_0_001011011101;
      patterns[14938] = 29'b0_011101001011_010_0_111010010110;
      patterns[14939] = 29'b0_011101001011_011_1_110100101100;
      patterns[14940] = 29'b0_011101001011_100_1_001110100101;
      patterns[14941] = 29'b0_011101001011_101_1_100111010010;
      patterns[14942] = 29'b0_011101001011_110_0_011101001011;
      patterns[14943] = 29'b0_011101001011_111_0_011101001011;
      patterns[14944] = 29'b0_011101001100_000_0_011101001100;
      patterns[14945] = 29'b0_011101001100_001_0_001100011101;
      patterns[14946] = 29'b0_011101001100_010_0_111010011000;
      patterns[14947] = 29'b0_011101001100_011_1_110100110000;
      patterns[14948] = 29'b0_011101001100_100_0_001110100110;
      patterns[14949] = 29'b0_011101001100_101_0_000111010011;
      patterns[14950] = 29'b0_011101001100_110_0_011101001100;
      patterns[14951] = 29'b0_011101001100_111_0_011101001100;
      patterns[14952] = 29'b0_011101001101_000_0_011101001101;
      patterns[14953] = 29'b0_011101001101_001_0_001101011101;
      patterns[14954] = 29'b0_011101001101_010_0_111010011010;
      patterns[14955] = 29'b0_011101001101_011_1_110100110100;
      patterns[14956] = 29'b0_011101001101_100_1_001110100110;
      patterns[14957] = 29'b0_011101001101_101_0_100111010011;
      patterns[14958] = 29'b0_011101001101_110_0_011101001101;
      patterns[14959] = 29'b0_011101001101_111_0_011101001101;
      patterns[14960] = 29'b0_011101001110_000_0_011101001110;
      patterns[14961] = 29'b0_011101001110_001_0_001110011101;
      patterns[14962] = 29'b0_011101001110_010_0_111010011100;
      patterns[14963] = 29'b0_011101001110_011_1_110100111000;
      patterns[14964] = 29'b0_011101001110_100_0_001110100111;
      patterns[14965] = 29'b0_011101001110_101_1_000111010011;
      patterns[14966] = 29'b0_011101001110_110_0_011101001110;
      patterns[14967] = 29'b0_011101001110_111_0_011101001110;
      patterns[14968] = 29'b0_011101001111_000_0_011101001111;
      patterns[14969] = 29'b0_011101001111_001_0_001111011101;
      patterns[14970] = 29'b0_011101001111_010_0_111010011110;
      patterns[14971] = 29'b0_011101001111_011_1_110100111100;
      patterns[14972] = 29'b0_011101001111_100_1_001110100111;
      patterns[14973] = 29'b0_011101001111_101_1_100111010011;
      patterns[14974] = 29'b0_011101001111_110_0_011101001111;
      patterns[14975] = 29'b0_011101001111_111_0_011101001111;
      patterns[14976] = 29'b0_011101010000_000_0_011101010000;
      patterns[14977] = 29'b0_011101010000_001_0_010000011101;
      patterns[14978] = 29'b0_011101010000_010_0_111010100000;
      patterns[14979] = 29'b0_011101010000_011_1_110101000000;
      patterns[14980] = 29'b0_011101010000_100_0_001110101000;
      patterns[14981] = 29'b0_011101010000_101_0_000111010100;
      patterns[14982] = 29'b0_011101010000_110_0_011101010000;
      patterns[14983] = 29'b0_011101010000_111_0_011101010000;
      patterns[14984] = 29'b0_011101010001_000_0_011101010001;
      patterns[14985] = 29'b0_011101010001_001_0_010001011101;
      patterns[14986] = 29'b0_011101010001_010_0_111010100010;
      patterns[14987] = 29'b0_011101010001_011_1_110101000100;
      patterns[14988] = 29'b0_011101010001_100_1_001110101000;
      patterns[14989] = 29'b0_011101010001_101_0_100111010100;
      patterns[14990] = 29'b0_011101010001_110_0_011101010001;
      patterns[14991] = 29'b0_011101010001_111_0_011101010001;
      patterns[14992] = 29'b0_011101010010_000_0_011101010010;
      patterns[14993] = 29'b0_011101010010_001_0_010010011101;
      patterns[14994] = 29'b0_011101010010_010_0_111010100100;
      patterns[14995] = 29'b0_011101010010_011_1_110101001000;
      patterns[14996] = 29'b0_011101010010_100_0_001110101001;
      patterns[14997] = 29'b0_011101010010_101_1_000111010100;
      patterns[14998] = 29'b0_011101010010_110_0_011101010010;
      patterns[14999] = 29'b0_011101010010_111_0_011101010010;
      patterns[15000] = 29'b0_011101010011_000_0_011101010011;
      patterns[15001] = 29'b0_011101010011_001_0_010011011101;
      patterns[15002] = 29'b0_011101010011_010_0_111010100110;
      patterns[15003] = 29'b0_011101010011_011_1_110101001100;
      patterns[15004] = 29'b0_011101010011_100_1_001110101001;
      patterns[15005] = 29'b0_011101010011_101_1_100111010100;
      patterns[15006] = 29'b0_011101010011_110_0_011101010011;
      patterns[15007] = 29'b0_011101010011_111_0_011101010011;
      patterns[15008] = 29'b0_011101010100_000_0_011101010100;
      patterns[15009] = 29'b0_011101010100_001_0_010100011101;
      patterns[15010] = 29'b0_011101010100_010_0_111010101000;
      patterns[15011] = 29'b0_011101010100_011_1_110101010000;
      patterns[15012] = 29'b0_011101010100_100_0_001110101010;
      patterns[15013] = 29'b0_011101010100_101_0_000111010101;
      patterns[15014] = 29'b0_011101010100_110_0_011101010100;
      patterns[15015] = 29'b0_011101010100_111_0_011101010100;
      patterns[15016] = 29'b0_011101010101_000_0_011101010101;
      patterns[15017] = 29'b0_011101010101_001_0_010101011101;
      patterns[15018] = 29'b0_011101010101_010_0_111010101010;
      patterns[15019] = 29'b0_011101010101_011_1_110101010100;
      patterns[15020] = 29'b0_011101010101_100_1_001110101010;
      patterns[15021] = 29'b0_011101010101_101_0_100111010101;
      patterns[15022] = 29'b0_011101010101_110_0_011101010101;
      patterns[15023] = 29'b0_011101010101_111_0_011101010101;
      patterns[15024] = 29'b0_011101010110_000_0_011101010110;
      patterns[15025] = 29'b0_011101010110_001_0_010110011101;
      patterns[15026] = 29'b0_011101010110_010_0_111010101100;
      patterns[15027] = 29'b0_011101010110_011_1_110101011000;
      patterns[15028] = 29'b0_011101010110_100_0_001110101011;
      patterns[15029] = 29'b0_011101010110_101_1_000111010101;
      patterns[15030] = 29'b0_011101010110_110_0_011101010110;
      patterns[15031] = 29'b0_011101010110_111_0_011101010110;
      patterns[15032] = 29'b0_011101010111_000_0_011101010111;
      patterns[15033] = 29'b0_011101010111_001_0_010111011101;
      patterns[15034] = 29'b0_011101010111_010_0_111010101110;
      patterns[15035] = 29'b0_011101010111_011_1_110101011100;
      patterns[15036] = 29'b0_011101010111_100_1_001110101011;
      patterns[15037] = 29'b0_011101010111_101_1_100111010101;
      patterns[15038] = 29'b0_011101010111_110_0_011101010111;
      patterns[15039] = 29'b0_011101010111_111_0_011101010111;
      patterns[15040] = 29'b0_011101011000_000_0_011101011000;
      patterns[15041] = 29'b0_011101011000_001_0_011000011101;
      patterns[15042] = 29'b0_011101011000_010_0_111010110000;
      patterns[15043] = 29'b0_011101011000_011_1_110101100000;
      patterns[15044] = 29'b0_011101011000_100_0_001110101100;
      patterns[15045] = 29'b0_011101011000_101_0_000111010110;
      patterns[15046] = 29'b0_011101011000_110_0_011101011000;
      patterns[15047] = 29'b0_011101011000_111_0_011101011000;
      patterns[15048] = 29'b0_011101011001_000_0_011101011001;
      patterns[15049] = 29'b0_011101011001_001_0_011001011101;
      patterns[15050] = 29'b0_011101011001_010_0_111010110010;
      patterns[15051] = 29'b0_011101011001_011_1_110101100100;
      patterns[15052] = 29'b0_011101011001_100_1_001110101100;
      patterns[15053] = 29'b0_011101011001_101_0_100111010110;
      patterns[15054] = 29'b0_011101011001_110_0_011101011001;
      patterns[15055] = 29'b0_011101011001_111_0_011101011001;
      patterns[15056] = 29'b0_011101011010_000_0_011101011010;
      patterns[15057] = 29'b0_011101011010_001_0_011010011101;
      patterns[15058] = 29'b0_011101011010_010_0_111010110100;
      patterns[15059] = 29'b0_011101011010_011_1_110101101000;
      patterns[15060] = 29'b0_011101011010_100_0_001110101101;
      patterns[15061] = 29'b0_011101011010_101_1_000111010110;
      patterns[15062] = 29'b0_011101011010_110_0_011101011010;
      patterns[15063] = 29'b0_011101011010_111_0_011101011010;
      patterns[15064] = 29'b0_011101011011_000_0_011101011011;
      patterns[15065] = 29'b0_011101011011_001_0_011011011101;
      patterns[15066] = 29'b0_011101011011_010_0_111010110110;
      patterns[15067] = 29'b0_011101011011_011_1_110101101100;
      patterns[15068] = 29'b0_011101011011_100_1_001110101101;
      patterns[15069] = 29'b0_011101011011_101_1_100111010110;
      patterns[15070] = 29'b0_011101011011_110_0_011101011011;
      patterns[15071] = 29'b0_011101011011_111_0_011101011011;
      patterns[15072] = 29'b0_011101011100_000_0_011101011100;
      patterns[15073] = 29'b0_011101011100_001_0_011100011101;
      patterns[15074] = 29'b0_011101011100_010_0_111010111000;
      patterns[15075] = 29'b0_011101011100_011_1_110101110000;
      patterns[15076] = 29'b0_011101011100_100_0_001110101110;
      patterns[15077] = 29'b0_011101011100_101_0_000111010111;
      patterns[15078] = 29'b0_011101011100_110_0_011101011100;
      patterns[15079] = 29'b0_011101011100_111_0_011101011100;
      patterns[15080] = 29'b0_011101011101_000_0_011101011101;
      patterns[15081] = 29'b0_011101011101_001_0_011101011101;
      patterns[15082] = 29'b0_011101011101_010_0_111010111010;
      patterns[15083] = 29'b0_011101011101_011_1_110101110100;
      patterns[15084] = 29'b0_011101011101_100_1_001110101110;
      patterns[15085] = 29'b0_011101011101_101_0_100111010111;
      patterns[15086] = 29'b0_011101011101_110_0_011101011101;
      patterns[15087] = 29'b0_011101011101_111_0_011101011101;
      patterns[15088] = 29'b0_011101011110_000_0_011101011110;
      patterns[15089] = 29'b0_011101011110_001_0_011110011101;
      patterns[15090] = 29'b0_011101011110_010_0_111010111100;
      patterns[15091] = 29'b0_011101011110_011_1_110101111000;
      patterns[15092] = 29'b0_011101011110_100_0_001110101111;
      patterns[15093] = 29'b0_011101011110_101_1_000111010111;
      patterns[15094] = 29'b0_011101011110_110_0_011101011110;
      patterns[15095] = 29'b0_011101011110_111_0_011101011110;
      patterns[15096] = 29'b0_011101011111_000_0_011101011111;
      patterns[15097] = 29'b0_011101011111_001_0_011111011101;
      patterns[15098] = 29'b0_011101011111_010_0_111010111110;
      patterns[15099] = 29'b0_011101011111_011_1_110101111100;
      patterns[15100] = 29'b0_011101011111_100_1_001110101111;
      patterns[15101] = 29'b0_011101011111_101_1_100111010111;
      patterns[15102] = 29'b0_011101011111_110_0_011101011111;
      patterns[15103] = 29'b0_011101011111_111_0_011101011111;
      patterns[15104] = 29'b0_011101100000_000_0_011101100000;
      patterns[15105] = 29'b0_011101100000_001_0_100000011101;
      patterns[15106] = 29'b0_011101100000_010_0_111011000000;
      patterns[15107] = 29'b0_011101100000_011_1_110110000000;
      patterns[15108] = 29'b0_011101100000_100_0_001110110000;
      patterns[15109] = 29'b0_011101100000_101_0_000111011000;
      patterns[15110] = 29'b0_011101100000_110_0_011101100000;
      patterns[15111] = 29'b0_011101100000_111_0_011101100000;
      patterns[15112] = 29'b0_011101100001_000_0_011101100001;
      patterns[15113] = 29'b0_011101100001_001_0_100001011101;
      patterns[15114] = 29'b0_011101100001_010_0_111011000010;
      patterns[15115] = 29'b0_011101100001_011_1_110110000100;
      patterns[15116] = 29'b0_011101100001_100_1_001110110000;
      patterns[15117] = 29'b0_011101100001_101_0_100111011000;
      patterns[15118] = 29'b0_011101100001_110_0_011101100001;
      patterns[15119] = 29'b0_011101100001_111_0_011101100001;
      patterns[15120] = 29'b0_011101100010_000_0_011101100010;
      patterns[15121] = 29'b0_011101100010_001_0_100010011101;
      patterns[15122] = 29'b0_011101100010_010_0_111011000100;
      patterns[15123] = 29'b0_011101100010_011_1_110110001000;
      patterns[15124] = 29'b0_011101100010_100_0_001110110001;
      patterns[15125] = 29'b0_011101100010_101_1_000111011000;
      patterns[15126] = 29'b0_011101100010_110_0_011101100010;
      patterns[15127] = 29'b0_011101100010_111_0_011101100010;
      patterns[15128] = 29'b0_011101100011_000_0_011101100011;
      patterns[15129] = 29'b0_011101100011_001_0_100011011101;
      patterns[15130] = 29'b0_011101100011_010_0_111011000110;
      patterns[15131] = 29'b0_011101100011_011_1_110110001100;
      patterns[15132] = 29'b0_011101100011_100_1_001110110001;
      patterns[15133] = 29'b0_011101100011_101_1_100111011000;
      patterns[15134] = 29'b0_011101100011_110_0_011101100011;
      patterns[15135] = 29'b0_011101100011_111_0_011101100011;
      patterns[15136] = 29'b0_011101100100_000_0_011101100100;
      patterns[15137] = 29'b0_011101100100_001_0_100100011101;
      patterns[15138] = 29'b0_011101100100_010_0_111011001000;
      patterns[15139] = 29'b0_011101100100_011_1_110110010000;
      patterns[15140] = 29'b0_011101100100_100_0_001110110010;
      patterns[15141] = 29'b0_011101100100_101_0_000111011001;
      patterns[15142] = 29'b0_011101100100_110_0_011101100100;
      patterns[15143] = 29'b0_011101100100_111_0_011101100100;
      patterns[15144] = 29'b0_011101100101_000_0_011101100101;
      patterns[15145] = 29'b0_011101100101_001_0_100101011101;
      patterns[15146] = 29'b0_011101100101_010_0_111011001010;
      patterns[15147] = 29'b0_011101100101_011_1_110110010100;
      patterns[15148] = 29'b0_011101100101_100_1_001110110010;
      patterns[15149] = 29'b0_011101100101_101_0_100111011001;
      patterns[15150] = 29'b0_011101100101_110_0_011101100101;
      patterns[15151] = 29'b0_011101100101_111_0_011101100101;
      patterns[15152] = 29'b0_011101100110_000_0_011101100110;
      patterns[15153] = 29'b0_011101100110_001_0_100110011101;
      patterns[15154] = 29'b0_011101100110_010_0_111011001100;
      patterns[15155] = 29'b0_011101100110_011_1_110110011000;
      patterns[15156] = 29'b0_011101100110_100_0_001110110011;
      patterns[15157] = 29'b0_011101100110_101_1_000111011001;
      patterns[15158] = 29'b0_011101100110_110_0_011101100110;
      patterns[15159] = 29'b0_011101100110_111_0_011101100110;
      patterns[15160] = 29'b0_011101100111_000_0_011101100111;
      patterns[15161] = 29'b0_011101100111_001_0_100111011101;
      patterns[15162] = 29'b0_011101100111_010_0_111011001110;
      patterns[15163] = 29'b0_011101100111_011_1_110110011100;
      patterns[15164] = 29'b0_011101100111_100_1_001110110011;
      patterns[15165] = 29'b0_011101100111_101_1_100111011001;
      patterns[15166] = 29'b0_011101100111_110_0_011101100111;
      patterns[15167] = 29'b0_011101100111_111_0_011101100111;
      patterns[15168] = 29'b0_011101101000_000_0_011101101000;
      patterns[15169] = 29'b0_011101101000_001_0_101000011101;
      patterns[15170] = 29'b0_011101101000_010_0_111011010000;
      patterns[15171] = 29'b0_011101101000_011_1_110110100000;
      patterns[15172] = 29'b0_011101101000_100_0_001110110100;
      patterns[15173] = 29'b0_011101101000_101_0_000111011010;
      patterns[15174] = 29'b0_011101101000_110_0_011101101000;
      patterns[15175] = 29'b0_011101101000_111_0_011101101000;
      patterns[15176] = 29'b0_011101101001_000_0_011101101001;
      patterns[15177] = 29'b0_011101101001_001_0_101001011101;
      patterns[15178] = 29'b0_011101101001_010_0_111011010010;
      patterns[15179] = 29'b0_011101101001_011_1_110110100100;
      patterns[15180] = 29'b0_011101101001_100_1_001110110100;
      patterns[15181] = 29'b0_011101101001_101_0_100111011010;
      patterns[15182] = 29'b0_011101101001_110_0_011101101001;
      patterns[15183] = 29'b0_011101101001_111_0_011101101001;
      patterns[15184] = 29'b0_011101101010_000_0_011101101010;
      patterns[15185] = 29'b0_011101101010_001_0_101010011101;
      patterns[15186] = 29'b0_011101101010_010_0_111011010100;
      patterns[15187] = 29'b0_011101101010_011_1_110110101000;
      patterns[15188] = 29'b0_011101101010_100_0_001110110101;
      patterns[15189] = 29'b0_011101101010_101_1_000111011010;
      patterns[15190] = 29'b0_011101101010_110_0_011101101010;
      patterns[15191] = 29'b0_011101101010_111_0_011101101010;
      patterns[15192] = 29'b0_011101101011_000_0_011101101011;
      patterns[15193] = 29'b0_011101101011_001_0_101011011101;
      patterns[15194] = 29'b0_011101101011_010_0_111011010110;
      patterns[15195] = 29'b0_011101101011_011_1_110110101100;
      patterns[15196] = 29'b0_011101101011_100_1_001110110101;
      patterns[15197] = 29'b0_011101101011_101_1_100111011010;
      patterns[15198] = 29'b0_011101101011_110_0_011101101011;
      patterns[15199] = 29'b0_011101101011_111_0_011101101011;
      patterns[15200] = 29'b0_011101101100_000_0_011101101100;
      patterns[15201] = 29'b0_011101101100_001_0_101100011101;
      patterns[15202] = 29'b0_011101101100_010_0_111011011000;
      patterns[15203] = 29'b0_011101101100_011_1_110110110000;
      patterns[15204] = 29'b0_011101101100_100_0_001110110110;
      patterns[15205] = 29'b0_011101101100_101_0_000111011011;
      patterns[15206] = 29'b0_011101101100_110_0_011101101100;
      patterns[15207] = 29'b0_011101101100_111_0_011101101100;
      patterns[15208] = 29'b0_011101101101_000_0_011101101101;
      patterns[15209] = 29'b0_011101101101_001_0_101101011101;
      patterns[15210] = 29'b0_011101101101_010_0_111011011010;
      patterns[15211] = 29'b0_011101101101_011_1_110110110100;
      patterns[15212] = 29'b0_011101101101_100_1_001110110110;
      patterns[15213] = 29'b0_011101101101_101_0_100111011011;
      patterns[15214] = 29'b0_011101101101_110_0_011101101101;
      patterns[15215] = 29'b0_011101101101_111_0_011101101101;
      patterns[15216] = 29'b0_011101101110_000_0_011101101110;
      patterns[15217] = 29'b0_011101101110_001_0_101110011101;
      patterns[15218] = 29'b0_011101101110_010_0_111011011100;
      patterns[15219] = 29'b0_011101101110_011_1_110110111000;
      patterns[15220] = 29'b0_011101101110_100_0_001110110111;
      patterns[15221] = 29'b0_011101101110_101_1_000111011011;
      patterns[15222] = 29'b0_011101101110_110_0_011101101110;
      patterns[15223] = 29'b0_011101101110_111_0_011101101110;
      patterns[15224] = 29'b0_011101101111_000_0_011101101111;
      patterns[15225] = 29'b0_011101101111_001_0_101111011101;
      patterns[15226] = 29'b0_011101101111_010_0_111011011110;
      patterns[15227] = 29'b0_011101101111_011_1_110110111100;
      patterns[15228] = 29'b0_011101101111_100_1_001110110111;
      patterns[15229] = 29'b0_011101101111_101_1_100111011011;
      patterns[15230] = 29'b0_011101101111_110_0_011101101111;
      patterns[15231] = 29'b0_011101101111_111_0_011101101111;
      patterns[15232] = 29'b0_011101110000_000_0_011101110000;
      patterns[15233] = 29'b0_011101110000_001_0_110000011101;
      patterns[15234] = 29'b0_011101110000_010_0_111011100000;
      patterns[15235] = 29'b0_011101110000_011_1_110111000000;
      patterns[15236] = 29'b0_011101110000_100_0_001110111000;
      patterns[15237] = 29'b0_011101110000_101_0_000111011100;
      patterns[15238] = 29'b0_011101110000_110_0_011101110000;
      patterns[15239] = 29'b0_011101110000_111_0_011101110000;
      patterns[15240] = 29'b0_011101110001_000_0_011101110001;
      patterns[15241] = 29'b0_011101110001_001_0_110001011101;
      patterns[15242] = 29'b0_011101110001_010_0_111011100010;
      patterns[15243] = 29'b0_011101110001_011_1_110111000100;
      patterns[15244] = 29'b0_011101110001_100_1_001110111000;
      patterns[15245] = 29'b0_011101110001_101_0_100111011100;
      patterns[15246] = 29'b0_011101110001_110_0_011101110001;
      patterns[15247] = 29'b0_011101110001_111_0_011101110001;
      patterns[15248] = 29'b0_011101110010_000_0_011101110010;
      patterns[15249] = 29'b0_011101110010_001_0_110010011101;
      patterns[15250] = 29'b0_011101110010_010_0_111011100100;
      patterns[15251] = 29'b0_011101110010_011_1_110111001000;
      patterns[15252] = 29'b0_011101110010_100_0_001110111001;
      patterns[15253] = 29'b0_011101110010_101_1_000111011100;
      patterns[15254] = 29'b0_011101110010_110_0_011101110010;
      patterns[15255] = 29'b0_011101110010_111_0_011101110010;
      patterns[15256] = 29'b0_011101110011_000_0_011101110011;
      patterns[15257] = 29'b0_011101110011_001_0_110011011101;
      patterns[15258] = 29'b0_011101110011_010_0_111011100110;
      patterns[15259] = 29'b0_011101110011_011_1_110111001100;
      patterns[15260] = 29'b0_011101110011_100_1_001110111001;
      patterns[15261] = 29'b0_011101110011_101_1_100111011100;
      patterns[15262] = 29'b0_011101110011_110_0_011101110011;
      patterns[15263] = 29'b0_011101110011_111_0_011101110011;
      patterns[15264] = 29'b0_011101110100_000_0_011101110100;
      patterns[15265] = 29'b0_011101110100_001_0_110100011101;
      patterns[15266] = 29'b0_011101110100_010_0_111011101000;
      patterns[15267] = 29'b0_011101110100_011_1_110111010000;
      patterns[15268] = 29'b0_011101110100_100_0_001110111010;
      patterns[15269] = 29'b0_011101110100_101_0_000111011101;
      patterns[15270] = 29'b0_011101110100_110_0_011101110100;
      patterns[15271] = 29'b0_011101110100_111_0_011101110100;
      patterns[15272] = 29'b0_011101110101_000_0_011101110101;
      patterns[15273] = 29'b0_011101110101_001_0_110101011101;
      patterns[15274] = 29'b0_011101110101_010_0_111011101010;
      patterns[15275] = 29'b0_011101110101_011_1_110111010100;
      patterns[15276] = 29'b0_011101110101_100_1_001110111010;
      patterns[15277] = 29'b0_011101110101_101_0_100111011101;
      patterns[15278] = 29'b0_011101110101_110_0_011101110101;
      patterns[15279] = 29'b0_011101110101_111_0_011101110101;
      patterns[15280] = 29'b0_011101110110_000_0_011101110110;
      patterns[15281] = 29'b0_011101110110_001_0_110110011101;
      patterns[15282] = 29'b0_011101110110_010_0_111011101100;
      patterns[15283] = 29'b0_011101110110_011_1_110111011000;
      patterns[15284] = 29'b0_011101110110_100_0_001110111011;
      patterns[15285] = 29'b0_011101110110_101_1_000111011101;
      patterns[15286] = 29'b0_011101110110_110_0_011101110110;
      patterns[15287] = 29'b0_011101110110_111_0_011101110110;
      patterns[15288] = 29'b0_011101110111_000_0_011101110111;
      patterns[15289] = 29'b0_011101110111_001_0_110111011101;
      patterns[15290] = 29'b0_011101110111_010_0_111011101110;
      patterns[15291] = 29'b0_011101110111_011_1_110111011100;
      patterns[15292] = 29'b0_011101110111_100_1_001110111011;
      patterns[15293] = 29'b0_011101110111_101_1_100111011101;
      patterns[15294] = 29'b0_011101110111_110_0_011101110111;
      patterns[15295] = 29'b0_011101110111_111_0_011101110111;
      patterns[15296] = 29'b0_011101111000_000_0_011101111000;
      patterns[15297] = 29'b0_011101111000_001_0_111000011101;
      patterns[15298] = 29'b0_011101111000_010_0_111011110000;
      patterns[15299] = 29'b0_011101111000_011_1_110111100000;
      patterns[15300] = 29'b0_011101111000_100_0_001110111100;
      patterns[15301] = 29'b0_011101111000_101_0_000111011110;
      patterns[15302] = 29'b0_011101111000_110_0_011101111000;
      patterns[15303] = 29'b0_011101111000_111_0_011101111000;
      patterns[15304] = 29'b0_011101111001_000_0_011101111001;
      patterns[15305] = 29'b0_011101111001_001_0_111001011101;
      patterns[15306] = 29'b0_011101111001_010_0_111011110010;
      patterns[15307] = 29'b0_011101111001_011_1_110111100100;
      patterns[15308] = 29'b0_011101111001_100_1_001110111100;
      patterns[15309] = 29'b0_011101111001_101_0_100111011110;
      patterns[15310] = 29'b0_011101111001_110_0_011101111001;
      patterns[15311] = 29'b0_011101111001_111_0_011101111001;
      patterns[15312] = 29'b0_011101111010_000_0_011101111010;
      patterns[15313] = 29'b0_011101111010_001_0_111010011101;
      patterns[15314] = 29'b0_011101111010_010_0_111011110100;
      patterns[15315] = 29'b0_011101111010_011_1_110111101000;
      patterns[15316] = 29'b0_011101111010_100_0_001110111101;
      patterns[15317] = 29'b0_011101111010_101_1_000111011110;
      patterns[15318] = 29'b0_011101111010_110_0_011101111010;
      patterns[15319] = 29'b0_011101111010_111_0_011101111010;
      patterns[15320] = 29'b0_011101111011_000_0_011101111011;
      patterns[15321] = 29'b0_011101111011_001_0_111011011101;
      patterns[15322] = 29'b0_011101111011_010_0_111011110110;
      patterns[15323] = 29'b0_011101111011_011_1_110111101100;
      patterns[15324] = 29'b0_011101111011_100_1_001110111101;
      patterns[15325] = 29'b0_011101111011_101_1_100111011110;
      patterns[15326] = 29'b0_011101111011_110_0_011101111011;
      patterns[15327] = 29'b0_011101111011_111_0_011101111011;
      patterns[15328] = 29'b0_011101111100_000_0_011101111100;
      patterns[15329] = 29'b0_011101111100_001_0_111100011101;
      patterns[15330] = 29'b0_011101111100_010_0_111011111000;
      patterns[15331] = 29'b0_011101111100_011_1_110111110000;
      patterns[15332] = 29'b0_011101111100_100_0_001110111110;
      patterns[15333] = 29'b0_011101111100_101_0_000111011111;
      patterns[15334] = 29'b0_011101111100_110_0_011101111100;
      patterns[15335] = 29'b0_011101111100_111_0_011101111100;
      patterns[15336] = 29'b0_011101111101_000_0_011101111101;
      patterns[15337] = 29'b0_011101111101_001_0_111101011101;
      patterns[15338] = 29'b0_011101111101_010_0_111011111010;
      patterns[15339] = 29'b0_011101111101_011_1_110111110100;
      patterns[15340] = 29'b0_011101111101_100_1_001110111110;
      patterns[15341] = 29'b0_011101111101_101_0_100111011111;
      patterns[15342] = 29'b0_011101111101_110_0_011101111101;
      patterns[15343] = 29'b0_011101111101_111_0_011101111101;
      patterns[15344] = 29'b0_011101111110_000_0_011101111110;
      patterns[15345] = 29'b0_011101111110_001_0_111110011101;
      patterns[15346] = 29'b0_011101111110_010_0_111011111100;
      patterns[15347] = 29'b0_011101111110_011_1_110111111000;
      patterns[15348] = 29'b0_011101111110_100_0_001110111111;
      patterns[15349] = 29'b0_011101111110_101_1_000111011111;
      patterns[15350] = 29'b0_011101111110_110_0_011101111110;
      patterns[15351] = 29'b0_011101111110_111_0_011101111110;
      patterns[15352] = 29'b0_011101111111_000_0_011101111111;
      patterns[15353] = 29'b0_011101111111_001_0_111111011101;
      patterns[15354] = 29'b0_011101111111_010_0_111011111110;
      patterns[15355] = 29'b0_011101111111_011_1_110111111100;
      patterns[15356] = 29'b0_011101111111_100_1_001110111111;
      patterns[15357] = 29'b0_011101111111_101_1_100111011111;
      patterns[15358] = 29'b0_011101111111_110_0_011101111111;
      patterns[15359] = 29'b0_011101111111_111_0_011101111111;
      patterns[15360] = 29'b0_011110000000_000_0_011110000000;
      patterns[15361] = 29'b0_011110000000_001_0_000000011110;
      patterns[15362] = 29'b0_011110000000_010_0_111100000000;
      patterns[15363] = 29'b0_011110000000_011_1_111000000000;
      patterns[15364] = 29'b0_011110000000_100_0_001111000000;
      patterns[15365] = 29'b0_011110000000_101_0_000111100000;
      patterns[15366] = 29'b0_011110000000_110_0_011110000000;
      patterns[15367] = 29'b0_011110000000_111_0_011110000000;
      patterns[15368] = 29'b0_011110000001_000_0_011110000001;
      patterns[15369] = 29'b0_011110000001_001_0_000001011110;
      patterns[15370] = 29'b0_011110000001_010_0_111100000010;
      patterns[15371] = 29'b0_011110000001_011_1_111000000100;
      patterns[15372] = 29'b0_011110000001_100_1_001111000000;
      patterns[15373] = 29'b0_011110000001_101_0_100111100000;
      patterns[15374] = 29'b0_011110000001_110_0_011110000001;
      patterns[15375] = 29'b0_011110000001_111_0_011110000001;
      patterns[15376] = 29'b0_011110000010_000_0_011110000010;
      patterns[15377] = 29'b0_011110000010_001_0_000010011110;
      patterns[15378] = 29'b0_011110000010_010_0_111100000100;
      patterns[15379] = 29'b0_011110000010_011_1_111000001000;
      patterns[15380] = 29'b0_011110000010_100_0_001111000001;
      patterns[15381] = 29'b0_011110000010_101_1_000111100000;
      patterns[15382] = 29'b0_011110000010_110_0_011110000010;
      patterns[15383] = 29'b0_011110000010_111_0_011110000010;
      patterns[15384] = 29'b0_011110000011_000_0_011110000011;
      patterns[15385] = 29'b0_011110000011_001_0_000011011110;
      patterns[15386] = 29'b0_011110000011_010_0_111100000110;
      patterns[15387] = 29'b0_011110000011_011_1_111000001100;
      patterns[15388] = 29'b0_011110000011_100_1_001111000001;
      patterns[15389] = 29'b0_011110000011_101_1_100111100000;
      patterns[15390] = 29'b0_011110000011_110_0_011110000011;
      patterns[15391] = 29'b0_011110000011_111_0_011110000011;
      patterns[15392] = 29'b0_011110000100_000_0_011110000100;
      patterns[15393] = 29'b0_011110000100_001_0_000100011110;
      patterns[15394] = 29'b0_011110000100_010_0_111100001000;
      patterns[15395] = 29'b0_011110000100_011_1_111000010000;
      patterns[15396] = 29'b0_011110000100_100_0_001111000010;
      patterns[15397] = 29'b0_011110000100_101_0_000111100001;
      patterns[15398] = 29'b0_011110000100_110_0_011110000100;
      patterns[15399] = 29'b0_011110000100_111_0_011110000100;
      patterns[15400] = 29'b0_011110000101_000_0_011110000101;
      patterns[15401] = 29'b0_011110000101_001_0_000101011110;
      patterns[15402] = 29'b0_011110000101_010_0_111100001010;
      patterns[15403] = 29'b0_011110000101_011_1_111000010100;
      patterns[15404] = 29'b0_011110000101_100_1_001111000010;
      patterns[15405] = 29'b0_011110000101_101_0_100111100001;
      patterns[15406] = 29'b0_011110000101_110_0_011110000101;
      patterns[15407] = 29'b0_011110000101_111_0_011110000101;
      patterns[15408] = 29'b0_011110000110_000_0_011110000110;
      patterns[15409] = 29'b0_011110000110_001_0_000110011110;
      patterns[15410] = 29'b0_011110000110_010_0_111100001100;
      patterns[15411] = 29'b0_011110000110_011_1_111000011000;
      patterns[15412] = 29'b0_011110000110_100_0_001111000011;
      patterns[15413] = 29'b0_011110000110_101_1_000111100001;
      patterns[15414] = 29'b0_011110000110_110_0_011110000110;
      patterns[15415] = 29'b0_011110000110_111_0_011110000110;
      patterns[15416] = 29'b0_011110000111_000_0_011110000111;
      patterns[15417] = 29'b0_011110000111_001_0_000111011110;
      patterns[15418] = 29'b0_011110000111_010_0_111100001110;
      patterns[15419] = 29'b0_011110000111_011_1_111000011100;
      patterns[15420] = 29'b0_011110000111_100_1_001111000011;
      patterns[15421] = 29'b0_011110000111_101_1_100111100001;
      patterns[15422] = 29'b0_011110000111_110_0_011110000111;
      patterns[15423] = 29'b0_011110000111_111_0_011110000111;
      patterns[15424] = 29'b0_011110001000_000_0_011110001000;
      patterns[15425] = 29'b0_011110001000_001_0_001000011110;
      patterns[15426] = 29'b0_011110001000_010_0_111100010000;
      patterns[15427] = 29'b0_011110001000_011_1_111000100000;
      patterns[15428] = 29'b0_011110001000_100_0_001111000100;
      patterns[15429] = 29'b0_011110001000_101_0_000111100010;
      patterns[15430] = 29'b0_011110001000_110_0_011110001000;
      patterns[15431] = 29'b0_011110001000_111_0_011110001000;
      patterns[15432] = 29'b0_011110001001_000_0_011110001001;
      patterns[15433] = 29'b0_011110001001_001_0_001001011110;
      patterns[15434] = 29'b0_011110001001_010_0_111100010010;
      patterns[15435] = 29'b0_011110001001_011_1_111000100100;
      patterns[15436] = 29'b0_011110001001_100_1_001111000100;
      patterns[15437] = 29'b0_011110001001_101_0_100111100010;
      patterns[15438] = 29'b0_011110001001_110_0_011110001001;
      patterns[15439] = 29'b0_011110001001_111_0_011110001001;
      patterns[15440] = 29'b0_011110001010_000_0_011110001010;
      patterns[15441] = 29'b0_011110001010_001_0_001010011110;
      patterns[15442] = 29'b0_011110001010_010_0_111100010100;
      patterns[15443] = 29'b0_011110001010_011_1_111000101000;
      patterns[15444] = 29'b0_011110001010_100_0_001111000101;
      patterns[15445] = 29'b0_011110001010_101_1_000111100010;
      patterns[15446] = 29'b0_011110001010_110_0_011110001010;
      patterns[15447] = 29'b0_011110001010_111_0_011110001010;
      patterns[15448] = 29'b0_011110001011_000_0_011110001011;
      patterns[15449] = 29'b0_011110001011_001_0_001011011110;
      patterns[15450] = 29'b0_011110001011_010_0_111100010110;
      patterns[15451] = 29'b0_011110001011_011_1_111000101100;
      patterns[15452] = 29'b0_011110001011_100_1_001111000101;
      patterns[15453] = 29'b0_011110001011_101_1_100111100010;
      patterns[15454] = 29'b0_011110001011_110_0_011110001011;
      patterns[15455] = 29'b0_011110001011_111_0_011110001011;
      patterns[15456] = 29'b0_011110001100_000_0_011110001100;
      patterns[15457] = 29'b0_011110001100_001_0_001100011110;
      patterns[15458] = 29'b0_011110001100_010_0_111100011000;
      patterns[15459] = 29'b0_011110001100_011_1_111000110000;
      patterns[15460] = 29'b0_011110001100_100_0_001111000110;
      patterns[15461] = 29'b0_011110001100_101_0_000111100011;
      patterns[15462] = 29'b0_011110001100_110_0_011110001100;
      patterns[15463] = 29'b0_011110001100_111_0_011110001100;
      patterns[15464] = 29'b0_011110001101_000_0_011110001101;
      patterns[15465] = 29'b0_011110001101_001_0_001101011110;
      patterns[15466] = 29'b0_011110001101_010_0_111100011010;
      patterns[15467] = 29'b0_011110001101_011_1_111000110100;
      patterns[15468] = 29'b0_011110001101_100_1_001111000110;
      patterns[15469] = 29'b0_011110001101_101_0_100111100011;
      patterns[15470] = 29'b0_011110001101_110_0_011110001101;
      patterns[15471] = 29'b0_011110001101_111_0_011110001101;
      patterns[15472] = 29'b0_011110001110_000_0_011110001110;
      patterns[15473] = 29'b0_011110001110_001_0_001110011110;
      patterns[15474] = 29'b0_011110001110_010_0_111100011100;
      patterns[15475] = 29'b0_011110001110_011_1_111000111000;
      patterns[15476] = 29'b0_011110001110_100_0_001111000111;
      patterns[15477] = 29'b0_011110001110_101_1_000111100011;
      patterns[15478] = 29'b0_011110001110_110_0_011110001110;
      patterns[15479] = 29'b0_011110001110_111_0_011110001110;
      patterns[15480] = 29'b0_011110001111_000_0_011110001111;
      patterns[15481] = 29'b0_011110001111_001_0_001111011110;
      patterns[15482] = 29'b0_011110001111_010_0_111100011110;
      patterns[15483] = 29'b0_011110001111_011_1_111000111100;
      patterns[15484] = 29'b0_011110001111_100_1_001111000111;
      patterns[15485] = 29'b0_011110001111_101_1_100111100011;
      patterns[15486] = 29'b0_011110001111_110_0_011110001111;
      patterns[15487] = 29'b0_011110001111_111_0_011110001111;
      patterns[15488] = 29'b0_011110010000_000_0_011110010000;
      patterns[15489] = 29'b0_011110010000_001_0_010000011110;
      patterns[15490] = 29'b0_011110010000_010_0_111100100000;
      patterns[15491] = 29'b0_011110010000_011_1_111001000000;
      patterns[15492] = 29'b0_011110010000_100_0_001111001000;
      patterns[15493] = 29'b0_011110010000_101_0_000111100100;
      patterns[15494] = 29'b0_011110010000_110_0_011110010000;
      patterns[15495] = 29'b0_011110010000_111_0_011110010000;
      patterns[15496] = 29'b0_011110010001_000_0_011110010001;
      patterns[15497] = 29'b0_011110010001_001_0_010001011110;
      patterns[15498] = 29'b0_011110010001_010_0_111100100010;
      patterns[15499] = 29'b0_011110010001_011_1_111001000100;
      patterns[15500] = 29'b0_011110010001_100_1_001111001000;
      patterns[15501] = 29'b0_011110010001_101_0_100111100100;
      patterns[15502] = 29'b0_011110010001_110_0_011110010001;
      patterns[15503] = 29'b0_011110010001_111_0_011110010001;
      patterns[15504] = 29'b0_011110010010_000_0_011110010010;
      patterns[15505] = 29'b0_011110010010_001_0_010010011110;
      patterns[15506] = 29'b0_011110010010_010_0_111100100100;
      patterns[15507] = 29'b0_011110010010_011_1_111001001000;
      patterns[15508] = 29'b0_011110010010_100_0_001111001001;
      patterns[15509] = 29'b0_011110010010_101_1_000111100100;
      patterns[15510] = 29'b0_011110010010_110_0_011110010010;
      patterns[15511] = 29'b0_011110010010_111_0_011110010010;
      patterns[15512] = 29'b0_011110010011_000_0_011110010011;
      patterns[15513] = 29'b0_011110010011_001_0_010011011110;
      patterns[15514] = 29'b0_011110010011_010_0_111100100110;
      patterns[15515] = 29'b0_011110010011_011_1_111001001100;
      patterns[15516] = 29'b0_011110010011_100_1_001111001001;
      patterns[15517] = 29'b0_011110010011_101_1_100111100100;
      patterns[15518] = 29'b0_011110010011_110_0_011110010011;
      patterns[15519] = 29'b0_011110010011_111_0_011110010011;
      patterns[15520] = 29'b0_011110010100_000_0_011110010100;
      patterns[15521] = 29'b0_011110010100_001_0_010100011110;
      patterns[15522] = 29'b0_011110010100_010_0_111100101000;
      patterns[15523] = 29'b0_011110010100_011_1_111001010000;
      patterns[15524] = 29'b0_011110010100_100_0_001111001010;
      patterns[15525] = 29'b0_011110010100_101_0_000111100101;
      patterns[15526] = 29'b0_011110010100_110_0_011110010100;
      patterns[15527] = 29'b0_011110010100_111_0_011110010100;
      patterns[15528] = 29'b0_011110010101_000_0_011110010101;
      patterns[15529] = 29'b0_011110010101_001_0_010101011110;
      patterns[15530] = 29'b0_011110010101_010_0_111100101010;
      patterns[15531] = 29'b0_011110010101_011_1_111001010100;
      patterns[15532] = 29'b0_011110010101_100_1_001111001010;
      patterns[15533] = 29'b0_011110010101_101_0_100111100101;
      patterns[15534] = 29'b0_011110010101_110_0_011110010101;
      patterns[15535] = 29'b0_011110010101_111_0_011110010101;
      patterns[15536] = 29'b0_011110010110_000_0_011110010110;
      patterns[15537] = 29'b0_011110010110_001_0_010110011110;
      patterns[15538] = 29'b0_011110010110_010_0_111100101100;
      patterns[15539] = 29'b0_011110010110_011_1_111001011000;
      patterns[15540] = 29'b0_011110010110_100_0_001111001011;
      patterns[15541] = 29'b0_011110010110_101_1_000111100101;
      patterns[15542] = 29'b0_011110010110_110_0_011110010110;
      patterns[15543] = 29'b0_011110010110_111_0_011110010110;
      patterns[15544] = 29'b0_011110010111_000_0_011110010111;
      patterns[15545] = 29'b0_011110010111_001_0_010111011110;
      patterns[15546] = 29'b0_011110010111_010_0_111100101110;
      patterns[15547] = 29'b0_011110010111_011_1_111001011100;
      patterns[15548] = 29'b0_011110010111_100_1_001111001011;
      patterns[15549] = 29'b0_011110010111_101_1_100111100101;
      patterns[15550] = 29'b0_011110010111_110_0_011110010111;
      patterns[15551] = 29'b0_011110010111_111_0_011110010111;
      patterns[15552] = 29'b0_011110011000_000_0_011110011000;
      patterns[15553] = 29'b0_011110011000_001_0_011000011110;
      patterns[15554] = 29'b0_011110011000_010_0_111100110000;
      patterns[15555] = 29'b0_011110011000_011_1_111001100000;
      patterns[15556] = 29'b0_011110011000_100_0_001111001100;
      patterns[15557] = 29'b0_011110011000_101_0_000111100110;
      patterns[15558] = 29'b0_011110011000_110_0_011110011000;
      patterns[15559] = 29'b0_011110011000_111_0_011110011000;
      patterns[15560] = 29'b0_011110011001_000_0_011110011001;
      patterns[15561] = 29'b0_011110011001_001_0_011001011110;
      patterns[15562] = 29'b0_011110011001_010_0_111100110010;
      patterns[15563] = 29'b0_011110011001_011_1_111001100100;
      patterns[15564] = 29'b0_011110011001_100_1_001111001100;
      patterns[15565] = 29'b0_011110011001_101_0_100111100110;
      patterns[15566] = 29'b0_011110011001_110_0_011110011001;
      patterns[15567] = 29'b0_011110011001_111_0_011110011001;
      patterns[15568] = 29'b0_011110011010_000_0_011110011010;
      patterns[15569] = 29'b0_011110011010_001_0_011010011110;
      patterns[15570] = 29'b0_011110011010_010_0_111100110100;
      patterns[15571] = 29'b0_011110011010_011_1_111001101000;
      patterns[15572] = 29'b0_011110011010_100_0_001111001101;
      patterns[15573] = 29'b0_011110011010_101_1_000111100110;
      patterns[15574] = 29'b0_011110011010_110_0_011110011010;
      patterns[15575] = 29'b0_011110011010_111_0_011110011010;
      patterns[15576] = 29'b0_011110011011_000_0_011110011011;
      patterns[15577] = 29'b0_011110011011_001_0_011011011110;
      patterns[15578] = 29'b0_011110011011_010_0_111100110110;
      patterns[15579] = 29'b0_011110011011_011_1_111001101100;
      patterns[15580] = 29'b0_011110011011_100_1_001111001101;
      patterns[15581] = 29'b0_011110011011_101_1_100111100110;
      patterns[15582] = 29'b0_011110011011_110_0_011110011011;
      patterns[15583] = 29'b0_011110011011_111_0_011110011011;
      patterns[15584] = 29'b0_011110011100_000_0_011110011100;
      patterns[15585] = 29'b0_011110011100_001_0_011100011110;
      patterns[15586] = 29'b0_011110011100_010_0_111100111000;
      patterns[15587] = 29'b0_011110011100_011_1_111001110000;
      patterns[15588] = 29'b0_011110011100_100_0_001111001110;
      patterns[15589] = 29'b0_011110011100_101_0_000111100111;
      patterns[15590] = 29'b0_011110011100_110_0_011110011100;
      patterns[15591] = 29'b0_011110011100_111_0_011110011100;
      patterns[15592] = 29'b0_011110011101_000_0_011110011101;
      patterns[15593] = 29'b0_011110011101_001_0_011101011110;
      patterns[15594] = 29'b0_011110011101_010_0_111100111010;
      patterns[15595] = 29'b0_011110011101_011_1_111001110100;
      patterns[15596] = 29'b0_011110011101_100_1_001111001110;
      patterns[15597] = 29'b0_011110011101_101_0_100111100111;
      patterns[15598] = 29'b0_011110011101_110_0_011110011101;
      patterns[15599] = 29'b0_011110011101_111_0_011110011101;
      patterns[15600] = 29'b0_011110011110_000_0_011110011110;
      patterns[15601] = 29'b0_011110011110_001_0_011110011110;
      patterns[15602] = 29'b0_011110011110_010_0_111100111100;
      patterns[15603] = 29'b0_011110011110_011_1_111001111000;
      patterns[15604] = 29'b0_011110011110_100_0_001111001111;
      patterns[15605] = 29'b0_011110011110_101_1_000111100111;
      patterns[15606] = 29'b0_011110011110_110_0_011110011110;
      patterns[15607] = 29'b0_011110011110_111_0_011110011110;
      patterns[15608] = 29'b0_011110011111_000_0_011110011111;
      patterns[15609] = 29'b0_011110011111_001_0_011111011110;
      patterns[15610] = 29'b0_011110011111_010_0_111100111110;
      patterns[15611] = 29'b0_011110011111_011_1_111001111100;
      patterns[15612] = 29'b0_011110011111_100_1_001111001111;
      patterns[15613] = 29'b0_011110011111_101_1_100111100111;
      patterns[15614] = 29'b0_011110011111_110_0_011110011111;
      patterns[15615] = 29'b0_011110011111_111_0_011110011111;
      patterns[15616] = 29'b0_011110100000_000_0_011110100000;
      patterns[15617] = 29'b0_011110100000_001_0_100000011110;
      patterns[15618] = 29'b0_011110100000_010_0_111101000000;
      patterns[15619] = 29'b0_011110100000_011_1_111010000000;
      patterns[15620] = 29'b0_011110100000_100_0_001111010000;
      patterns[15621] = 29'b0_011110100000_101_0_000111101000;
      patterns[15622] = 29'b0_011110100000_110_0_011110100000;
      patterns[15623] = 29'b0_011110100000_111_0_011110100000;
      patterns[15624] = 29'b0_011110100001_000_0_011110100001;
      patterns[15625] = 29'b0_011110100001_001_0_100001011110;
      patterns[15626] = 29'b0_011110100001_010_0_111101000010;
      patterns[15627] = 29'b0_011110100001_011_1_111010000100;
      patterns[15628] = 29'b0_011110100001_100_1_001111010000;
      patterns[15629] = 29'b0_011110100001_101_0_100111101000;
      patterns[15630] = 29'b0_011110100001_110_0_011110100001;
      patterns[15631] = 29'b0_011110100001_111_0_011110100001;
      patterns[15632] = 29'b0_011110100010_000_0_011110100010;
      patterns[15633] = 29'b0_011110100010_001_0_100010011110;
      patterns[15634] = 29'b0_011110100010_010_0_111101000100;
      patterns[15635] = 29'b0_011110100010_011_1_111010001000;
      patterns[15636] = 29'b0_011110100010_100_0_001111010001;
      patterns[15637] = 29'b0_011110100010_101_1_000111101000;
      patterns[15638] = 29'b0_011110100010_110_0_011110100010;
      patterns[15639] = 29'b0_011110100010_111_0_011110100010;
      patterns[15640] = 29'b0_011110100011_000_0_011110100011;
      patterns[15641] = 29'b0_011110100011_001_0_100011011110;
      patterns[15642] = 29'b0_011110100011_010_0_111101000110;
      patterns[15643] = 29'b0_011110100011_011_1_111010001100;
      patterns[15644] = 29'b0_011110100011_100_1_001111010001;
      patterns[15645] = 29'b0_011110100011_101_1_100111101000;
      patterns[15646] = 29'b0_011110100011_110_0_011110100011;
      patterns[15647] = 29'b0_011110100011_111_0_011110100011;
      patterns[15648] = 29'b0_011110100100_000_0_011110100100;
      patterns[15649] = 29'b0_011110100100_001_0_100100011110;
      patterns[15650] = 29'b0_011110100100_010_0_111101001000;
      patterns[15651] = 29'b0_011110100100_011_1_111010010000;
      patterns[15652] = 29'b0_011110100100_100_0_001111010010;
      patterns[15653] = 29'b0_011110100100_101_0_000111101001;
      patterns[15654] = 29'b0_011110100100_110_0_011110100100;
      patterns[15655] = 29'b0_011110100100_111_0_011110100100;
      patterns[15656] = 29'b0_011110100101_000_0_011110100101;
      patterns[15657] = 29'b0_011110100101_001_0_100101011110;
      patterns[15658] = 29'b0_011110100101_010_0_111101001010;
      patterns[15659] = 29'b0_011110100101_011_1_111010010100;
      patterns[15660] = 29'b0_011110100101_100_1_001111010010;
      patterns[15661] = 29'b0_011110100101_101_0_100111101001;
      patterns[15662] = 29'b0_011110100101_110_0_011110100101;
      patterns[15663] = 29'b0_011110100101_111_0_011110100101;
      patterns[15664] = 29'b0_011110100110_000_0_011110100110;
      patterns[15665] = 29'b0_011110100110_001_0_100110011110;
      patterns[15666] = 29'b0_011110100110_010_0_111101001100;
      patterns[15667] = 29'b0_011110100110_011_1_111010011000;
      patterns[15668] = 29'b0_011110100110_100_0_001111010011;
      patterns[15669] = 29'b0_011110100110_101_1_000111101001;
      patterns[15670] = 29'b0_011110100110_110_0_011110100110;
      patterns[15671] = 29'b0_011110100110_111_0_011110100110;
      patterns[15672] = 29'b0_011110100111_000_0_011110100111;
      patterns[15673] = 29'b0_011110100111_001_0_100111011110;
      patterns[15674] = 29'b0_011110100111_010_0_111101001110;
      patterns[15675] = 29'b0_011110100111_011_1_111010011100;
      patterns[15676] = 29'b0_011110100111_100_1_001111010011;
      patterns[15677] = 29'b0_011110100111_101_1_100111101001;
      patterns[15678] = 29'b0_011110100111_110_0_011110100111;
      patterns[15679] = 29'b0_011110100111_111_0_011110100111;
      patterns[15680] = 29'b0_011110101000_000_0_011110101000;
      patterns[15681] = 29'b0_011110101000_001_0_101000011110;
      patterns[15682] = 29'b0_011110101000_010_0_111101010000;
      patterns[15683] = 29'b0_011110101000_011_1_111010100000;
      patterns[15684] = 29'b0_011110101000_100_0_001111010100;
      patterns[15685] = 29'b0_011110101000_101_0_000111101010;
      patterns[15686] = 29'b0_011110101000_110_0_011110101000;
      patterns[15687] = 29'b0_011110101000_111_0_011110101000;
      patterns[15688] = 29'b0_011110101001_000_0_011110101001;
      patterns[15689] = 29'b0_011110101001_001_0_101001011110;
      patterns[15690] = 29'b0_011110101001_010_0_111101010010;
      patterns[15691] = 29'b0_011110101001_011_1_111010100100;
      patterns[15692] = 29'b0_011110101001_100_1_001111010100;
      patterns[15693] = 29'b0_011110101001_101_0_100111101010;
      patterns[15694] = 29'b0_011110101001_110_0_011110101001;
      patterns[15695] = 29'b0_011110101001_111_0_011110101001;
      patterns[15696] = 29'b0_011110101010_000_0_011110101010;
      patterns[15697] = 29'b0_011110101010_001_0_101010011110;
      patterns[15698] = 29'b0_011110101010_010_0_111101010100;
      patterns[15699] = 29'b0_011110101010_011_1_111010101000;
      patterns[15700] = 29'b0_011110101010_100_0_001111010101;
      patterns[15701] = 29'b0_011110101010_101_1_000111101010;
      patterns[15702] = 29'b0_011110101010_110_0_011110101010;
      patterns[15703] = 29'b0_011110101010_111_0_011110101010;
      patterns[15704] = 29'b0_011110101011_000_0_011110101011;
      patterns[15705] = 29'b0_011110101011_001_0_101011011110;
      patterns[15706] = 29'b0_011110101011_010_0_111101010110;
      patterns[15707] = 29'b0_011110101011_011_1_111010101100;
      patterns[15708] = 29'b0_011110101011_100_1_001111010101;
      patterns[15709] = 29'b0_011110101011_101_1_100111101010;
      patterns[15710] = 29'b0_011110101011_110_0_011110101011;
      patterns[15711] = 29'b0_011110101011_111_0_011110101011;
      patterns[15712] = 29'b0_011110101100_000_0_011110101100;
      patterns[15713] = 29'b0_011110101100_001_0_101100011110;
      patterns[15714] = 29'b0_011110101100_010_0_111101011000;
      patterns[15715] = 29'b0_011110101100_011_1_111010110000;
      patterns[15716] = 29'b0_011110101100_100_0_001111010110;
      patterns[15717] = 29'b0_011110101100_101_0_000111101011;
      patterns[15718] = 29'b0_011110101100_110_0_011110101100;
      patterns[15719] = 29'b0_011110101100_111_0_011110101100;
      patterns[15720] = 29'b0_011110101101_000_0_011110101101;
      patterns[15721] = 29'b0_011110101101_001_0_101101011110;
      patterns[15722] = 29'b0_011110101101_010_0_111101011010;
      patterns[15723] = 29'b0_011110101101_011_1_111010110100;
      patterns[15724] = 29'b0_011110101101_100_1_001111010110;
      patterns[15725] = 29'b0_011110101101_101_0_100111101011;
      patterns[15726] = 29'b0_011110101101_110_0_011110101101;
      patterns[15727] = 29'b0_011110101101_111_0_011110101101;
      patterns[15728] = 29'b0_011110101110_000_0_011110101110;
      patterns[15729] = 29'b0_011110101110_001_0_101110011110;
      patterns[15730] = 29'b0_011110101110_010_0_111101011100;
      patterns[15731] = 29'b0_011110101110_011_1_111010111000;
      patterns[15732] = 29'b0_011110101110_100_0_001111010111;
      patterns[15733] = 29'b0_011110101110_101_1_000111101011;
      patterns[15734] = 29'b0_011110101110_110_0_011110101110;
      patterns[15735] = 29'b0_011110101110_111_0_011110101110;
      patterns[15736] = 29'b0_011110101111_000_0_011110101111;
      patterns[15737] = 29'b0_011110101111_001_0_101111011110;
      patterns[15738] = 29'b0_011110101111_010_0_111101011110;
      patterns[15739] = 29'b0_011110101111_011_1_111010111100;
      patterns[15740] = 29'b0_011110101111_100_1_001111010111;
      patterns[15741] = 29'b0_011110101111_101_1_100111101011;
      patterns[15742] = 29'b0_011110101111_110_0_011110101111;
      patterns[15743] = 29'b0_011110101111_111_0_011110101111;
      patterns[15744] = 29'b0_011110110000_000_0_011110110000;
      patterns[15745] = 29'b0_011110110000_001_0_110000011110;
      patterns[15746] = 29'b0_011110110000_010_0_111101100000;
      patterns[15747] = 29'b0_011110110000_011_1_111011000000;
      patterns[15748] = 29'b0_011110110000_100_0_001111011000;
      patterns[15749] = 29'b0_011110110000_101_0_000111101100;
      patterns[15750] = 29'b0_011110110000_110_0_011110110000;
      patterns[15751] = 29'b0_011110110000_111_0_011110110000;
      patterns[15752] = 29'b0_011110110001_000_0_011110110001;
      patterns[15753] = 29'b0_011110110001_001_0_110001011110;
      patterns[15754] = 29'b0_011110110001_010_0_111101100010;
      patterns[15755] = 29'b0_011110110001_011_1_111011000100;
      patterns[15756] = 29'b0_011110110001_100_1_001111011000;
      patterns[15757] = 29'b0_011110110001_101_0_100111101100;
      patterns[15758] = 29'b0_011110110001_110_0_011110110001;
      patterns[15759] = 29'b0_011110110001_111_0_011110110001;
      patterns[15760] = 29'b0_011110110010_000_0_011110110010;
      patterns[15761] = 29'b0_011110110010_001_0_110010011110;
      patterns[15762] = 29'b0_011110110010_010_0_111101100100;
      patterns[15763] = 29'b0_011110110010_011_1_111011001000;
      patterns[15764] = 29'b0_011110110010_100_0_001111011001;
      patterns[15765] = 29'b0_011110110010_101_1_000111101100;
      patterns[15766] = 29'b0_011110110010_110_0_011110110010;
      patterns[15767] = 29'b0_011110110010_111_0_011110110010;
      patterns[15768] = 29'b0_011110110011_000_0_011110110011;
      patterns[15769] = 29'b0_011110110011_001_0_110011011110;
      patterns[15770] = 29'b0_011110110011_010_0_111101100110;
      patterns[15771] = 29'b0_011110110011_011_1_111011001100;
      patterns[15772] = 29'b0_011110110011_100_1_001111011001;
      patterns[15773] = 29'b0_011110110011_101_1_100111101100;
      patterns[15774] = 29'b0_011110110011_110_0_011110110011;
      patterns[15775] = 29'b0_011110110011_111_0_011110110011;
      patterns[15776] = 29'b0_011110110100_000_0_011110110100;
      patterns[15777] = 29'b0_011110110100_001_0_110100011110;
      patterns[15778] = 29'b0_011110110100_010_0_111101101000;
      patterns[15779] = 29'b0_011110110100_011_1_111011010000;
      patterns[15780] = 29'b0_011110110100_100_0_001111011010;
      patterns[15781] = 29'b0_011110110100_101_0_000111101101;
      patterns[15782] = 29'b0_011110110100_110_0_011110110100;
      patterns[15783] = 29'b0_011110110100_111_0_011110110100;
      patterns[15784] = 29'b0_011110110101_000_0_011110110101;
      patterns[15785] = 29'b0_011110110101_001_0_110101011110;
      patterns[15786] = 29'b0_011110110101_010_0_111101101010;
      patterns[15787] = 29'b0_011110110101_011_1_111011010100;
      patterns[15788] = 29'b0_011110110101_100_1_001111011010;
      patterns[15789] = 29'b0_011110110101_101_0_100111101101;
      patterns[15790] = 29'b0_011110110101_110_0_011110110101;
      patterns[15791] = 29'b0_011110110101_111_0_011110110101;
      patterns[15792] = 29'b0_011110110110_000_0_011110110110;
      patterns[15793] = 29'b0_011110110110_001_0_110110011110;
      patterns[15794] = 29'b0_011110110110_010_0_111101101100;
      patterns[15795] = 29'b0_011110110110_011_1_111011011000;
      patterns[15796] = 29'b0_011110110110_100_0_001111011011;
      patterns[15797] = 29'b0_011110110110_101_1_000111101101;
      patterns[15798] = 29'b0_011110110110_110_0_011110110110;
      patterns[15799] = 29'b0_011110110110_111_0_011110110110;
      patterns[15800] = 29'b0_011110110111_000_0_011110110111;
      patterns[15801] = 29'b0_011110110111_001_0_110111011110;
      patterns[15802] = 29'b0_011110110111_010_0_111101101110;
      patterns[15803] = 29'b0_011110110111_011_1_111011011100;
      patterns[15804] = 29'b0_011110110111_100_1_001111011011;
      patterns[15805] = 29'b0_011110110111_101_1_100111101101;
      patterns[15806] = 29'b0_011110110111_110_0_011110110111;
      patterns[15807] = 29'b0_011110110111_111_0_011110110111;
      patterns[15808] = 29'b0_011110111000_000_0_011110111000;
      patterns[15809] = 29'b0_011110111000_001_0_111000011110;
      patterns[15810] = 29'b0_011110111000_010_0_111101110000;
      patterns[15811] = 29'b0_011110111000_011_1_111011100000;
      patterns[15812] = 29'b0_011110111000_100_0_001111011100;
      patterns[15813] = 29'b0_011110111000_101_0_000111101110;
      patterns[15814] = 29'b0_011110111000_110_0_011110111000;
      patterns[15815] = 29'b0_011110111000_111_0_011110111000;
      patterns[15816] = 29'b0_011110111001_000_0_011110111001;
      patterns[15817] = 29'b0_011110111001_001_0_111001011110;
      patterns[15818] = 29'b0_011110111001_010_0_111101110010;
      patterns[15819] = 29'b0_011110111001_011_1_111011100100;
      patterns[15820] = 29'b0_011110111001_100_1_001111011100;
      patterns[15821] = 29'b0_011110111001_101_0_100111101110;
      patterns[15822] = 29'b0_011110111001_110_0_011110111001;
      patterns[15823] = 29'b0_011110111001_111_0_011110111001;
      patterns[15824] = 29'b0_011110111010_000_0_011110111010;
      patterns[15825] = 29'b0_011110111010_001_0_111010011110;
      patterns[15826] = 29'b0_011110111010_010_0_111101110100;
      patterns[15827] = 29'b0_011110111010_011_1_111011101000;
      patterns[15828] = 29'b0_011110111010_100_0_001111011101;
      patterns[15829] = 29'b0_011110111010_101_1_000111101110;
      patterns[15830] = 29'b0_011110111010_110_0_011110111010;
      patterns[15831] = 29'b0_011110111010_111_0_011110111010;
      patterns[15832] = 29'b0_011110111011_000_0_011110111011;
      patterns[15833] = 29'b0_011110111011_001_0_111011011110;
      patterns[15834] = 29'b0_011110111011_010_0_111101110110;
      patterns[15835] = 29'b0_011110111011_011_1_111011101100;
      patterns[15836] = 29'b0_011110111011_100_1_001111011101;
      patterns[15837] = 29'b0_011110111011_101_1_100111101110;
      patterns[15838] = 29'b0_011110111011_110_0_011110111011;
      patterns[15839] = 29'b0_011110111011_111_0_011110111011;
      patterns[15840] = 29'b0_011110111100_000_0_011110111100;
      patterns[15841] = 29'b0_011110111100_001_0_111100011110;
      patterns[15842] = 29'b0_011110111100_010_0_111101111000;
      patterns[15843] = 29'b0_011110111100_011_1_111011110000;
      patterns[15844] = 29'b0_011110111100_100_0_001111011110;
      patterns[15845] = 29'b0_011110111100_101_0_000111101111;
      patterns[15846] = 29'b0_011110111100_110_0_011110111100;
      patterns[15847] = 29'b0_011110111100_111_0_011110111100;
      patterns[15848] = 29'b0_011110111101_000_0_011110111101;
      patterns[15849] = 29'b0_011110111101_001_0_111101011110;
      patterns[15850] = 29'b0_011110111101_010_0_111101111010;
      patterns[15851] = 29'b0_011110111101_011_1_111011110100;
      patterns[15852] = 29'b0_011110111101_100_1_001111011110;
      patterns[15853] = 29'b0_011110111101_101_0_100111101111;
      patterns[15854] = 29'b0_011110111101_110_0_011110111101;
      patterns[15855] = 29'b0_011110111101_111_0_011110111101;
      patterns[15856] = 29'b0_011110111110_000_0_011110111110;
      patterns[15857] = 29'b0_011110111110_001_0_111110011110;
      patterns[15858] = 29'b0_011110111110_010_0_111101111100;
      patterns[15859] = 29'b0_011110111110_011_1_111011111000;
      patterns[15860] = 29'b0_011110111110_100_0_001111011111;
      patterns[15861] = 29'b0_011110111110_101_1_000111101111;
      patterns[15862] = 29'b0_011110111110_110_0_011110111110;
      patterns[15863] = 29'b0_011110111110_111_0_011110111110;
      patterns[15864] = 29'b0_011110111111_000_0_011110111111;
      patterns[15865] = 29'b0_011110111111_001_0_111111011110;
      patterns[15866] = 29'b0_011110111111_010_0_111101111110;
      patterns[15867] = 29'b0_011110111111_011_1_111011111100;
      patterns[15868] = 29'b0_011110111111_100_1_001111011111;
      patterns[15869] = 29'b0_011110111111_101_1_100111101111;
      patterns[15870] = 29'b0_011110111111_110_0_011110111111;
      patterns[15871] = 29'b0_011110111111_111_0_011110111111;
      patterns[15872] = 29'b0_011111000000_000_0_011111000000;
      patterns[15873] = 29'b0_011111000000_001_0_000000011111;
      patterns[15874] = 29'b0_011111000000_010_0_111110000000;
      patterns[15875] = 29'b0_011111000000_011_1_111100000000;
      patterns[15876] = 29'b0_011111000000_100_0_001111100000;
      patterns[15877] = 29'b0_011111000000_101_0_000111110000;
      patterns[15878] = 29'b0_011111000000_110_0_011111000000;
      patterns[15879] = 29'b0_011111000000_111_0_011111000000;
      patterns[15880] = 29'b0_011111000001_000_0_011111000001;
      patterns[15881] = 29'b0_011111000001_001_0_000001011111;
      patterns[15882] = 29'b0_011111000001_010_0_111110000010;
      patterns[15883] = 29'b0_011111000001_011_1_111100000100;
      patterns[15884] = 29'b0_011111000001_100_1_001111100000;
      patterns[15885] = 29'b0_011111000001_101_0_100111110000;
      patterns[15886] = 29'b0_011111000001_110_0_011111000001;
      patterns[15887] = 29'b0_011111000001_111_0_011111000001;
      patterns[15888] = 29'b0_011111000010_000_0_011111000010;
      patterns[15889] = 29'b0_011111000010_001_0_000010011111;
      patterns[15890] = 29'b0_011111000010_010_0_111110000100;
      patterns[15891] = 29'b0_011111000010_011_1_111100001000;
      patterns[15892] = 29'b0_011111000010_100_0_001111100001;
      patterns[15893] = 29'b0_011111000010_101_1_000111110000;
      patterns[15894] = 29'b0_011111000010_110_0_011111000010;
      patterns[15895] = 29'b0_011111000010_111_0_011111000010;
      patterns[15896] = 29'b0_011111000011_000_0_011111000011;
      patterns[15897] = 29'b0_011111000011_001_0_000011011111;
      patterns[15898] = 29'b0_011111000011_010_0_111110000110;
      patterns[15899] = 29'b0_011111000011_011_1_111100001100;
      patterns[15900] = 29'b0_011111000011_100_1_001111100001;
      patterns[15901] = 29'b0_011111000011_101_1_100111110000;
      patterns[15902] = 29'b0_011111000011_110_0_011111000011;
      patterns[15903] = 29'b0_011111000011_111_0_011111000011;
      patterns[15904] = 29'b0_011111000100_000_0_011111000100;
      patterns[15905] = 29'b0_011111000100_001_0_000100011111;
      patterns[15906] = 29'b0_011111000100_010_0_111110001000;
      patterns[15907] = 29'b0_011111000100_011_1_111100010000;
      patterns[15908] = 29'b0_011111000100_100_0_001111100010;
      patterns[15909] = 29'b0_011111000100_101_0_000111110001;
      patterns[15910] = 29'b0_011111000100_110_0_011111000100;
      patterns[15911] = 29'b0_011111000100_111_0_011111000100;
      patterns[15912] = 29'b0_011111000101_000_0_011111000101;
      patterns[15913] = 29'b0_011111000101_001_0_000101011111;
      patterns[15914] = 29'b0_011111000101_010_0_111110001010;
      patterns[15915] = 29'b0_011111000101_011_1_111100010100;
      patterns[15916] = 29'b0_011111000101_100_1_001111100010;
      patterns[15917] = 29'b0_011111000101_101_0_100111110001;
      patterns[15918] = 29'b0_011111000101_110_0_011111000101;
      patterns[15919] = 29'b0_011111000101_111_0_011111000101;
      patterns[15920] = 29'b0_011111000110_000_0_011111000110;
      patterns[15921] = 29'b0_011111000110_001_0_000110011111;
      patterns[15922] = 29'b0_011111000110_010_0_111110001100;
      patterns[15923] = 29'b0_011111000110_011_1_111100011000;
      patterns[15924] = 29'b0_011111000110_100_0_001111100011;
      patterns[15925] = 29'b0_011111000110_101_1_000111110001;
      patterns[15926] = 29'b0_011111000110_110_0_011111000110;
      patterns[15927] = 29'b0_011111000110_111_0_011111000110;
      patterns[15928] = 29'b0_011111000111_000_0_011111000111;
      patterns[15929] = 29'b0_011111000111_001_0_000111011111;
      patterns[15930] = 29'b0_011111000111_010_0_111110001110;
      patterns[15931] = 29'b0_011111000111_011_1_111100011100;
      patterns[15932] = 29'b0_011111000111_100_1_001111100011;
      patterns[15933] = 29'b0_011111000111_101_1_100111110001;
      patterns[15934] = 29'b0_011111000111_110_0_011111000111;
      patterns[15935] = 29'b0_011111000111_111_0_011111000111;
      patterns[15936] = 29'b0_011111001000_000_0_011111001000;
      patterns[15937] = 29'b0_011111001000_001_0_001000011111;
      patterns[15938] = 29'b0_011111001000_010_0_111110010000;
      patterns[15939] = 29'b0_011111001000_011_1_111100100000;
      patterns[15940] = 29'b0_011111001000_100_0_001111100100;
      patterns[15941] = 29'b0_011111001000_101_0_000111110010;
      patterns[15942] = 29'b0_011111001000_110_0_011111001000;
      patterns[15943] = 29'b0_011111001000_111_0_011111001000;
      patterns[15944] = 29'b0_011111001001_000_0_011111001001;
      patterns[15945] = 29'b0_011111001001_001_0_001001011111;
      patterns[15946] = 29'b0_011111001001_010_0_111110010010;
      patterns[15947] = 29'b0_011111001001_011_1_111100100100;
      patterns[15948] = 29'b0_011111001001_100_1_001111100100;
      patterns[15949] = 29'b0_011111001001_101_0_100111110010;
      patterns[15950] = 29'b0_011111001001_110_0_011111001001;
      patterns[15951] = 29'b0_011111001001_111_0_011111001001;
      patterns[15952] = 29'b0_011111001010_000_0_011111001010;
      patterns[15953] = 29'b0_011111001010_001_0_001010011111;
      patterns[15954] = 29'b0_011111001010_010_0_111110010100;
      patterns[15955] = 29'b0_011111001010_011_1_111100101000;
      patterns[15956] = 29'b0_011111001010_100_0_001111100101;
      patterns[15957] = 29'b0_011111001010_101_1_000111110010;
      patterns[15958] = 29'b0_011111001010_110_0_011111001010;
      patterns[15959] = 29'b0_011111001010_111_0_011111001010;
      patterns[15960] = 29'b0_011111001011_000_0_011111001011;
      patterns[15961] = 29'b0_011111001011_001_0_001011011111;
      patterns[15962] = 29'b0_011111001011_010_0_111110010110;
      patterns[15963] = 29'b0_011111001011_011_1_111100101100;
      patterns[15964] = 29'b0_011111001011_100_1_001111100101;
      patterns[15965] = 29'b0_011111001011_101_1_100111110010;
      patterns[15966] = 29'b0_011111001011_110_0_011111001011;
      patterns[15967] = 29'b0_011111001011_111_0_011111001011;
      patterns[15968] = 29'b0_011111001100_000_0_011111001100;
      patterns[15969] = 29'b0_011111001100_001_0_001100011111;
      patterns[15970] = 29'b0_011111001100_010_0_111110011000;
      patterns[15971] = 29'b0_011111001100_011_1_111100110000;
      patterns[15972] = 29'b0_011111001100_100_0_001111100110;
      patterns[15973] = 29'b0_011111001100_101_0_000111110011;
      patterns[15974] = 29'b0_011111001100_110_0_011111001100;
      patterns[15975] = 29'b0_011111001100_111_0_011111001100;
      patterns[15976] = 29'b0_011111001101_000_0_011111001101;
      patterns[15977] = 29'b0_011111001101_001_0_001101011111;
      patterns[15978] = 29'b0_011111001101_010_0_111110011010;
      patterns[15979] = 29'b0_011111001101_011_1_111100110100;
      patterns[15980] = 29'b0_011111001101_100_1_001111100110;
      patterns[15981] = 29'b0_011111001101_101_0_100111110011;
      patterns[15982] = 29'b0_011111001101_110_0_011111001101;
      patterns[15983] = 29'b0_011111001101_111_0_011111001101;
      patterns[15984] = 29'b0_011111001110_000_0_011111001110;
      patterns[15985] = 29'b0_011111001110_001_0_001110011111;
      patterns[15986] = 29'b0_011111001110_010_0_111110011100;
      patterns[15987] = 29'b0_011111001110_011_1_111100111000;
      patterns[15988] = 29'b0_011111001110_100_0_001111100111;
      patterns[15989] = 29'b0_011111001110_101_1_000111110011;
      patterns[15990] = 29'b0_011111001110_110_0_011111001110;
      patterns[15991] = 29'b0_011111001110_111_0_011111001110;
      patterns[15992] = 29'b0_011111001111_000_0_011111001111;
      patterns[15993] = 29'b0_011111001111_001_0_001111011111;
      patterns[15994] = 29'b0_011111001111_010_0_111110011110;
      patterns[15995] = 29'b0_011111001111_011_1_111100111100;
      patterns[15996] = 29'b0_011111001111_100_1_001111100111;
      patterns[15997] = 29'b0_011111001111_101_1_100111110011;
      patterns[15998] = 29'b0_011111001111_110_0_011111001111;
      patterns[15999] = 29'b0_011111001111_111_0_011111001111;
      patterns[16000] = 29'b0_011111010000_000_0_011111010000;
      patterns[16001] = 29'b0_011111010000_001_0_010000011111;
      patterns[16002] = 29'b0_011111010000_010_0_111110100000;
      patterns[16003] = 29'b0_011111010000_011_1_111101000000;
      patterns[16004] = 29'b0_011111010000_100_0_001111101000;
      patterns[16005] = 29'b0_011111010000_101_0_000111110100;
      patterns[16006] = 29'b0_011111010000_110_0_011111010000;
      patterns[16007] = 29'b0_011111010000_111_0_011111010000;
      patterns[16008] = 29'b0_011111010001_000_0_011111010001;
      patterns[16009] = 29'b0_011111010001_001_0_010001011111;
      patterns[16010] = 29'b0_011111010001_010_0_111110100010;
      patterns[16011] = 29'b0_011111010001_011_1_111101000100;
      patterns[16012] = 29'b0_011111010001_100_1_001111101000;
      patterns[16013] = 29'b0_011111010001_101_0_100111110100;
      patterns[16014] = 29'b0_011111010001_110_0_011111010001;
      patterns[16015] = 29'b0_011111010001_111_0_011111010001;
      patterns[16016] = 29'b0_011111010010_000_0_011111010010;
      patterns[16017] = 29'b0_011111010010_001_0_010010011111;
      patterns[16018] = 29'b0_011111010010_010_0_111110100100;
      patterns[16019] = 29'b0_011111010010_011_1_111101001000;
      patterns[16020] = 29'b0_011111010010_100_0_001111101001;
      patterns[16021] = 29'b0_011111010010_101_1_000111110100;
      patterns[16022] = 29'b0_011111010010_110_0_011111010010;
      patterns[16023] = 29'b0_011111010010_111_0_011111010010;
      patterns[16024] = 29'b0_011111010011_000_0_011111010011;
      patterns[16025] = 29'b0_011111010011_001_0_010011011111;
      patterns[16026] = 29'b0_011111010011_010_0_111110100110;
      patterns[16027] = 29'b0_011111010011_011_1_111101001100;
      patterns[16028] = 29'b0_011111010011_100_1_001111101001;
      patterns[16029] = 29'b0_011111010011_101_1_100111110100;
      patterns[16030] = 29'b0_011111010011_110_0_011111010011;
      patterns[16031] = 29'b0_011111010011_111_0_011111010011;
      patterns[16032] = 29'b0_011111010100_000_0_011111010100;
      patterns[16033] = 29'b0_011111010100_001_0_010100011111;
      patterns[16034] = 29'b0_011111010100_010_0_111110101000;
      patterns[16035] = 29'b0_011111010100_011_1_111101010000;
      patterns[16036] = 29'b0_011111010100_100_0_001111101010;
      patterns[16037] = 29'b0_011111010100_101_0_000111110101;
      patterns[16038] = 29'b0_011111010100_110_0_011111010100;
      patterns[16039] = 29'b0_011111010100_111_0_011111010100;
      patterns[16040] = 29'b0_011111010101_000_0_011111010101;
      patterns[16041] = 29'b0_011111010101_001_0_010101011111;
      patterns[16042] = 29'b0_011111010101_010_0_111110101010;
      patterns[16043] = 29'b0_011111010101_011_1_111101010100;
      patterns[16044] = 29'b0_011111010101_100_1_001111101010;
      patterns[16045] = 29'b0_011111010101_101_0_100111110101;
      patterns[16046] = 29'b0_011111010101_110_0_011111010101;
      patterns[16047] = 29'b0_011111010101_111_0_011111010101;
      patterns[16048] = 29'b0_011111010110_000_0_011111010110;
      patterns[16049] = 29'b0_011111010110_001_0_010110011111;
      patterns[16050] = 29'b0_011111010110_010_0_111110101100;
      patterns[16051] = 29'b0_011111010110_011_1_111101011000;
      patterns[16052] = 29'b0_011111010110_100_0_001111101011;
      patterns[16053] = 29'b0_011111010110_101_1_000111110101;
      patterns[16054] = 29'b0_011111010110_110_0_011111010110;
      patterns[16055] = 29'b0_011111010110_111_0_011111010110;
      patterns[16056] = 29'b0_011111010111_000_0_011111010111;
      patterns[16057] = 29'b0_011111010111_001_0_010111011111;
      patterns[16058] = 29'b0_011111010111_010_0_111110101110;
      patterns[16059] = 29'b0_011111010111_011_1_111101011100;
      patterns[16060] = 29'b0_011111010111_100_1_001111101011;
      patterns[16061] = 29'b0_011111010111_101_1_100111110101;
      patterns[16062] = 29'b0_011111010111_110_0_011111010111;
      patterns[16063] = 29'b0_011111010111_111_0_011111010111;
      patterns[16064] = 29'b0_011111011000_000_0_011111011000;
      patterns[16065] = 29'b0_011111011000_001_0_011000011111;
      patterns[16066] = 29'b0_011111011000_010_0_111110110000;
      patterns[16067] = 29'b0_011111011000_011_1_111101100000;
      patterns[16068] = 29'b0_011111011000_100_0_001111101100;
      patterns[16069] = 29'b0_011111011000_101_0_000111110110;
      patterns[16070] = 29'b0_011111011000_110_0_011111011000;
      patterns[16071] = 29'b0_011111011000_111_0_011111011000;
      patterns[16072] = 29'b0_011111011001_000_0_011111011001;
      patterns[16073] = 29'b0_011111011001_001_0_011001011111;
      patterns[16074] = 29'b0_011111011001_010_0_111110110010;
      patterns[16075] = 29'b0_011111011001_011_1_111101100100;
      patterns[16076] = 29'b0_011111011001_100_1_001111101100;
      patterns[16077] = 29'b0_011111011001_101_0_100111110110;
      patterns[16078] = 29'b0_011111011001_110_0_011111011001;
      patterns[16079] = 29'b0_011111011001_111_0_011111011001;
      patterns[16080] = 29'b0_011111011010_000_0_011111011010;
      patterns[16081] = 29'b0_011111011010_001_0_011010011111;
      patterns[16082] = 29'b0_011111011010_010_0_111110110100;
      patterns[16083] = 29'b0_011111011010_011_1_111101101000;
      patterns[16084] = 29'b0_011111011010_100_0_001111101101;
      patterns[16085] = 29'b0_011111011010_101_1_000111110110;
      patterns[16086] = 29'b0_011111011010_110_0_011111011010;
      patterns[16087] = 29'b0_011111011010_111_0_011111011010;
      patterns[16088] = 29'b0_011111011011_000_0_011111011011;
      patterns[16089] = 29'b0_011111011011_001_0_011011011111;
      patterns[16090] = 29'b0_011111011011_010_0_111110110110;
      patterns[16091] = 29'b0_011111011011_011_1_111101101100;
      patterns[16092] = 29'b0_011111011011_100_1_001111101101;
      patterns[16093] = 29'b0_011111011011_101_1_100111110110;
      patterns[16094] = 29'b0_011111011011_110_0_011111011011;
      patterns[16095] = 29'b0_011111011011_111_0_011111011011;
      patterns[16096] = 29'b0_011111011100_000_0_011111011100;
      patterns[16097] = 29'b0_011111011100_001_0_011100011111;
      patterns[16098] = 29'b0_011111011100_010_0_111110111000;
      patterns[16099] = 29'b0_011111011100_011_1_111101110000;
      patterns[16100] = 29'b0_011111011100_100_0_001111101110;
      patterns[16101] = 29'b0_011111011100_101_0_000111110111;
      patterns[16102] = 29'b0_011111011100_110_0_011111011100;
      patterns[16103] = 29'b0_011111011100_111_0_011111011100;
      patterns[16104] = 29'b0_011111011101_000_0_011111011101;
      patterns[16105] = 29'b0_011111011101_001_0_011101011111;
      patterns[16106] = 29'b0_011111011101_010_0_111110111010;
      patterns[16107] = 29'b0_011111011101_011_1_111101110100;
      patterns[16108] = 29'b0_011111011101_100_1_001111101110;
      patterns[16109] = 29'b0_011111011101_101_0_100111110111;
      patterns[16110] = 29'b0_011111011101_110_0_011111011101;
      patterns[16111] = 29'b0_011111011101_111_0_011111011101;
      patterns[16112] = 29'b0_011111011110_000_0_011111011110;
      patterns[16113] = 29'b0_011111011110_001_0_011110011111;
      patterns[16114] = 29'b0_011111011110_010_0_111110111100;
      patterns[16115] = 29'b0_011111011110_011_1_111101111000;
      patterns[16116] = 29'b0_011111011110_100_0_001111101111;
      patterns[16117] = 29'b0_011111011110_101_1_000111110111;
      patterns[16118] = 29'b0_011111011110_110_0_011111011110;
      patterns[16119] = 29'b0_011111011110_111_0_011111011110;
      patterns[16120] = 29'b0_011111011111_000_0_011111011111;
      patterns[16121] = 29'b0_011111011111_001_0_011111011111;
      patterns[16122] = 29'b0_011111011111_010_0_111110111110;
      patterns[16123] = 29'b0_011111011111_011_1_111101111100;
      patterns[16124] = 29'b0_011111011111_100_1_001111101111;
      patterns[16125] = 29'b0_011111011111_101_1_100111110111;
      patterns[16126] = 29'b0_011111011111_110_0_011111011111;
      patterns[16127] = 29'b0_011111011111_111_0_011111011111;
      patterns[16128] = 29'b0_011111100000_000_0_011111100000;
      patterns[16129] = 29'b0_011111100000_001_0_100000011111;
      patterns[16130] = 29'b0_011111100000_010_0_111111000000;
      patterns[16131] = 29'b0_011111100000_011_1_111110000000;
      patterns[16132] = 29'b0_011111100000_100_0_001111110000;
      patterns[16133] = 29'b0_011111100000_101_0_000111111000;
      patterns[16134] = 29'b0_011111100000_110_0_011111100000;
      patterns[16135] = 29'b0_011111100000_111_0_011111100000;
      patterns[16136] = 29'b0_011111100001_000_0_011111100001;
      patterns[16137] = 29'b0_011111100001_001_0_100001011111;
      patterns[16138] = 29'b0_011111100001_010_0_111111000010;
      patterns[16139] = 29'b0_011111100001_011_1_111110000100;
      patterns[16140] = 29'b0_011111100001_100_1_001111110000;
      patterns[16141] = 29'b0_011111100001_101_0_100111111000;
      patterns[16142] = 29'b0_011111100001_110_0_011111100001;
      patterns[16143] = 29'b0_011111100001_111_0_011111100001;
      patterns[16144] = 29'b0_011111100010_000_0_011111100010;
      patterns[16145] = 29'b0_011111100010_001_0_100010011111;
      patterns[16146] = 29'b0_011111100010_010_0_111111000100;
      patterns[16147] = 29'b0_011111100010_011_1_111110001000;
      patterns[16148] = 29'b0_011111100010_100_0_001111110001;
      patterns[16149] = 29'b0_011111100010_101_1_000111111000;
      patterns[16150] = 29'b0_011111100010_110_0_011111100010;
      patterns[16151] = 29'b0_011111100010_111_0_011111100010;
      patterns[16152] = 29'b0_011111100011_000_0_011111100011;
      patterns[16153] = 29'b0_011111100011_001_0_100011011111;
      patterns[16154] = 29'b0_011111100011_010_0_111111000110;
      patterns[16155] = 29'b0_011111100011_011_1_111110001100;
      patterns[16156] = 29'b0_011111100011_100_1_001111110001;
      patterns[16157] = 29'b0_011111100011_101_1_100111111000;
      patterns[16158] = 29'b0_011111100011_110_0_011111100011;
      patterns[16159] = 29'b0_011111100011_111_0_011111100011;
      patterns[16160] = 29'b0_011111100100_000_0_011111100100;
      patterns[16161] = 29'b0_011111100100_001_0_100100011111;
      patterns[16162] = 29'b0_011111100100_010_0_111111001000;
      patterns[16163] = 29'b0_011111100100_011_1_111110010000;
      patterns[16164] = 29'b0_011111100100_100_0_001111110010;
      patterns[16165] = 29'b0_011111100100_101_0_000111111001;
      patterns[16166] = 29'b0_011111100100_110_0_011111100100;
      patterns[16167] = 29'b0_011111100100_111_0_011111100100;
      patterns[16168] = 29'b0_011111100101_000_0_011111100101;
      patterns[16169] = 29'b0_011111100101_001_0_100101011111;
      patterns[16170] = 29'b0_011111100101_010_0_111111001010;
      patterns[16171] = 29'b0_011111100101_011_1_111110010100;
      patterns[16172] = 29'b0_011111100101_100_1_001111110010;
      patterns[16173] = 29'b0_011111100101_101_0_100111111001;
      patterns[16174] = 29'b0_011111100101_110_0_011111100101;
      patterns[16175] = 29'b0_011111100101_111_0_011111100101;
      patterns[16176] = 29'b0_011111100110_000_0_011111100110;
      patterns[16177] = 29'b0_011111100110_001_0_100110011111;
      patterns[16178] = 29'b0_011111100110_010_0_111111001100;
      patterns[16179] = 29'b0_011111100110_011_1_111110011000;
      patterns[16180] = 29'b0_011111100110_100_0_001111110011;
      patterns[16181] = 29'b0_011111100110_101_1_000111111001;
      patterns[16182] = 29'b0_011111100110_110_0_011111100110;
      patterns[16183] = 29'b0_011111100110_111_0_011111100110;
      patterns[16184] = 29'b0_011111100111_000_0_011111100111;
      patterns[16185] = 29'b0_011111100111_001_0_100111011111;
      patterns[16186] = 29'b0_011111100111_010_0_111111001110;
      patterns[16187] = 29'b0_011111100111_011_1_111110011100;
      patterns[16188] = 29'b0_011111100111_100_1_001111110011;
      patterns[16189] = 29'b0_011111100111_101_1_100111111001;
      patterns[16190] = 29'b0_011111100111_110_0_011111100111;
      patterns[16191] = 29'b0_011111100111_111_0_011111100111;
      patterns[16192] = 29'b0_011111101000_000_0_011111101000;
      patterns[16193] = 29'b0_011111101000_001_0_101000011111;
      patterns[16194] = 29'b0_011111101000_010_0_111111010000;
      patterns[16195] = 29'b0_011111101000_011_1_111110100000;
      patterns[16196] = 29'b0_011111101000_100_0_001111110100;
      patterns[16197] = 29'b0_011111101000_101_0_000111111010;
      patterns[16198] = 29'b0_011111101000_110_0_011111101000;
      patterns[16199] = 29'b0_011111101000_111_0_011111101000;
      patterns[16200] = 29'b0_011111101001_000_0_011111101001;
      patterns[16201] = 29'b0_011111101001_001_0_101001011111;
      patterns[16202] = 29'b0_011111101001_010_0_111111010010;
      patterns[16203] = 29'b0_011111101001_011_1_111110100100;
      patterns[16204] = 29'b0_011111101001_100_1_001111110100;
      patterns[16205] = 29'b0_011111101001_101_0_100111111010;
      patterns[16206] = 29'b0_011111101001_110_0_011111101001;
      patterns[16207] = 29'b0_011111101001_111_0_011111101001;
      patterns[16208] = 29'b0_011111101010_000_0_011111101010;
      patterns[16209] = 29'b0_011111101010_001_0_101010011111;
      patterns[16210] = 29'b0_011111101010_010_0_111111010100;
      patterns[16211] = 29'b0_011111101010_011_1_111110101000;
      patterns[16212] = 29'b0_011111101010_100_0_001111110101;
      patterns[16213] = 29'b0_011111101010_101_1_000111111010;
      patterns[16214] = 29'b0_011111101010_110_0_011111101010;
      patterns[16215] = 29'b0_011111101010_111_0_011111101010;
      patterns[16216] = 29'b0_011111101011_000_0_011111101011;
      patterns[16217] = 29'b0_011111101011_001_0_101011011111;
      patterns[16218] = 29'b0_011111101011_010_0_111111010110;
      patterns[16219] = 29'b0_011111101011_011_1_111110101100;
      patterns[16220] = 29'b0_011111101011_100_1_001111110101;
      patterns[16221] = 29'b0_011111101011_101_1_100111111010;
      patterns[16222] = 29'b0_011111101011_110_0_011111101011;
      patterns[16223] = 29'b0_011111101011_111_0_011111101011;
      patterns[16224] = 29'b0_011111101100_000_0_011111101100;
      patterns[16225] = 29'b0_011111101100_001_0_101100011111;
      patterns[16226] = 29'b0_011111101100_010_0_111111011000;
      patterns[16227] = 29'b0_011111101100_011_1_111110110000;
      patterns[16228] = 29'b0_011111101100_100_0_001111110110;
      patterns[16229] = 29'b0_011111101100_101_0_000111111011;
      patterns[16230] = 29'b0_011111101100_110_0_011111101100;
      patterns[16231] = 29'b0_011111101100_111_0_011111101100;
      patterns[16232] = 29'b0_011111101101_000_0_011111101101;
      patterns[16233] = 29'b0_011111101101_001_0_101101011111;
      patterns[16234] = 29'b0_011111101101_010_0_111111011010;
      patterns[16235] = 29'b0_011111101101_011_1_111110110100;
      patterns[16236] = 29'b0_011111101101_100_1_001111110110;
      patterns[16237] = 29'b0_011111101101_101_0_100111111011;
      patterns[16238] = 29'b0_011111101101_110_0_011111101101;
      patterns[16239] = 29'b0_011111101101_111_0_011111101101;
      patterns[16240] = 29'b0_011111101110_000_0_011111101110;
      patterns[16241] = 29'b0_011111101110_001_0_101110011111;
      patterns[16242] = 29'b0_011111101110_010_0_111111011100;
      patterns[16243] = 29'b0_011111101110_011_1_111110111000;
      patterns[16244] = 29'b0_011111101110_100_0_001111110111;
      patterns[16245] = 29'b0_011111101110_101_1_000111111011;
      patterns[16246] = 29'b0_011111101110_110_0_011111101110;
      patterns[16247] = 29'b0_011111101110_111_0_011111101110;
      patterns[16248] = 29'b0_011111101111_000_0_011111101111;
      patterns[16249] = 29'b0_011111101111_001_0_101111011111;
      patterns[16250] = 29'b0_011111101111_010_0_111111011110;
      patterns[16251] = 29'b0_011111101111_011_1_111110111100;
      patterns[16252] = 29'b0_011111101111_100_1_001111110111;
      patterns[16253] = 29'b0_011111101111_101_1_100111111011;
      patterns[16254] = 29'b0_011111101111_110_0_011111101111;
      patterns[16255] = 29'b0_011111101111_111_0_011111101111;
      patterns[16256] = 29'b0_011111110000_000_0_011111110000;
      patterns[16257] = 29'b0_011111110000_001_0_110000011111;
      patterns[16258] = 29'b0_011111110000_010_0_111111100000;
      patterns[16259] = 29'b0_011111110000_011_1_111111000000;
      patterns[16260] = 29'b0_011111110000_100_0_001111111000;
      patterns[16261] = 29'b0_011111110000_101_0_000111111100;
      patterns[16262] = 29'b0_011111110000_110_0_011111110000;
      patterns[16263] = 29'b0_011111110000_111_0_011111110000;
      patterns[16264] = 29'b0_011111110001_000_0_011111110001;
      patterns[16265] = 29'b0_011111110001_001_0_110001011111;
      patterns[16266] = 29'b0_011111110001_010_0_111111100010;
      patterns[16267] = 29'b0_011111110001_011_1_111111000100;
      patterns[16268] = 29'b0_011111110001_100_1_001111111000;
      patterns[16269] = 29'b0_011111110001_101_0_100111111100;
      patterns[16270] = 29'b0_011111110001_110_0_011111110001;
      patterns[16271] = 29'b0_011111110001_111_0_011111110001;
      patterns[16272] = 29'b0_011111110010_000_0_011111110010;
      patterns[16273] = 29'b0_011111110010_001_0_110010011111;
      patterns[16274] = 29'b0_011111110010_010_0_111111100100;
      patterns[16275] = 29'b0_011111110010_011_1_111111001000;
      patterns[16276] = 29'b0_011111110010_100_0_001111111001;
      patterns[16277] = 29'b0_011111110010_101_1_000111111100;
      patterns[16278] = 29'b0_011111110010_110_0_011111110010;
      patterns[16279] = 29'b0_011111110010_111_0_011111110010;
      patterns[16280] = 29'b0_011111110011_000_0_011111110011;
      patterns[16281] = 29'b0_011111110011_001_0_110011011111;
      patterns[16282] = 29'b0_011111110011_010_0_111111100110;
      patterns[16283] = 29'b0_011111110011_011_1_111111001100;
      patterns[16284] = 29'b0_011111110011_100_1_001111111001;
      patterns[16285] = 29'b0_011111110011_101_1_100111111100;
      patterns[16286] = 29'b0_011111110011_110_0_011111110011;
      patterns[16287] = 29'b0_011111110011_111_0_011111110011;
      patterns[16288] = 29'b0_011111110100_000_0_011111110100;
      patterns[16289] = 29'b0_011111110100_001_0_110100011111;
      patterns[16290] = 29'b0_011111110100_010_0_111111101000;
      patterns[16291] = 29'b0_011111110100_011_1_111111010000;
      patterns[16292] = 29'b0_011111110100_100_0_001111111010;
      patterns[16293] = 29'b0_011111110100_101_0_000111111101;
      patterns[16294] = 29'b0_011111110100_110_0_011111110100;
      patterns[16295] = 29'b0_011111110100_111_0_011111110100;
      patterns[16296] = 29'b0_011111110101_000_0_011111110101;
      patterns[16297] = 29'b0_011111110101_001_0_110101011111;
      patterns[16298] = 29'b0_011111110101_010_0_111111101010;
      patterns[16299] = 29'b0_011111110101_011_1_111111010100;
      patterns[16300] = 29'b0_011111110101_100_1_001111111010;
      patterns[16301] = 29'b0_011111110101_101_0_100111111101;
      patterns[16302] = 29'b0_011111110101_110_0_011111110101;
      patterns[16303] = 29'b0_011111110101_111_0_011111110101;
      patterns[16304] = 29'b0_011111110110_000_0_011111110110;
      patterns[16305] = 29'b0_011111110110_001_0_110110011111;
      patterns[16306] = 29'b0_011111110110_010_0_111111101100;
      patterns[16307] = 29'b0_011111110110_011_1_111111011000;
      patterns[16308] = 29'b0_011111110110_100_0_001111111011;
      patterns[16309] = 29'b0_011111110110_101_1_000111111101;
      patterns[16310] = 29'b0_011111110110_110_0_011111110110;
      patterns[16311] = 29'b0_011111110110_111_0_011111110110;
      patterns[16312] = 29'b0_011111110111_000_0_011111110111;
      patterns[16313] = 29'b0_011111110111_001_0_110111011111;
      patterns[16314] = 29'b0_011111110111_010_0_111111101110;
      patterns[16315] = 29'b0_011111110111_011_1_111111011100;
      patterns[16316] = 29'b0_011111110111_100_1_001111111011;
      patterns[16317] = 29'b0_011111110111_101_1_100111111101;
      patterns[16318] = 29'b0_011111110111_110_0_011111110111;
      patterns[16319] = 29'b0_011111110111_111_0_011111110111;
      patterns[16320] = 29'b0_011111111000_000_0_011111111000;
      patterns[16321] = 29'b0_011111111000_001_0_111000011111;
      patterns[16322] = 29'b0_011111111000_010_0_111111110000;
      patterns[16323] = 29'b0_011111111000_011_1_111111100000;
      patterns[16324] = 29'b0_011111111000_100_0_001111111100;
      patterns[16325] = 29'b0_011111111000_101_0_000111111110;
      patterns[16326] = 29'b0_011111111000_110_0_011111111000;
      patterns[16327] = 29'b0_011111111000_111_0_011111111000;
      patterns[16328] = 29'b0_011111111001_000_0_011111111001;
      patterns[16329] = 29'b0_011111111001_001_0_111001011111;
      patterns[16330] = 29'b0_011111111001_010_0_111111110010;
      patterns[16331] = 29'b0_011111111001_011_1_111111100100;
      patterns[16332] = 29'b0_011111111001_100_1_001111111100;
      patterns[16333] = 29'b0_011111111001_101_0_100111111110;
      patterns[16334] = 29'b0_011111111001_110_0_011111111001;
      patterns[16335] = 29'b0_011111111001_111_0_011111111001;
      patterns[16336] = 29'b0_011111111010_000_0_011111111010;
      patterns[16337] = 29'b0_011111111010_001_0_111010011111;
      patterns[16338] = 29'b0_011111111010_010_0_111111110100;
      patterns[16339] = 29'b0_011111111010_011_1_111111101000;
      patterns[16340] = 29'b0_011111111010_100_0_001111111101;
      patterns[16341] = 29'b0_011111111010_101_1_000111111110;
      patterns[16342] = 29'b0_011111111010_110_0_011111111010;
      patterns[16343] = 29'b0_011111111010_111_0_011111111010;
      patterns[16344] = 29'b0_011111111011_000_0_011111111011;
      patterns[16345] = 29'b0_011111111011_001_0_111011011111;
      patterns[16346] = 29'b0_011111111011_010_0_111111110110;
      patterns[16347] = 29'b0_011111111011_011_1_111111101100;
      patterns[16348] = 29'b0_011111111011_100_1_001111111101;
      patterns[16349] = 29'b0_011111111011_101_1_100111111110;
      patterns[16350] = 29'b0_011111111011_110_0_011111111011;
      patterns[16351] = 29'b0_011111111011_111_0_011111111011;
      patterns[16352] = 29'b0_011111111100_000_0_011111111100;
      patterns[16353] = 29'b0_011111111100_001_0_111100011111;
      patterns[16354] = 29'b0_011111111100_010_0_111111111000;
      patterns[16355] = 29'b0_011111111100_011_1_111111110000;
      patterns[16356] = 29'b0_011111111100_100_0_001111111110;
      patterns[16357] = 29'b0_011111111100_101_0_000111111111;
      patterns[16358] = 29'b0_011111111100_110_0_011111111100;
      patterns[16359] = 29'b0_011111111100_111_0_011111111100;
      patterns[16360] = 29'b0_011111111101_000_0_011111111101;
      patterns[16361] = 29'b0_011111111101_001_0_111101011111;
      patterns[16362] = 29'b0_011111111101_010_0_111111111010;
      patterns[16363] = 29'b0_011111111101_011_1_111111110100;
      patterns[16364] = 29'b0_011111111101_100_1_001111111110;
      patterns[16365] = 29'b0_011111111101_101_0_100111111111;
      patterns[16366] = 29'b0_011111111101_110_0_011111111101;
      patterns[16367] = 29'b0_011111111101_111_0_011111111101;
      patterns[16368] = 29'b0_011111111110_000_0_011111111110;
      patterns[16369] = 29'b0_011111111110_001_0_111110011111;
      patterns[16370] = 29'b0_011111111110_010_0_111111111100;
      patterns[16371] = 29'b0_011111111110_011_1_111111111000;
      patterns[16372] = 29'b0_011111111110_100_0_001111111111;
      patterns[16373] = 29'b0_011111111110_101_1_000111111111;
      patterns[16374] = 29'b0_011111111110_110_0_011111111110;
      patterns[16375] = 29'b0_011111111110_111_0_011111111110;
      patterns[16376] = 29'b0_011111111111_000_0_011111111111;
      patterns[16377] = 29'b0_011111111111_001_0_111111011111;
      patterns[16378] = 29'b0_011111111111_010_0_111111111110;
      patterns[16379] = 29'b0_011111111111_011_1_111111111100;
      patterns[16380] = 29'b0_011111111111_100_1_001111111111;
      patterns[16381] = 29'b0_011111111111_101_1_100111111111;
      patterns[16382] = 29'b0_011111111111_110_0_011111111111;
      patterns[16383] = 29'b0_011111111111_111_0_011111111111;
      patterns[16384] = 29'b0_100000000000_000_0_100000000000;
      patterns[16385] = 29'b0_100000000000_001_0_000000100000;
      patterns[16386] = 29'b0_100000000000_010_1_000000000000;
      patterns[16387] = 29'b0_100000000000_011_0_000000000001;
      patterns[16388] = 29'b0_100000000000_100_0_010000000000;
      patterns[16389] = 29'b0_100000000000_101_0_001000000000;
      patterns[16390] = 29'b0_100000000000_110_0_100000000000;
      patterns[16391] = 29'b0_100000000000_111_0_100000000000;
      patterns[16392] = 29'b0_100000000001_000_0_100000000001;
      patterns[16393] = 29'b0_100000000001_001_0_000001100000;
      patterns[16394] = 29'b0_100000000001_010_1_000000000010;
      patterns[16395] = 29'b0_100000000001_011_0_000000000101;
      patterns[16396] = 29'b0_100000000001_100_1_010000000000;
      patterns[16397] = 29'b0_100000000001_101_0_101000000000;
      patterns[16398] = 29'b0_100000000001_110_0_100000000001;
      patterns[16399] = 29'b0_100000000001_111_0_100000000001;
      patterns[16400] = 29'b0_100000000010_000_0_100000000010;
      patterns[16401] = 29'b0_100000000010_001_0_000010100000;
      patterns[16402] = 29'b0_100000000010_010_1_000000000100;
      patterns[16403] = 29'b0_100000000010_011_0_000000001001;
      patterns[16404] = 29'b0_100000000010_100_0_010000000001;
      patterns[16405] = 29'b0_100000000010_101_1_001000000000;
      patterns[16406] = 29'b0_100000000010_110_0_100000000010;
      patterns[16407] = 29'b0_100000000010_111_0_100000000010;
      patterns[16408] = 29'b0_100000000011_000_0_100000000011;
      patterns[16409] = 29'b0_100000000011_001_0_000011100000;
      patterns[16410] = 29'b0_100000000011_010_1_000000000110;
      patterns[16411] = 29'b0_100000000011_011_0_000000001101;
      patterns[16412] = 29'b0_100000000011_100_1_010000000001;
      patterns[16413] = 29'b0_100000000011_101_1_101000000000;
      patterns[16414] = 29'b0_100000000011_110_0_100000000011;
      patterns[16415] = 29'b0_100000000011_111_0_100000000011;
      patterns[16416] = 29'b0_100000000100_000_0_100000000100;
      patterns[16417] = 29'b0_100000000100_001_0_000100100000;
      patterns[16418] = 29'b0_100000000100_010_1_000000001000;
      patterns[16419] = 29'b0_100000000100_011_0_000000010001;
      patterns[16420] = 29'b0_100000000100_100_0_010000000010;
      patterns[16421] = 29'b0_100000000100_101_0_001000000001;
      patterns[16422] = 29'b0_100000000100_110_0_100000000100;
      patterns[16423] = 29'b0_100000000100_111_0_100000000100;
      patterns[16424] = 29'b0_100000000101_000_0_100000000101;
      patterns[16425] = 29'b0_100000000101_001_0_000101100000;
      patterns[16426] = 29'b0_100000000101_010_1_000000001010;
      patterns[16427] = 29'b0_100000000101_011_0_000000010101;
      patterns[16428] = 29'b0_100000000101_100_1_010000000010;
      patterns[16429] = 29'b0_100000000101_101_0_101000000001;
      patterns[16430] = 29'b0_100000000101_110_0_100000000101;
      patterns[16431] = 29'b0_100000000101_111_0_100000000101;
      patterns[16432] = 29'b0_100000000110_000_0_100000000110;
      patterns[16433] = 29'b0_100000000110_001_0_000110100000;
      patterns[16434] = 29'b0_100000000110_010_1_000000001100;
      patterns[16435] = 29'b0_100000000110_011_0_000000011001;
      patterns[16436] = 29'b0_100000000110_100_0_010000000011;
      patterns[16437] = 29'b0_100000000110_101_1_001000000001;
      patterns[16438] = 29'b0_100000000110_110_0_100000000110;
      patterns[16439] = 29'b0_100000000110_111_0_100000000110;
      patterns[16440] = 29'b0_100000000111_000_0_100000000111;
      patterns[16441] = 29'b0_100000000111_001_0_000111100000;
      patterns[16442] = 29'b0_100000000111_010_1_000000001110;
      patterns[16443] = 29'b0_100000000111_011_0_000000011101;
      patterns[16444] = 29'b0_100000000111_100_1_010000000011;
      patterns[16445] = 29'b0_100000000111_101_1_101000000001;
      patterns[16446] = 29'b0_100000000111_110_0_100000000111;
      patterns[16447] = 29'b0_100000000111_111_0_100000000111;
      patterns[16448] = 29'b0_100000001000_000_0_100000001000;
      patterns[16449] = 29'b0_100000001000_001_0_001000100000;
      patterns[16450] = 29'b0_100000001000_010_1_000000010000;
      patterns[16451] = 29'b0_100000001000_011_0_000000100001;
      patterns[16452] = 29'b0_100000001000_100_0_010000000100;
      patterns[16453] = 29'b0_100000001000_101_0_001000000010;
      patterns[16454] = 29'b0_100000001000_110_0_100000001000;
      patterns[16455] = 29'b0_100000001000_111_0_100000001000;
      patterns[16456] = 29'b0_100000001001_000_0_100000001001;
      patterns[16457] = 29'b0_100000001001_001_0_001001100000;
      patterns[16458] = 29'b0_100000001001_010_1_000000010010;
      patterns[16459] = 29'b0_100000001001_011_0_000000100101;
      patterns[16460] = 29'b0_100000001001_100_1_010000000100;
      patterns[16461] = 29'b0_100000001001_101_0_101000000010;
      patterns[16462] = 29'b0_100000001001_110_0_100000001001;
      patterns[16463] = 29'b0_100000001001_111_0_100000001001;
      patterns[16464] = 29'b0_100000001010_000_0_100000001010;
      patterns[16465] = 29'b0_100000001010_001_0_001010100000;
      patterns[16466] = 29'b0_100000001010_010_1_000000010100;
      patterns[16467] = 29'b0_100000001010_011_0_000000101001;
      patterns[16468] = 29'b0_100000001010_100_0_010000000101;
      patterns[16469] = 29'b0_100000001010_101_1_001000000010;
      patterns[16470] = 29'b0_100000001010_110_0_100000001010;
      patterns[16471] = 29'b0_100000001010_111_0_100000001010;
      patterns[16472] = 29'b0_100000001011_000_0_100000001011;
      patterns[16473] = 29'b0_100000001011_001_0_001011100000;
      patterns[16474] = 29'b0_100000001011_010_1_000000010110;
      patterns[16475] = 29'b0_100000001011_011_0_000000101101;
      patterns[16476] = 29'b0_100000001011_100_1_010000000101;
      patterns[16477] = 29'b0_100000001011_101_1_101000000010;
      patterns[16478] = 29'b0_100000001011_110_0_100000001011;
      patterns[16479] = 29'b0_100000001011_111_0_100000001011;
      patterns[16480] = 29'b0_100000001100_000_0_100000001100;
      patterns[16481] = 29'b0_100000001100_001_0_001100100000;
      patterns[16482] = 29'b0_100000001100_010_1_000000011000;
      patterns[16483] = 29'b0_100000001100_011_0_000000110001;
      patterns[16484] = 29'b0_100000001100_100_0_010000000110;
      patterns[16485] = 29'b0_100000001100_101_0_001000000011;
      patterns[16486] = 29'b0_100000001100_110_0_100000001100;
      patterns[16487] = 29'b0_100000001100_111_0_100000001100;
      patterns[16488] = 29'b0_100000001101_000_0_100000001101;
      patterns[16489] = 29'b0_100000001101_001_0_001101100000;
      patterns[16490] = 29'b0_100000001101_010_1_000000011010;
      patterns[16491] = 29'b0_100000001101_011_0_000000110101;
      patterns[16492] = 29'b0_100000001101_100_1_010000000110;
      patterns[16493] = 29'b0_100000001101_101_0_101000000011;
      patterns[16494] = 29'b0_100000001101_110_0_100000001101;
      patterns[16495] = 29'b0_100000001101_111_0_100000001101;
      patterns[16496] = 29'b0_100000001110_000_0_100000001110;
      patterns[16497] = 29'b0_100000001110_001_0_001110100000;
      patterns[16498] = 29'b0_100000001110_010_1_000000011100;
      patterns[16499] = 29'b0_100000001110_011_0_000000111001;
      patterns[16500] = 29'b0_100000001110_100_0_010000000111;
      patterns[16501] = 29'b0_100000001110_101_1_001000000011;
      patterns[16502] = 29'b0_100000001110_110_0_100000001110;
      patterns[16503] = 29'b0_100000001110_111_0_100000001110;
      patterns[16504] = 29'b0_100000001111_000_0_100000001111;
      patterns[16505] = 29'b0_100000001111_001_0_001111100000;
      patterns[16506] = 29'b0_100000001111_010_1_000000011110;
      patterns[16507] = 29'b0_100000001111_011_0_000000111101;
      patterns[16508] = 29'b0_100000001111_100_1_010000000111;
      patterns[16509] = 29'b0_100000001111_101_1_101000000011;
      patterns[16510] = 29'b0_100000001111_110_0_100000001111;
      patterns[16511] = 29'b0_100000001111_111_0_100000001111;
      patterns[16512] = 29'b0_100000010000_000_0_100000010000;
      patterns[16513] = 29'b0_100000010000_001_0_010000100000;
      patterns[16514] = 29'b0_100000010000_010_1_000000100000;
      patterns[16515] = 29'b0_100000010000_011_0_000001000001;
      patterns[16516] = 29'b0_100000010000_100_0_010000001000;
      patterns[16517] = 29'b0_100000010000_101_0_001000000100;
      patterns[16518] = 29'b0_100000010000_110_0_100000010000;
      patterns[16519] = 29'b0_100000010000_111_0_100000010000;
      patterns[16520] = 29'b0_100000010001_000_0_100000010001;
      patterns[16521] = 29'b0_100000010001_001_0_010001100000;
      patterns[16522] = 29'b0_100000010001_010_1_000000100010;
      patterns[16523] = 29'b0_100000010001_011_0_000001000101;
      patterns[16524] = 29'b0_100000010001_100_1_010000001000;
      patterns[16525] = 29'b0_100000010001_101_0_101000000100;
      patterns[16526] = 29'b0_100000010001_110_0_100000010001;
      patterns[16527] = 29'b0_100000010001_111_0_100000010001;
      patterns[16528] = 29'b0_100000010010_000_0_100000010010;
      patterns[16529] = 29'b0_100000010010_001_0_010010100000;
      patterns[16530] = 29'b0_100000010010_010_1_000000100100;
      patterns[16531] = 29'b0_100000010010_011_0_000001001001;
      patterns[16532] = 29'b0_100000010010_100_0_010000001001;
      patterns[16533] = 29'b0_100000010010_101_1_001000000100;
      patterns[16534] = 29'b0_100000010010_110_0_100000010010;
      patterns[16535] = 29'b0_100000010010_111_0_100000010010;
      patterns[16536] = 29'b0_100000010011_000_0_100000010011;
      patterns[16537] = 29'b0_100000010011_001_0_010011100000;
      patterns[16538] = 29'b0_100000010011_010_1_000000100110;
      patterns[16539] = 29'b0_100000010011_011_0_000001001101;
      patterns[16540] = 29'b0_100000010011_100_1_010000001001;
      patterns[16541] = 29'b0_100000010011_101_1_101000000100;
      patterns[16542] = 29'b0_100000010011_110_0_100000010011;
      patterns[16543] = 29'b0_100000010011_111_0_100000010011;
      patterns[16544] = 29'b0_100000010100_000_0_100000010100;
      patterns[16545] = 29'b0_100000010100_001_0_010100100000;
      patterns[16546] = 29'b0_100000010100_010_1_000000101000;
      patterns[16547] = 29'b0_100000010100_011_0_000001010001;
      patterns[16548] = 29'b0_100000010100_100_0_010000001010;
      patterns[16549] = 29'b0_100000010100_101_0_001000000101;
      patterns[16550] = 29'b0_100000010100_110_0_100000010100;
      patterns[16551] = 29'b0_100000010100_111_0_100000010100;
      patterns[16552] = 29'b0_100000010101_000_0_100000010101;
      patterns[16553] = 29'b0_100000010101_001_0_010101100000;
      patterns[16554] = 29'b0_100000010101_010_1_000000101010;
      patterns[16555] = 29'b0_100000010101_011_0_000001010101;
      patterns[16556] = 29'b0_100000010101_100_1_010000001010;
      patterns[16557] = 29'b0_100000010101_101_0_101000000101;
      patterns[16558] = 29'b0_100000010101_110_0_100000010101;
      patterns[16559] = 29'b0_100000010101_111_0_100000010101;
      patterns[16560] = 29'b0_100000010110_000_0_100000010110;
      patterns[16561] = 29'b0_100000010110_001_0_010110100000;
      patterns[16562] = 29'b0_100000010110_010_1_000000101100;
      patterns[16563] = 29'b0_100000010110_011_0_000001011001;
      patterns[16564] = 29'b0_100000010110_100_0_010000001011;
      patterns[16565] = 29'b0_100000010110_101_1_001000000101;
      patterns[16566] = 29'b0_100000010110_110_0_100000010110;
      patterns[16567] = 29'b0_100000010110_111_0_100000010110;
      patterns[16568] = 29'b0_100000010111_000_0_100000010111;
      patterns[16569] = 29'b0_100000010111_001_0_010111100000;
      patterns[16570] = 29'b0_100000010111_010_1_000000101110;
      patterns[16571] = 29'b0_100000010111_011_0_000001011101;
      patterns[16572] = 29'b0_100000010111_100_1_010000001011;
      patterns[16573] = 29'b0_100000010111_101_1_101000000101;
      patterns[16574] = 29'b0_100000010111_110_0_100000010111;
      patterns[16575] = 29'b0_100000010111_111_0_100000010111;
      patterns[16576] = 29'b0_100000011000_000_0_100000011000;
      patterns[16577] = 29'b0_100000011000_001_0_011000100000;
      patterns[16578] = 29'b0_100000011000_010_1_000000110000;
      patterns[16579] = 29'b0_100000011000_011_0_000001100001;
      patterns[16580] = 29'b0_100000011000_100_0_010000001100;
      patterns[16581] = 29'b0_100000011000_101_0_001000000110;
      patterns[16582] = 29'b0_100000011000_110_0_100000011000;
      patterns[16583] = 29'b0_100000011000_111_0_100000011000;
      patterns[16584] = 29'b0_100000011001_000_0_100000011001;
      patterns[16585] = 29'b0_100000011001_001_0_011001100000;
      patterns[16586] = 29'b0_100000011001_010_1_000000110010;
      patterns[16587] = 29'b0_100000011001_011_0_000001100101;
      patterns[16588] = 29'b0_100000011001_100_1_010000001100;
      patterns[16589] = 29'b0_100000011001_101_0_101000000110;
      patterns[16590] = 29'b0_100000011001_110_0_100000011001;
      patterns[16591] = 29'b0_100000011001_111_0_100000011001;
      patterns[16592] = 29'b0_100000011010_000_0_100000011010;
      patterns[16593] = 29'b0_100000011010_001_0_011010100000;
      patterns[16594] = 29'b0_100000011010_010_1_000000110100;
      patterns[16595] = 29'b0_100000011010_011_0_000001101001;
      patterns[16596] = 29'b0_100000011010_100_0_010000001101;
      patterns[16597] = 29'b0_100000011010_101_1_001000000110;
      patterns[16598] = 29'b0_100000011010_110_0_100000011010;
      patterns[16599] = 29'b0_100000011010_111_0_100000011010;
      patterns[16600] = 29'b0_100000011011_000_0_100000011011;
      patterns[16601] = 29'b0_100000011011_001_0_011011100000;
      patterns[16602] = 29'b0_100000011011_010_1_000000110110;
      patterns[16603] = 29'b0_100000011011_011_0_000001101101;
      patterns[16604] = 29'b0_100000011011_100_1_010000001101;
      patterns[16605] = 29'b0_100000011011_101_1_101000000110;
      patterns[16606] = 29'b0_100000011011_110_0_100000011011;
      patterns[16607] = 29'b0_100000011011_111_0_100000011011;
      patterns[16608] = 29'b0_100000011100_000_0_100000011100;
      patterns[16609] = 29'b0_100000011100_001_0_011100100000;
      patterns[16610] = 29'b0_100000011100_010_1_000000111000;
      patterns[16611] = 29'b0_100000011100_011_0_000001110001;
      patterns[16612] = 29'b0_100000011100_100_0_010000001110;
      patterns[16613] = 29'b0_100000011100_101_0_001000000111;
      patterns[16614] = 29'b0_100000011100_110_0_100000011100;
      patterns[16615] = 29'b0_100000011100_111_0_100000011100;
      patterns[16616] = 29'b0_100000011101_000_0_100000011101;
      patterns[16617] = 29'b0_100000011101_001_0_011101100000;
      patterns[16618] = 29'b0_100000011101_010_1_000000111010;
      patterns[16619] = 29'b0_100000011101_011_0_000001110101;
      patterns[16620] = 29'b0_100000011101_100_1_010000001110;
      patterns[16621] = 29'b0_100000011101_101_0_101000000111;
      patterns[16622] = 29'b0_100000011101_110_0_100000011101;
      patterns[16623] = 29'b0_100000011101_111_0_100000011101;
      patterns[16624] = 29'b0_100000011110_000_0_100000011110;
      patterns[16625] = 29'b0_100000011110_001_0_011110100000;
      patterns[16626] = 29'b0_100000011110_010_1_000000111100;
      patterns[16627] = 29'b0_100000011110_011_0_000001111001;
      patterns[16628] = 29'b0_100000011110_100_0_010000001111;
      patterns[16629] = 29'b0_100000011110_101_1_001000000111;
      patterns[16630] = 29'b0_100000011110_110_0_100000011110;
      patterns[16631] = 29'b0_100000011110_111_0_100000011110;
      patterns[16632] = 29'b0_100000011111_000_0_100000011111;
      patterns[16633] = 29'b0_100000011111_001_0_011111100000;
      patterns[16634] = 29'b0_100000011111_010_1_000000111110;
      patterns[16635] = 29'b0_100000011111_011_0_000001111101;
      patterns[16636] = 29'b0_100000011111_100_1_010000001111;
      patterns[16637] = 29'b0_100000011111_101_1_101000000111;
      patterns[16638] = 29'b0_100000011111_110_0_100000011111;
      patterns[16639] = 29'b0_100000011111_111_0_100000011111;
      patterns[16640] = 29'b0_100000100000_000_0_100000100000;
      patterns[16641] = 29'b0_100000100000_001_0_100000100000;
      patterns[16642] = 29'b0_100000100000_010_1_000001000000;
      patterns[16643] = 29'b0_100000100000_011_0_000010000001;
      patterns[16644] = 29'b0_100000100000_100_0_010000010000;
      patterns[16645] = 29'b0_100000100000_101_0_001000001000;
      patterns[16646] = 29'b0_100000100000_110_0_100000100000;
      patterns[16647] = 29'b0_100000100000_111_0_100000100000;
      patterns[16648] = 29'b0_100000100001_000_0_100000100001;
      patterns[16649] = 29'b0_100000100001_001_0_100001100000;
      patterns[16650] = 29'b0_100000100001_010_1_000001000010;
      patterns[16651] = 29'b0_100000100001_011_0_000010000101;
      patterns[16652] = 29'b0_100000100001_100_1_010000010000;
      patterns[16653] = 29'b0_100000100001_101_0_101000001000;
      patterns[16654] = 29'b0_100000100001_110_0_100000100001;
      patterns[16655] = 29'b0_100000100001_111_0_100000100001;
      patterns[16656] = 29'b0_100000100010_000_0_100000100010;
      patterns[16657] = 29'b0_100000100010_001_0_100010100000;
      patterns[16658] = 29'b0_100000100010_010_1_000001000100;
      patterns[16659] = 29'b0_100000100010_011_0_000010001001;
      patterns[16660] = 29'b0_100000100010_100_0_010000010001;
      patterns[16661] = 29'b0_100000100010_101_1_001000001000;
      patterns[16662] = 29'b0_100000100010_110_0_100000100010;
      patterns[16663] = 29'b0_100000100010_111_0_100000100010;
      patterns[16664] = 29'b0_100000100011_000_0_100000100011;
      patterns[16665] = 29'b0_100000100011_001_0_100011100000;
      patterns[16666] = 29'b0_100000100011_010_1_000001000110;
      patterns[16667] = 29'b0_100000100011_011_0_000010001101;
      patterns[16668] = 29'b0_100000100011_100_1_010000010001;
      patterns[16669] = 29'b0_100000100011_101_1_101000001000;
      patterns[16670] = 29'b0_100000100011_110_0_100000100011;
      patterns[16671] = 29'b0_100000100011_111_0_100000100011;
      patterns[16672] = 29'b0_100000100100_000_0_100000100100;
      patterns[16673] = 29'b0_100000100100_001_0_100100100000;
      patterns[16674] = 29'b0_100000100100_010_1_000001001000;
      patterns[16675] = 29'b0_100000100100_011_0_000010010001;
      patterns[16676] = 29'b0_100000100100_100_0_010000010010;
      patterns[16677] = 29'b0_100000100100_101_0_001000001001;
      patterns[16678] = 29'b0_100000100100_110_0_100000100100;
      patterns[16679] = 29'b0_100000100100_111_0_100000100100;
      patterns[16680] = 29'b0_100000100101_000_0_100000100101;
      patterns[16681] = 29'b0_100000100101_001_0_100101100000;
      patterns[16682] = 29'b0_100000100101_010_1_000001001010;
      patterns[16683] = 29'b0_100000100101_011_0_000010010101;
      patterns[16684] = 29'b0_100000100101_100_1_010000010010;
      patterns[16685] = 29'b0_100000100101_101_0_101000001001;
      patterns[16686] = 29'b0_100000100101_110_0_100000100101;
      patterns[16687] = 29'b0_100000100101_111_0_100000100101;
      patterns[16688] = 29'b0_100000100110_000_0_100000100110;
      patterns[16689] = 29'b0_100000100110_001_0_100110100000;
      patterns[16690] = 29'b0_100000100110_010_1_000001001100;
      patterns[16691] = 29'b0_100000100110_011_0_000010011001;
      patterns[16692] = 29'b0_100000100110_100_0_010000010011;
      patterns[16693] = 29'b0_100000100110_101_1_001000001001;
      patterns[16694] = 29'b0_100000100110_110_0_100000100110;
      patterns[16695] = 29'b0_100000100110_111_0_100000100110;
      patterns[16696] = 29'b0_100000100111_000_0_100000100111;
      patterns[16697] = 29'b0_100000100111_001_0_100111100000;
      patterns[16698] = 29'b0_100000100111_010_1_000001001110;
      patterns[16699] = 29'b0_100000100111_011_0_000010011101;
      patterns[16700] = 29'b0_100000100111_100_1_010000010011;
      patterns[16701] = 29'b0_100000100111_101_1_101000001001;
      patterns[16702] = 29'b0_100000100111_110_0_100000100111;
      patterns[16703] = 29'b0_100000100111_111_0_100000100111;
      patterns[16704] = 29'b0_100000101000_000_0_100000101000;
      patterns[16705] = 29'b0_100000101000_001_0_101000100000;
      patterns[16706] = 29'b0_100000101000_010_1_000001010000;
      patterns[16707] = 29'b0_100000101000_011_0_000010100001;
      patterns[16708] = 29'b0_100000101000_100_0_010000010100;
      patterns[16709] = 29'b0_100000101000_101_0_001000001010;
      patterns[16710] = 29'b0_100000101000_110_0_100000101000;
      patterns[16711] = 29'b0_100000101000_111_0_100000101000;
      patterns[16712] = 29'b0_100000101001_000_0_100000101001;
      patterns[16713] = 29'b0_100000101001_001_0_101001100000;
      patterns[16714] = 29'b0_100000101001_010_1_000001010010;
      patterns[16715] = 29'b0_100000101001_011_0_000010100101;
      patterns[16716] = 29'b0_100000101001_100_1_010000010100;
      patterns[16717] = 29'b0_100000101001_101_0_101000001010;
      patterns[16718] = 29'b0_100000101001_110_0_100000101001;
      patterns[16719] = 29'b0_100000101001_111_0_100000101001;
      patterns[16720] = 29'b0_100000101010_000_0_100000101010;
      patterns[16721] = 29'b0_100000101010_001_0_101010100000;
      patterns[16722] = 29'b0_100000101010_010_1_000001010100;
      patterns[16723] = 29'b0_100000101010_011_0_000010101001;
      patterns[16724] = 29'b0_100000101010_100_0_010000010101;
      patterns[16725] = 29'b0_100000101010_101_1_001000001010;
      patterns[16726] = 29'b0_100000101010_110_0_100000101010;
      patterns[16727] = 29'b0_100000101010_111_0_100000101010;
      patterns[16728] = 29'b0_100000101011_000_0_100000101011;
      patterns[16729] = 29'b0_100000101011_001_0_101011100000;
      patterns[16730] = 29'b0_100000101011_010_1_000001010110;
      patterns[16731] = 29'b0_100000101011_011_0_000010101101;
      patterns[16732] = 29'b0_100000101011_100_1_010000010101;
      patterns[16733] = 29'b0_100000101011_101_1_101000001010;
      patterns[16734] = 29'b0_100000101011_110_0_100000101011;
      patterns[16735] = 29'b0_100000101011_111_0_100000101011;
      patterns[16736] = 29'b0_100000101100_000_0_100000101100;
      patterns[16737] = 29'b0_100000101100_001_0_101100100000;
      patterns[16738] = 29'b0_100000101100_010_1_000001011000;
      patterns[16739] = 29'b0_100000101100_011_0_000010110001;
      patterns[16740] = 29'b0_100000101100_100_0_010000010110;
      patterns[16741] = 29'b0_100000101100_101_0_001000001011;
      patterns[16742] = 29'b0_100000101100_110_0_100000101100;
      patterns[16743] = 29'b0_100000101100_111_0_100000101100;
      patterns[16744] = 29'b0_100000101101_000_0_100000101101;
      patterns[16745] = 29'b0_100000101101_001_0_101101100000;
      patterns[16746] = 29'b0_100000101101_010_1_000001011010;
      patterns[16747] = 29'b0_100000101101_011_0_000010110101;
      patterns[16748] = 29'b0_100000101101_100_1_010000010110;
      patterns[16749] = 29'b0_100000101101_101_0_101000001011;
      patterns[16750] = 29'b0_100000101101_110_0_100000101101;
      patterns[16751] = 29'b0_100000101101_111_0_100000101101;
      patterns[16752] = 29'b0_100000101110_000_0_100000101110;
      patterns[16753] = 29'b0_100000101110_001_0_101110100000;
      patterns[16754] = 29'b0_100000101110_010_1_000001011100;
      patterns[16755] = 29'b0_100000101110_011_0_000010111001;
      patterns[16756] = 29'b0_100000101110_100_0_010000010111;
      patterns[16757] = 29'b0_100000101110_101_1_001000001011;
      patterns[16758] = 29'b0_100000101110_110_0_100000101110;
      patterns[16759] = 29'b0_100000101110_111_0_100000101110;
      patterns[16760] = 29'b0_100000101111_000_0_100000101111;
      patterns[16761] = 29'b0_100000101111_001_0_101111100000;
      patterns[16762] = 29'b0_100000101111_010_1_000001011110;
      patterns[16763] = 29'b0_100000101111_011_0_000010111101;
      patterns[16764] = 29'b0_100000101111_100_1_010000010111;
      patterns[16765] = 29'b0_100000101111_101_1_101000001011;
      patterns[16766] = 29'b0_100000101111_110_0_100000101111;
      patterns[16767] = 29'b0_100000101111_111_0_100000101111;
      patterns[16768] = 29'b0_100000110000_000_0_100000110000;
      patterns[16769] = 29'b0_100000110000_001_0_110000100000;
      patterns[16770] = 29'b0_100000110000_010_1_000001100000;
      patterns[16771] = 29'b0_100000110000_011_0_000011000001;
      patterns[16772] = 29'b0_100000110000_100_0_010000011000;
      patterns[16773] = 29'b0_100000110000_101_0_001000001100;
      patterns[16774] = 29'b0_100000110000_110_0_100000110000;
      patterns[16775] = 29'b0_100000110000_111_0_100000110000;
      patterns[16776] = 29'b0_100000110001_000_0_100000110001;
      patterns[16777] = 29'b0_100000110001_001_0_110001100000;
      patterns[16778] = 29'b0_100000110001_010_1_000001100010;
      patterns[16779] = 29'b0_100000110001_011_0_000011000101;
      patterns[16780] = 29'b0_100000110001_100_1_010000011000;
      patterns[16781] = 29'b0_100000110001_101_0_101000001100;
      patterns[16782] = 29'b0_100000110001_110_0_100000110001;
      patterns[16783] = 29'b0_100000110001_111_0_100000110001;
      patterns[16784] = 29'b0_100000110010_000_0_100000110010;
      patterns[16785] = 29'b0_100000110010_001_0_110010100000;
      patterns[16786] = 29'b0_100000110010_010_1_000001100100;
      patterns[16787] = 29'b0_100000110010_011_0_000011001001;
      patterns[16788] = 29'b0_100000110010_100_0_010000011001;
      patterns[16789] = 29'b0_100000110010_101_1_001000001100;
      patterns[16790] = 29'b0_100000110010_110_0_100000110010;
      patterns[16791] = 29'b0_100000110010_111_0_100000110010;
      patterns[16792] = 29'b0_100000110011_000_0_100000110011;
      patterns[16793] = 29'b0_100000110011_001_0_110011100000;
      patterns[16794] = 29'b0_100000110011_010_1_000001100110;
      patterns[16795] = 29'b0_100000110011_011_0_000011001101;
      patterns[16796] = 29'b0_100000110011_100_1_010000011001;
      patterns[16797] = 29'b0_100000110011_101_1_101000001100;
      patterns[16798] = 29'b0_100000110011_110_0_100000110011;
      patterns[16799] = 29'b0_100000110011_111_0_100000110011;
      patterns[16800] = 29'b0_100000110100_000_0_100000110100;
      patterns[16801] = 29'b0_100000110100_001_0_110100100000;
      patterns[16802] = 29'b0_100000110100_010_1_000001101000;
      patterns[16803] = 29'b0_100000110100_011_0_000011010001;
      patterns[16804] = 29'b0_100000110100_100_0_010000011010;
      patterns[16805] = 29'b0_100000110100_101_0_001000001101;
      patterns[16806] = 29'b0_100000110100_110_0_100000110100;
      patterns[16807] = 29'b0_100000110100_111_0_100000110100;
      patterns[16808] = 29'b0_100000110101_000_0_100000110101;
      patterns[16809] = 29'b0_100000110101_001_0_110101100000;
      patterns[16810] = 29'b0_100000110101_010_1_000001101010;
      patterns[16811] = 29'b0_100000110101_011_0_000011010101;
      patterns[16812] = 29'b0_100000110101_100_1_010000011010;
      patterns[16813] = 29'b0_100000110101_101_0_101000001101;
      patterns[16814] = 29'b0_100000110101_110_0_100000110101;
      patterns[16815] = 29'b0_100000110101_111_0_100000110101;
      patterns[16816] = 29'b0_100000110110_000_0_100000110110;
      patterns[16817] = 29'b0_100000110110_001_0_110110100000;
      patterns[16818] = 29'b0_100000110110_010_1_000001101100;
      patterns[16819] = 29'b0_100000110110_011_0_000011011001;
      patterns[16820] = 29'b0_100000110110_100_0_010000011011;
      patterns[16821] = 29'b0_100000110110_101_1_001000001101;
      patterns[16822] = 29'b0_100000110110_110_0_100000110110;
      patterns[16823] = 29'b0_100000110110_111_0_100000110110;
      patterns[16824] = 29'b0_100000110111_000_0_100000110111;
      patterns[16825] = 29'b0_100000110111_001_0_110111100000;
      patterns[16826] = 29'b0_100000110111_010_1_000001101110;
      patterns[16827] = 29'b0_100000110111_011_0_000011011101;
      patterns[16828] = 29'b0_100000110111_100_1_010000011011;
      patterns[16829] = 29'b0_100000110111_101_1_101000001101;
      patterns[16830] = 29'b0_100000110111_110_0_100000110111;
      patterns[16831] = 29'b0_100000110111_111_0_100000110111;
      patterns[16832] = 29'b0_100000111000_000_0_100000111000;
      patterns[16833] = 29'b0_100000111000_001_0_111000100000;
      patterns[16834] = 29'b0_100000111000_010_1_000001110000;
      patterns[16835] = 29'b0_100000111000_011_0_000011100001;
      patterns[16836] = 29'b0_100000111000_100_0_010000011100;
      patterns[16837] = 29'b0_100000111000_101_0_001000001110;
      patterns[16838] = 29'b0_100000111000_110_0_100000111000;
      patterns[16839] = 29'b0_100000111000_111_0_100000111000;
      patterns[16840] = 29'b0_100000111001_000_0_100000111001;
      patterns[16841] = 29'b0_100000111001_001_0_111001100000;
      patterns[16842] = 29'b0_100000111001_010_1_000001110010;
      patterns[16843] = 29'b0_100000111001_011_0_000011100101;
      patterns[16844] = 29'b0_100000111001_100_1_010000011100;
      patterns[16845] = 29'b0_100000111001_101_0_101000001110;
      patterns[16846] = 29'b0_100000111001_110_0_100000111001;
      patterns[16847] = 29'b0_100000111001_111_0_100000111001;
      patterns[16848] = 29'b0_100000111010_000_0_100000111010;
      patterns[16849] = 29'b0_100000111010_001_0_111010100000;
      patterns[16850] = 29'b0_100000111010_010_1_000001110100;
      patterns[16851] = 29'b0_100000111010_011_0_000011101001;
      patterns[16852] = 29'b0_100000111010_100_0_010000011101;
      patterns[16853] = 29'b0_100000111010_101_1_001000001110;
      patterns[16854] = 29'b0_100000111010_110_0_100000111010;
      patterns[16855] = 29'b0_100000111010_111_0_100000111010;
      patterns[16856] = 29'b0_100000111011_000_0_100000111011;
      patterns[16857] = 29'b0_100000111011_001_0_111011100000;
      patterns[16858] = 29'b0_100000111011_010_1_000001110110;
      patterns[16859] = 29'b0_100000111011_011_0_000011101101;
      patterns[16860] = 29'b0_100000111011_100_1_010000011101;
      patterns[16861] = 29'b0_100000111011_101_1_101000001110;
      patterns[16862] = 29'b0_100000111011_110_0_100000111011;
      patterns[16863] = 29'b0_100000111011_111_0_100000111011;
      patterns[16864] = 29'b0_100000111100_000_0_100000111100;
      patterns[16865] = 29'b0_100000111100_001_0_111100100000;
      patterns[16866] = 29'b0_100000111100_010_1_000001111000;
      patterns[16867] = 29'b0_100000111100_011_0_000011110001;
      patterns[16868] = 29'b0_100000111100_100_0_010000011110;
      patterns[16869] = 29'b0_100000111100_101_0_001000001111;
      patterns[16870] = 29'b0_100000111100_110_0_100000111100;
      patterns[16871] = 29'b0_100000111100_111_0_100000111100;
      patterns[16872] = 29'b0_100000111101_000_0_100000111101;
      patterns[16873] = 29'b0_100000111101_001_0_111101100000;
      patterns[16874] = 29'b0_100000111101_010_1_000001111010;
      patterns[16875] = 29'b0_100000111101_011_0_000011110101;
      patterns[16876] = 29'b0_100000111101_100_1_010000011110;
      patterns[16877] = 29'b0_100000111101_101_0_101000001111;
      patterns[16878] = 29'b0_100000111101_110_0_100000111101;
      patterns[16879] = 29'b0_100000111101_111_0_100000111101;
      patterns[16880] = 29'b0_100000111110_000_0_100000111110;
      patterns[16881] = 29'b0_100000111110_001_0_111110100000;
      patterns[16882] = 29'b0_100000111110_010_1_000001111100;
      patterns[16883] = 29'b0_100000111110_011_0_000011111001;
      patterns[16884] = 29'b0_100000111110_100_0_010000011111;
      patterns[16885] = 29'b0_100000111110_101_1_001000001111;
      patterns[16886] = 29'b0_100000111110_110_0_100000111110;
      patterns[16887] = 29'b0_100000111110_111_0_100000111110;
      patterns[16888] = 29'b0_100000111111_000_0_100000111111;
      patterns[16889] = 29'b0_100000111111_001_0_111111100000;
      patterns[16890] = 29'b0_100000111111_010_1_000001111110;
      patterns[16891] = 29'b0_100000111111_011_0_000011111101;
      patterns[16892] = 29'b0_100000111111_100_1_010000011111;
      patterns[16893] = 29'b0_100000111111_101_1_101000001111;
      patterns[16894] = 29'b0_100000111111_110_0_100000111111;
      patterns[16895] = 29'b0_100000111111_111_0_100000111111;
      patterns[16896] = 29'b0_100001000000_000_0_100001000000;
      patterns[16897] = 29'b0_100001000000_001_0_000000100001;
      patterns[16898] = 29'b0_100001000000_010_1_000010000000;
      patterns[16899] = 29'b0_100001000000_011_0_000100000001;
      patterns[16900] = 29'b0_100001000000_100_0_010000100000;
      patterns[16901] = 29'b0_100001000000_101_0_001000010000;
      patterns[16902] = 29'b0_100001000000_110_0_100001000000;
      patterns[16903] = 29'b0_100001000000_111_0_100001000000;
      patterns[16904] = 29'b0_100001000001_000_0_100001000001;
      patterns[16905] = 29'b0_100001000001_001_0_000001100001;
      patterns[16906] = 29'b0_100001000001_010_1_000010000010;
      patterns[16907] = 29'b0_100001000001_011_0_000100000101;
      patterns[16908] = 29'b0_100001000001_100_1_010000100000;
      patterns[16909] = 29'b0_100001000001_101_0_101000010000;
      patterns[16910] = 29'b0_100001000001_110_0_100001000001;
      patterns[16911] = 29'b0_100001000001_111_0_100001000001;
      patterns[16912] = 29'b0_100001000010_000_0_100001000010;
      patterns[16913] = 29'b0_100001000010_001_0_000010100001;
      patterns[16914] = 29'b0_100001000010_010_1_000010000100;
      patterns[16915] = 29'b0_100001000010_011_0_000100001001;
      patterns[16916] = 29'b0_100001000010_100_0_010000100001;
      patterns[16917] = 29'b0_100001000010_101_1_001000010000;
      patterns[16918] = 29'b0_100001000010_110_0_100001000010;
      patterns[16919] = 29'b0_100001000010_111_0_100001000010;
      patterns[16920] = 29'b0_100001000011_000_0_100001000011;
      patterns[16921] = 29'b0_100001000011_001_0_000011100001;
      patterns[16922] = 29'b0_100001000011_010_1_000010000110;
      patterns[16923] = 29'b0_100001000011_011_0_000100001101;
      patterns[16924] = 29'b0_100001000011_100_1_010000100001;
      patterns[16925] = 29'b0_100001000011_101_1_101000010000;
      patterns[16926] = 29'b0_100001000011_110_0_100001000011;
      patterns[16927] = 29'b0_100001000011_111_0_100001000011;
      patterns[16928] = 29'b0_100001000100_000_0_100001000100;
      patterns[16929] = 29'b0_100001000100_001_0_000100100001;
      patterns[16930] = 29'b0_100001000100_010_1_000010001000;
      patterns[16931] = 29'b0_100001000100_011_0_000100010001;
      patterns[16932] = 29'b0_100001000100_100_0_010000100010;
      patterns[16933] = 29'b0_100001000100_101_0_001000010001;
      patterns[16934] = 29'b0_100001000100_110_0_100001000100;
      patterns[16935] = 29'b0_100001000100_111_0_100001000100;
      patterns[16936] = 29'b0_100001000101_000_0_100001000101;
      patterns[16937] = 29'b0_100001000101_001_0_000101100001;
      patterns[16938] = 29'b0_100001000101_010_1_000010001010;
      patterns[16939] = 29'b0_100001000101_011_0_000100010101;
      patterns[16940] = 29'b0_100001000101_100_1_010000100010;
      patterns[16941] = 29'b0_100001000101_101_0_101000010001;
      patterns[16942] = 29'b0_100001000101_110_0_100001000101;
      patterns[16943] = 29'b0_100001000101_111_0_100001000101;
      patterns[16944] = 29'b0_100001000110_000_0_100001000110;
      patterns[16945] = 29'b0_100001000110_001_0_000110100001;
      patterns[16946] = 29'b0_100001000110_010_1_000010001100;
      patterns[16947] = 29'b0_100001000110_011_0_000100011001;
      patterns[16948] = 29'b0_100001000110_100_0_010000100011;
      patterns[16949] = 29'b0_100001000110_101_1_001000010001;
      patterns[16950] = 29'b0_100001000110_110_0_100001000110;
      patterns[16951] = 29'b0_100001000110_111_0_100001000110;
      patterns[16952] = 29'b0_100001000111_000_0_100001000111;
      patterns[16953] = 29'b0_100001000111_001_0_000111100001;
      patterns[16954] = 29'b0_100001000111_010_1_000010001110;
      patterns[16955] = 29'b0_100001000111_011_0_000100011101;
      patterns[16956] = 29'b0_100001000111_100_1_010000100011;
      patterns[16957] = 29'b0_100001000111_101_1_101000010001;
      patterns[16958] = 29'b0_100001000111_110_0_100001000111;
      patterns[16959] = 29'b0_100001000111_111_0_100001000111;
      patterns[16960] = 29'b0_100001001000_000_0_100001001000;
      patterns[16961] = 29'b0_100001001000_001_0_001000100001;
      patterns[16962] = 29'b0_100001001000_010_1_000010010000;
      patterns[16963] = 29'b0_100001001000_011_0_000100100001;
      patterns[16964] = 29'b0_100001001000_100_0_010000100100;
      patterns[16965] = 29'b0_100001001000_101_0_001000010010;
      patterns[16966] = 29'b0_100001001000_110_0_100001001000;
      patterns[16967] = 29'b0_100001001000_111_0_100001001000;
      patterns[16968] = 29'b0_100001001001_000_0_100001001001;
      patterns[16969] = 29'b0_100001001001_001_0_001001100001;
      patterns[16970] = 29'b0_100001001001_010_1_000010010010;
      patterns[16971] = 29'b0_100001001001_011_0_000100100101;
      patterns[16972] = 29'b0_100001001001_100_1_010000100100;
      patterns[16973] = 29'b0_100001001001_101_0_101000010010;
      patterns[16974] = 29'b0_100001001001_110_0_100001001001;
      patterns[16975] = 29'b0_100001001001_111_0_100001001001;
      patterns[16976] = 29'b0_100001001010_000_0_100001001010;
      patterns[16977] = 29'b0_100001001010_001_0_001010100001;
      patterns[16978] = 29'b0_100001001010_010_1_000010010100;
      patterns[16979] = 29'b0_100001001010_011_0_000100101001;
      patterns[16980] = 29'b0_100001001010_100_0_010000100101;
      patterns[16981] = 29'b0_100001001010_101_1_001000010010;
      patterns[16982] = 29'b0_100001001010_110_0_100001001010;
      patterns[16983] = 29'b0_100001001010_111_0_100001001010;
      patterns[16984] = 29'b0_100001001011_000_0_100001001011;
      patterns[16985] = 29'b0_100001001011_001_0_001011100001;
      patterns[16986] = 29'b0_100001001011_010_1_000010010110;
      patterns[16987] = 29'b0_100001001011_011_0_000100101101;
      patterns[16988] = 29'b0_100001001011_100_1_010000100101;
      patterns[16989] = 29'b0_100001001011_101_1_101000010010;
      patterns[16990] = 29'b0_100001001011_110_0_100001001011;
      patterns[16991] = 29'b0_100001001011_111_0_100001001011;
      patterns[16992] = 29'b0_100001001100_000_0_100001001100;
      patterns[16993] = 29'b0_100001001100_001_0_001100100001;
      patterns[16994] = 29'b0_100001001100_010_1_000010011000;
      patterns[16995] = 29'b0_100001001100_011_0_000100110001;
      patterns[16996] = 29'b0_100001001100_100_0_010000100110;
      patterns[16997] = 29'b0_100001001100_101_0_001000010011;
      patterns[16998] = 29'b0_100001001100_110_0_100001001100;
      patterns[16999] = 29'b0_100001001100_111_0_100001001100;
      patterns[17000] = 29'b0_100001001101_000_0_100001001101;
      patterns[17001] = 29'b0_100001001101_001_0_001101100001;
      patterns[17002] = 29'b0_100001001101_010_1_000010011010;
      patterns[17003] = 29'b0_100001001101_011_0_000100110101;
      patterns[17004] = 29'b0_100001001101_100_1_010000100110;
      patterns[17005] = 29'b0_100001001101_101_0_101000010011;
      patterns[17006] = 29'b0_100001001101_110_0_100001001101;
      patterns[17007] = 29'b0_100001001101_111_0_100001001101;
      patterns[17008] = 29'b0_100001001110_000_0_100001001110;
      patterns[17009] = 29'b0_100001001110_001_0_001110100001;
      patterns[17010] = 29'b0_100001001110_010_1_000010011100;
      patterns[17011] = 29'b0_100001001110_011_0_000100111001;
      patterns[17012] = 29'b0_100001001110_100_0_010000100111;
      patterns[17013] = 29'b0_100001001110_101_1_001000010011;
      patterns[17014] = 29'b0_100001001110_110_0_100001001110;
      patterns[17015] = 29'b0_100001001110_111_0_100001001110;
      patterns[17016] = 29'b0_100001001111_000_0_100001001111;
      patterns[17017] = 29'b0_100001001111_001_0_001111100001;
      patterns[17018] = 29'b0_100001001111_010_1_000010011110;
      patterns[17019] = 29'b0_100001001111_011_0_000100111101;
      patterns[17020] = 29'b0_100001001111_100_1_010000100111;
      patterns[17021] = 29'b0_100001001111_101_1_101000010011;
      patterns[17022] = 29'b0_100001001111_110_0_100001001111;
      patterns[17023] = 29'b0_100001001111_111_0_100001001111;
      patterns[17024] = 29'b0_100001010000_000_0_100001010000;
      patterns[17025] = 29'b0_100001010000_001_0_010000100001;
      patterns[17026] = 29'b0_100001010000_010_1_000010100000;
      patterns[17027] = 29'b0_100001010000_011_0_000101000001;
      patterns[17028] = 29'b0_100001010000_100_0_010000101000;
      patterns[17029] = 29'b0_100001010000_101_0_001000010100;
      patterns[17030] = 29'b0_100001010000_110_0_100001010000;
      patterns[17031] = 29'b0_100001010000_111_0_100001010000;
      patterns[17032] = 29'b0_100001010001_000_0_100001010001;
      patterns[17033] = 29'b0_100001010001_001_0_010001100001;
      patterns[17034] = 29'b0_100001010001_010_1_000010100010;
      patterns[17035] = 29'b0_100001010001_011_0_000101000101;
      patterns[17036] = 29'b0_100001010001_100_1_010000101000;
      patterns[17037] = 29'b0_100001010001_101_0_101000010100;
      patterns[17038] = 29'b0_100001010001_110_0_100001010001;
      patterns[17039] = 29'b0_100001010001_111_0_100001010001;
      patterns[17040] = 29'b0_100001010010_000_0_100001010010;
      patterns[17041] = 29'b0_100001010010_001_0_010010100001;
      patterns[17042] = 29'b0_100001010010_010_1_000010100100;
      patterns[17043] = 29'b0_100001010010_011_0_000101001001;
      patterns[17044] = 29'b0_100001010010_100_0_010000101001;
      patterns[17045] = 29'b0_100001010010_101_1_001000010100;
      patterns[17046] = 29'b0_100001010010_110_0_100001010010;
      patterns[17047] = 29'b0_100001010010_111_0_100001010010;
      patterns[17048] = 29'b0_100001010011_000_0_100001010011;
      patterns[17049] = 29'b0_100001010011_001_0_010011100001;
      patterns[17050] = 29'b0_100001010011_010_1_000010100110;
      patterns[17051] = 29'b0_100001010011_011_0_000101001101;
      patterns[17052] = 29'b0_100001010011_100_1_010000101001;
      patterns[17053] = 29'b0_100001010011_101_1_101000010100;
      patterns[17054] = 29'b0_100001010011_110_0_100001010011;
      patterns[17055] = 29'b0_100001010011_111_0_100001010011;
      patterns[17056] = 29'b0_100001010100_000_0_100001010100;
      patterns[17057] = 29'b0_100001010100_001_0_010100100001;
      patterns[17058] = 29'b0_100001010100_010_1_000010101000;
      patterns[17059] = 29'b0_100001010100_011_0_000101010001;
      patterns[17060] = 29'b0_100001010100_100_0_010000101010;
      patterns[17061] = 29'b0_100001010100_101_0_001000010101;
      patterns[17062] = 29'b0_100001010100_110_0_100001010100;
      patterns[17063] = 29'b0_100001010100_111_0_100001010100;
      patterns[17064] = 29'b0_100001010101_000_0_100001010101;
      patterns[17065] = 29'b0_100001010101_001_0_010101100001;
      patterns[17066] = 29'b0_100001010101_010_1_000010101010;
      patterns[17067] = 29'b0_100001010101_011_0_000101010101;
      patterns[17068] = 29'b0_100001010101_100_1_010000101010;
      patterns[17069] = 29'b0_100001010101_101_0_101000010101;
      patterns[17070] = 29'b0_100001010101_110_0_100001010101;
      patterns[17071] = 29'b0_100001010101_111_0_100001010101;
      patterns[17072] = 29'b0_100001010110_000_0_100001010110;
      patterns[17073] = 29'b0_100001010110_001_0_010110100001;
      patterns[17074] = 29'b0_100001010110_010_1_000010101100;
      patterns[17075] = 29'b0_100001010110_011_0_000101011001;
      patterns[17076] = 29'b0_100001010110_100_0_010000101011;
      patterns[17077] = 29'b0_100001010110_101_1_001000010101;
      patterns[17078] = 29'b0_100001010110_110_0_100001010110;
      patterns[17079] = 29'b0_100001010110_111_0_100001010110;
      patterns[17080] = 29'b0_100001010111_000_0_100001010111;
      patterns[17081] = 29'b0_100001010111_001_0_010111100001;
      patterns[17082] = 29'b0_100001010111_010_1_000010101110;
      patterns[17083] = 29'b0_100001010111_011_0_000101011101;
      patterns[17084] = 29'b0_100001010111_100_1_010000101011;
      patterns[17085] = 29'b0_100001010111_101_1_101000010101;
      patterns[17086] = 29'b0_100001010111_110_0_100001010111;
      patterns[17087] = 29'b0_100001010111_111_0_100001010111;
      patterns[17088] = 29'b0_100001011000_000_0_100001011000;
      patterns[17089] = 29'b0_100001011000_001_0_011000100001;
      patterns[17090] = 29'b0_100001011000_010_1_000010110000;
      patterns[17091] = 29'b0_100001011000_011_0_000101100001;
      patterns[17092] = 29'b0_100001011000_100_0_010000101100;
      patterns[17093] = 29'b0_100001011000_101_0_001000010110;
      patterns[17094] = 29'b0_100001011000_110_0_100001011000;
      patterns[17095] = 29'b0_100001011000_111_0_100001011000;
      patterns[17096] = 29'b0_100001011001_000_0_100001011001;
      patterns[17097] = 29'b0_100001011001_001_0_011001100001;
      patterns[17098] = 29'b0_100001011001_010_1_000010110010;
      patterns[17099] = 29'b0_100001011001_011_0_000101100101;
      patterns[17100] = 29'b0_100001011001_100_1_010000101100;
      patterns[17101] = 29'b0_100001011001_101_0_101000010110;
      patterns[17102] = 29'b0_100001011001_110_0_100001011001;
      patterns[17103] = 29'b0_100001011001_111_0_100001011001;
      patterns[17104] = 29'b0_100001011010_000_0_100001011010;
      patterns[17105] = 29'b0_100001011010_001_0_011010100001;
      patterns[17106] = 29'b0_100001011010_010_1_000010110100;
      patterns[17107] = 29'b0_100001011010_011_0_000101101001;
      patterns[17108] = 29'b0_100001011010_100_0_010000101101;
      patterns[17109] = 29'b0_100001011010_101_1_001000010110;
      patterns[17110] = 29'b0_100001011010_110_0_100001011010;
      patterns[17111] = 29'b0_100001011010_111_0_100001011010;
      patterns[17112] = 29'b0_100001011011_000_0_100001011011;
      patterns[17113] = 29'b0_100001011011_001_0_011011100001;
      patterns[17114] = 29'b0_100001011011_010_1_000010110110;
      patterns[17115] = 29'b0_100001011011_011_0_000101101101;
      patterns[17116] = 29'b0_100001011011_100_1_010000101101;
      patterns[17117] = 29'b0_100001011011_101_1_101000010110;
      patterns[17118] = 29'b0_100001011011_110_0_100001011011;
      patterns[17119] = 29'b0_100001011011_111_0_100001011011;
      patterns[17120] = 29'b0_100001011100_000_0_100001011100;
      patterns[17121] = 29'b0_100001011100_001_0_011100100001;
      patterns[17122] = 29'b0_100001011100_010_1_000010111000;
      patterns[17123] = 29'b0_100001011100_011_0_000101110001;
      patterns[17124] = 29'b0_100001011100_100_0_010000101110;
      patterns[17125] = 29'b0_100001011100_101_0_001000010111;
      patterns[17126] = 29'b0_100001011100_110_0_100001011100;
      patterns[17127] = 29'b0_100001011100_111_0_100001011100;
      patterns[17128] = 29'b0_100001011101_000_0_100001011101;
      patterns[17129] = 29'b0_100001011101_001_0_011101100001;
      patterns[17130] = 29'b0_100001011101_010_1_000010111010;
      patterns[17131] = 29'b0_100001011101_011_0_000101110101;
      patterns[17132] = 29'b0_100001011101_100_1_010000101110;
      patterns[17133] = 29'b0_100001011101_101_0_101000010111;
      patterns[17134] = 29'b0_100001011101_110_0_100001011101;
      patterns[17135] = 29'b0_100001011101_111_0_100001011101;
      patterns[17136] = 29'b0_100001011110_000_0_100001011110;
      patterns[17137] = 29'b0_100001011110_001_0_011110100001;
      patterns[17138] = 29'b0_100001011110_010_1_000010111100;
      patterns[17139] = 29'b0_100001011110_011_0_000101111001;
      patterns[17140] = 29'b0_100001011110_100_0_010000101111;
      patterns[17141] = 29'b0_100001011110_101_1_001000010111;
      patterns[17142] = 29'b0_100001011110_110_0_100001011110;
      patterns[17143] = 29'b0_100001011110_111_0_100001011110;
      patterns[17144] = 29'b0_100001011111_000_0_100001011111;
      patterns[17145] = 29'b0_100001011111_001_0_011111100001;
      patterns[17146] = 29'b0_100001011111_010_1_000010111110;
      patterns[17147] = 29'b0_100001011111_011_0_000101111101;
      patterns[17148] = 29'b0_100001011111_100_1_010000101111;
      patterns[17149] = 29'b0_100001011111_101_1_101000010111;
      patterns[17150] = 29'b0_100001011111_110_0_100001011111;
      patterns[17151] = 29'b0_100001011111_111_0_100001011111;
      patterns[17152] = 29'b0_100001100000_000_0_100001100000;
      patterns[17153] = 29'b0_100001100000_001_0_100000100001;
      patterns[17154] = 29'b0_100001100000_010_1_000011000000;
      patterns[17155] = 29'b0_100001100000_011_0_000110000001;
      patterns[17156] = 29'b0_100001100000_100_0_010000110000;
      patterns[17157] = 29'b0_100001100000_101_0_001000011000;
      patterns[17158] = 29'b0_100001100000_110_0_100001100000;
      patterns[17159] = 29'b0_100001100000_111_0_100001100000;
      patterns[17160] = 29'b0_100001100001_000_0_100001100001;
      patterns[17161] = 29'b0_100001100001_001_0_100001100001;
      patterns[17162] = 29'b0_100001100001_010_1_000011000010;
      patterns[17163] = 29'b0_100001100001_011_0_000110000101;
      patterns[17164] = 29'b0_100001100001_100_1_010000110000;
      patterns[17165] = 29'b0_100001100001_101_0_101000011000;
      patterns[17166] = 29'b0_100001100001_110_0_100001100001;
      patterns[17167] = 29'b0_100001100001_111_0_100001100001;
      patterns[17168] = 29'b0_100001100010_000_0_100001100010;
      patterns[17169] = 29'b0_100001100010_001_0_100010100001;
      patterns[17170] = 29'b0_100001100010_010_1_000011000100;
      patterns[17171] = 29'b0_100001100010_011_0_000110001001;
      patterns[17172] = 29'b0_100001100010_100_0_010000110001;
      patterns[17173] = 29'b0_100001100010_101_1_001000011000;
      patterns[17174] = 29'b0_100001100010_110_0_100001100010;
      patterns[17175] = 29'b0_100001100010_111_0_100001100010;
      patterns[17176] = 29'b0_100001100011_000_0_100001100011;
      patterns[17177] = 29'b0_100001100011_001_0_100011100001;
      patterns[17178] = 29'b0_100001100011_010_1_000011000110;
      patterns[17179] = 29'b0_100001100011_011_0_000110001101;
      patterns[17180] = 29'b0_100001100011_100_1_010000110001;
      patterns[17181] = 29'b0_100001100011_101_1_101000011000;
      patterns[17182] = 29'b0_100001100011_110_0_100001100011;
      patterns[17183] = 29'b0_100001100011_111_0_100001100011;
      patterns[17184] = 29'b0_100001100100_000_0_100001100100;
      patterns[17185] = 29'b0_100001100100_001_0_100100100001;
      patterns[17186] = 29'b0_100001100100_010_1_000011001000;
      patterns[17187] = 29'b0_100001100100_011_0_000110010001;
      patterns[17188] = 29'b0_100001100100_100_0_010000110010;
      patterns[17189] = 29'b0_100001100100_101_0_001000011001;
      patterns[17190] = 29'b0_100001100100_110_0_100001100100;
      patterns[17191] = 29'b0_100001100100_111_0_100001100100;
      patterns[17192] = 29'b0_100001100101_000_0_100001100101;
      patterns[17193] = 29'b0_100001100101_001_0_100101100001;
      patterns[17194] = 29'b0_100001100101_010_1_000011001010;
      patterns[17195] = 29'b0_100001100101_011_0_000110010101;
      patterns[17196] = 29'b0_100001100101_100_1_010000110010;
      patterns[17197] = 29'b0_100001100101_101_0_101000011001;
      patterns[17198] = 29'b0_100001100101_110_0_100001100101;
      patterns[17199] = 29'b0_100001100101_111_0_100001100101;
      patterns[17200] = 29'b0_100001100110_000_0_100001100110;
      patterns[17201] = 29'b0_100001100110_001_0_100110100001;
      patterns[17202] = 29'b0_100001100110_010_1_000011001100;
      patterns[17203] = 29'b0_100001100110_011_0_000110011001;
      patterns[17204] = 29'b0_100001100110_100_0_010000110011;
      patterns[17205] = 29'b0_100001100110_101_1_001000011001;
      patterns[17206] = 29'b0_100001100110_110_0_100001100110;
      patterns[17207] = 29'b0_100001100110_111_0_100001100110;
      patterns[17208] = 29'b0_100001100111_000_0_100001100111;
      patterns[17209] = 29'b0_100001100111_001_0_100111100001;
      patterns[17210] = 29'b0_100001100111_010_1_000011001110;
      patterns[17211] = 29'b0_100001100111_011_0_000110011101;
      patterns[17212] = 29'b0_100001100111_100_1_010000110011;
      patterns[17213] = 29'b0_100001100111_101_1_101000011001;
      patterns[17214] = 29'b0_100001100111_110_0_100001100111;
      patterns[17215] = 29'b0_100001100111_111_0_100001100111;
      patterns[17216] = 29'b0_100001101000_000_0_100001101000;
      patterns[17217] = 29'b0_100001101000_001_0_101000100001;
      patterns[17218] = 29'b0_100001101000_010_1_000011010000;
      patterns[17219] = 29'b0_100001101000_011_0_000110100001;
      patterns[17220] = 29'b0_100001101000_100_0_010000110100;
      patterns[17221] = 29'b0_100001101000_101_0_001000011010;
      patterns[17222] = 29'b0_100001101000_110_0_100001101000;
      patterns[17223] = 29'b0_100001101000_111_0_100001101000;
      patterns[17224] = 29'b0_100001101001_000_0_100001101001;
      patterns[17225] = 29'b0_100001101001_001_0_101001100001;
      patterns[17226] = 29'b0_100001101001_010_1_000011010010;
      patterns[17227] = 29'b0_100001101001_011_0_000110100101;
      patterns[17228] = 29'b0_100001101001_100_1_010000110100;
      patterns[17229] = 29'b0_100001101001_101_0_101000011010;
      patterns[17230] = 29'b0_100001101001_110_0_100001101001;
      patterns[17231] = 29'b0_100001101001_111_0_100001101001;
      patterns[17232] = 29'b0_100001101010_000_0_100001101010;
      patterns[17233] = 29'b0_100001101010_001_0_101010100001;
      patterns[17234] = 29'b0_100001101010_010_1_000011010100;
      patterns[17235] = 29'b0_100001101010_011_0_000110101001;
      patterns[17236] = 29'b0_100001101010_100_0_010000110101;
      patterns[17237] = 29'b0_100001101010_101_1_001000011010;
      patterns[17238] = 29'b0_100001101010_110_0_100001101010;
      patterns[17239] = 29'b0_100001101010_111_0_100001101010;
      patterns[17240] = 29'b0_100001101011_000_0_100001101011;
      patterns[17241] = 29'b0_100001101011_001_0_101011100001;
      patterns[17242] = 29'b0_100001101011_010_1_000011010110;
      patterns[17243] = 29'b0_100001101011_011_0_000110101101;
      patterns[17244] = 29'b0_100001101011_100_1_010000110101;
      patterns[17245] = 29'b0_100001101011_101_1_101000011010;
      patterns[17246] = 29'b0_100001101011_110_0_100001101011;
      patterns[17247] = 29'b0_100001101011_111_0_100001101011;
      patterns[17248] = 29'b0_100001101100_000_0_100001101100;
      patterns[17249] = 29'b0_100001101100_001_0_101100100001;
      patterns[17250] = 29'b0_100001101100_010_1_000011011000;
      patterns[17251] = 29'b0_100001101100_011_0_000110110001;
      patterns[17252] = 29'b0_100001101100_100_0_010000110110;
      patterns[17253] = 29'b0_100001101100_101_0_001000011011;
      patterns[17254] = 29'b0_100001101100_110_0_100001101100;
      patterns[17255] = 29'b0_100001101100_111_0_100001101100;
      patterns[17256] = 29'b0_100001101101_000_0_100001101101;
      patterns[17257] = 29'b0_100001101101_001_0_101101100001;
      patterns[17258] = 29'b0_100001101101_010_1_000011011010;
      patterns[17259] = 29'b0_100001101101_011_0_000110110101;
      patterns[17260] = 29'b0_100001101101_100_1_010000110110;
      patterns[17261] = 29'b0_100001101101_101_0_101000011011;
      patterns[17262] = 29'b0_100001101101_110_0_100001101101;
      patterns[17263] = 29'b0_100001101101_111_0_100001101101;
      patterns[17264] = 29'b0_100001101110_000_0_100001101110;
      patterns[17265] = 29'b0_100001101110_001_0_101110100001;
      patterns[17266] = 29'b0_100001101110_010_1_000011011100;
      patterns[17267] = 29'b0_100001101110_011_0_000110111001;
      patterns[17268] = 29'b0_100001101110_100_0_010000110111;
      patterns[17269] = 29'b0_100001101110_101_1_001000011011;
      patterns[17270] = 29'b0_100001101110_110_0_100001101110;
      patterns[17271] = 29'b0_100001101110_111_0_100001101110;
      patterns[17272] = 29'b0_100001101111_000_0_100001101111;
      patterns[17273] = 29'b0_100001101111_001_0_101111100001;
      patterns[17274] = 29'b0_100001101111_010_1_000011011110;
      patterns[17275] = 29'b0_100001101111_011_0_000110111101;
      patterns[17276] = 29'b0_100001101111_100_1_010000110111;
      patterns[17277] = 29'b0_100001101111_101_1_101000011011;
      patterns[17278] = 29'b0_100001101111_110_0_100001101111;
      patterns[17279] = 29'b0_100001101111_111_0_100001101111;
      patterns[17280] = 29'b0_100001110000_000_0_100001110000;
      patterns[17281] = 29'b0_100001110000_001_0_110000100001;
      patterns[17282] = 29'b0_100001110000_010_1_000011100000;
      patterns[17283] = 29'b0_100001110000_011_0_000111000001;
      patterns[17284] = 29'b0_100001110000_100_0_010000111000;
      patterns[17285] = 29'b0_100001110000_101_0_001000011100;
      patterns[17286] = 29'b0_100001110000_110_0_100001110000;
      patterns[17287] = 29'b0_100001110000_111_0_100001110000;
      patterns[17288] = 29'b0_100001110001_000_0_100001110001;
      patterns[17289] = 29'b0_100001110001_001_0_110001100001;
      patterns[17290] = 29'b0_100001110001_010_1_000011100010;
      patterns[17291] = 29'b0_100001110001_011_0_000111000101;
      patterns[17292] = 29'b0_100001110001_100_1_010000111000;
      patterns[17293] = 29'b0_100001110001_101_0_101000011100;
      patterns[17294] = 29'b0_100001110001_110_0_100001110001;
      patterns[17295] = 29'b0_100001110001_111_0_100001110001;
      patterns[17296] = 29'b0_100001110010_000_0_100001110010;
      patterns[17297] = 29'b0_100001110010_001_0_110010100001;
      patterns[17298] = 29'b0_100001110010_010_1_000011100100;
      patterns[17299] = 29'b0_100001110010_011_0_000111001001;
      patterns[17300] = 29'b0_100001110010_100_0_010000111001;
      patterns[17301] = 29'b0_100001110010_101_1_001000011100;
      patterns[17302] = 29'b0_100001110010_110_0_100001110010;
      patterns[17303] = 29'b0_100001110010_111_0_100001110010;
      patterns[17304] = 29'b0_100001110011_000_0_100001110011;
      patterns[17305] = 29'b0_100001110011_001_0_110011100001;
      patterns[17306] = 29'b0_100001110011_010_1_000011100110;
      patterns[17307] = 29'b0_100001110011_011_0_000111001101;
      patterns[17308] = 29'b0_100001110011_100_1_010000111001;
      patterns[17309] = 29'b0_100001110011_101_1_101000011100;
      patterns[17310] = 29'b0_100001110011_110_0_100001110011;
      patterns[17311] = 29'b0_100001110011_111_0_100001110011;
      patterns[17312] = 29'b0_100001110100_000_0_100001110100;
      patterns[17313] = 29'b0_100001110100_001_0_110100100001;
      patterns[17314] = 29'b0_100001110100_010_1_000011101000;
      patterns[17315] = 29'b0_100001110100_011_0_000111010001;
      patterns[17316] = 29'b0_100001110100_100_0_010000111010;
      patterns[17317] = 29'b0_100001110100_101_0_001000011101;
      patterns[17318] = 29'b0_100001110100_110_0_100001110100;
      patterns[17319] = 29'b0_100001110100_111_0_100001110100;
      patterns[17320] = 29'b0_100001110101_000_0_100001110101;
      patterns[17321] = 29'b0_100001110101_001_0_110101100001;
      patterns[17322] = 29'b0_100001110101_010_1_000011101010;
      patterns[17323] = 29'b0_100001110101_011_0_000111010101;
      patterns[17324] = 29'b0_100001110101_100_1_010000111010;
      patterns[17325] = 29'b0_100001110101_101_0_101000011101;
      patterns[17326] = 29'b0_100001110101_110_0_100001110101;
      patterns[17327] = 29'b0_100001110101_111_0_100001110101;
      patterns[17328] = 29'b0_100001110110_000_0_100001110110;
      patterns[17329] = 29'b0_100001110110_001_0_110110100001;
      patterns[17330] = 29'b0_100001110110_010_1_000011101100;
      patterns[17331] = 29'b0_100001110110_011_0_000111011001;
      patterns[17332] = 29'b0_100001110110_100_0_010000111011;
      patterns[17333] = 29'b0_100001110110_101_1_001000011101;
      patterns[17334] = 29'b0_100001110110_110_0_100001110110;
      patterns[17335] = 29'b0_100001110110_111_0_100001110110;
      patterns[17336] = 29'b0_100001110111_000_0_100001110111;
      patterns[17337] = 29'b0_100001110111_001_0_110111100001;
      patterns[17338] = 29'b0_100001110111_010_1_000011101110;
      patterns[17339] = 29'b0_100001110111_011_0_000111011101;
      patterns[17340] = 29'b0_100001110111_100_1_010000111011;
      patterns[17341] = 29'b0_100001110111_101_1_101000011101;
      patterns[17342] = 29'b0_100001110111_110_0_100001110111;
      patterns[17343] = 29'b0_100001110111_111_0_100001110111;
      patterns[17344] = 29'b0_100001111000_000_0_100001111000;
      patterns[17345] = 29'b0_100001111000_001_0_111000100001;
      patterns[17346] = 29'b0_100001111000_010_1_000011110000;
      patterns[17347] = 29'b0_100001111000_011_0_000111100001;
      patterns[17348] = 29'b0_100001111000_100_0_010000111100;
      patterns[17349] = 29'b0_100001111000_101_0_001000011110;
      patterns[17350] = 29'b0_100001111000_110_0_100001111000;
      patterns[17351] = 29'b0_100001111000_111_0_100001111000;
      patterns[17352] = 29'b0_100001111001_000_0_100001111001;
      patterns[17353] = 29'b0_100001111001_001_0_111001100001;
      patterns[17354] = 29'b0_100001111001_010_1_000011110010;
      patterns[17355] = 29'b0_100001111001_011_0_000111100101;
      patterns[17356] = 29'b0_100001111001_100_1_010000111100;
      patterns[17357] = 29'b0_100001111001_101_0_101000011110;
      patterns[17358] = 29'b0_100001111001_110_0_100001111001;
      patterns[17359] = 29'b0_100001111001_111_0_100001111001;
      patterns[17360] = 29'b0_100001111010_000_0_100001111010;
      patterns[17361] = 29'b0_100001111010_001_0_111010100001;
      patterns[17362] = 29'b0_100001111010_010_1_000011110100;
      patterns[17363] = 29'b0_100001111010_011_0_000111101001;
      patterns[17364] = 29'b0_100001111010_100_0_010000111101;
      patterns[17365] = 29'b0_100001111010_101_1_001000011110;
      patterns[17366] = 29'b0_100001111010_110_0_100001111010;
      patterns[17367] = 29'b0_100001111010_111_0_100001111010;
      patterns[17368] = 29'b0_100001111011_000_0_100001111011;
      patterns[17369] = 29'b0_100001111011_001_0_111011100001;
      patterns[17370] = 29'b0_100001111011_010_1_000011110110;
      patterns[17371] = 29'b0_100001111011_011_0_000111101101;
      patterns[17372] = 29'b0_100001111011_100_1_010000111101;
      patterns[17373] = 29'b0_100001111011_101_1_101000011110;
      patterns[17374] = 29'b0_100001111011_110_0_100001111011;
      patterns[17375] = 29'b0_100001111011_111_0_100001111011;
      patterns[17376] = 29'b0_100001111100_000_0_100001111100;
      patterns[17377] = 29'b0_100001111100_001_0_111100100001;
      patterns[17378] = 29'b0_100001111100_010_1_000011111000;
      patterns[17379] = 29'b0_100001111100_011_0_000111110001;
      patterns[17380] = 29'b0_100001111100_100_0_010000111110;
      patterns[17381] = 29'b0_100001111100_101_0_001000011111;
      patterns[17382] = 29'b0_100001111100_110_0_100001111100;
      patterns[17383] = 29'b0_100001111100_111_0_100001111100;
      patterns[17384] = 29'b0_100001111101_000_0_100001111101;
      patterns[17385] = 29'b0_100001111101_001_0_111101100001;
      patterns[17386] = 29'b0_100001111101_010_1_000011111010;
      patterns[17387] = 29'b0_100001111101_011_0_000111110101;
      patterns[17388] = 29'b0_100001111101_100_1_010000111110;
      patterns[17389] = 29'b0_100001111101_101_0_101000011111;
      patterns[17390] = 29'b0_100001111101_110_0_100001111101;
      patterns[17391] = 29'b0_100001111101_111_0_100001111101;
      patterns[17392] = 29'b0_100001111110_000_0_100001111110;
      patterns[17393] = 29'b0_100001111110_001_0_111110100001;
      patterns[17394] = 29'b0_100001111110_010_1_000011111100;
      patterns[17395] = 29'b0_100001111110_011_0_000111111001;
      patterns[17396] = 29'b0_100001111110_100_0_010000111111;
      patterns[17397] = 29'b0_100001111110_101_1_001000011111;
      patterns[17398] = 29'b0_100001111110_110_0_100001111110;
      patterns[17399] = 29'b0_100001111110_111_0_100001111110;
      patterns[17400] = 29'b0_100001111111_000_0_100001111111;
      patterns[17401] = 29'b0_100001111111_001_0_111111100001;
      patterns[17402] = 29'b0_100001111111_010_1_000011111110;
      patterns[17403] = 29'b0_100001111111_011_0_000111111101;
      patterns[17404] = 29'b0_100001111111_100_1_010000111111;
      patterns[17405] = 29'b0_100001111111_101_1_101000011111;
      patterns[17406] = 29'b0_100001111111_110_0_100001111111;
      patterns[17407] = 29'b0_100001111111_111_0_100001111111;
      patterns[17408] = 29'b0_100010000000_000_0_100010000000;
      patterns[17409] = 29'b0_100010000000_001_0_000000100010;
      patterns[17410] = 29'b0_100010000000_010_1_000100000000;
      patterns[17411] = 29'b0_100010000000_011_0_001000000001;
      patterns[17412] = 29'b0_100010000000_100_0_010001000000;
      patterns[17413] = 29'b0_100010000000_101_0_001000100000;
      patterns[17414] = 29'b0_100010000000_110_0_100010000000;
      patterns[17415] = 29'b0_100010000000_111_0_100010000000;
      patterns[17416] = 29'b0_100010000001_000_0_100010000001;
      patterns[17417] = 29'b0_100010000001_001_0_000001100010;
      patterns[17418] = 29'b0_100010000001_010_1_000100000010;
      patterns[17419] = 29'b0_100010000001_011_0_001000000101;
      patterns[17420] = 29'b0_100010000001_100_1_010001000000;
      patterns[17421] = 29'b0_100010000001_101_0_101000100000;
      patterns[17422] = 29'b0_100010000001_110_0_100010000001;
      patterns[17423] = 29'b0_100010000001_111_0_100010000001;
      patterns[17424] = 29'b0_100010000010_000_0_100010000010;
      patterns[17425] = 29'b0_100010000010_001_0_000010100010;
      patterns[17426] = 29'b0_100010000010_010_1_000100000100;
      patterns[17427] = 29'b0_100010000010_011_0_001000001001;
      patterns[17428] = 29'b0_100010000010_100_0_010001000001;
      patterns[17429] = 29'b0_100010000010_101_1_001000100000;
      patterns[17430] = 29'b0_100010000010_110_0_100010000010;
      patterns[17431] = 29'b0_100010000010_111_0_100010000010;
      patterns[17432] = 29'b0_100010000011_000_0_100010000011;
      patterns[17433] = 29'b0_100010000011_001_0_000011100010;
      patterns[17434] = 29'b0_100010000011_010_1_000100000110;
      patterns[17435] = 29'b0_100010000011_011_0_001000001101;
      patterns[17436] = 29'b0_100010000011_100_1_010001000001;
      patterns[17437] = 29'b0_100010000011_101_1_101000100000;
      patterns[17438] = 29'b0_100010000011_110_0_100010000011;
      patterns[17439] = 29'b0_100010000011_111_0_100010000011;
      patterns[17440] = 29'b0_100010000100_000_0_100010000100;
      patterns[17441] = 29'b0_100010000100_001_0_000100100010;
      patterns[17442] = 29'b0_100010000100_010_1_000100001000;
      patterns[17443] = 29'b0_100010000100_011_0_001000010001;
      patterns[17444] = 29'b0_100010000100_100_0_010001000010;
      patterns[17445] = 29'b0_100010000100_101_0_001000100001;
      patterns[17446] = 29'b0_100010000100_110_0_100010000100;
      patterns[17447] = 29'b0_100010000100_111_0_100010000100;
      patterns[17448] = 29'b0_100010000101_000_0_100010000101;
      patterns[17449] = 29'b0_100010000101_001_0_000101100010;
      patterns[17450] = 29'b0_100010000101_010_1_000100001010;
      patterns[17451] = 29'b0_100010000101_011_0_001000010101;
      patterns[17452] = 29'b0_100010000101_100_1_010001000010;
      patterns[17453] = 29'b0_100010000101_101_0_101000100001;
      patterns[17454] = 29'b0_100010000101_110_0_100010000101;
      patterns[17455] = 29'b0_100010000101_111_0_100010000101;
      patterns[17456] = 29'b0_100010000110_000_0_100010000110;
      patterns[17457] = 29'b0_100010000110_001_0_000110100010;
      patterns[17458] = 29'b0_100010000110_010_1_000100001100;
      patterns[17459] = 29'b0_100010000110_011_0_001000011001;
      patterns[17460] = 29'b0_100010000110_100_0_010001000011;
      patterns[17461] = 29'b0_100010000110_101_1_001000100001;
      patterns[17462] = 29'b0_100010000110_110_0_100010000110;
      patterns[17463] = 29'b0_100010000110_111_0_100010000110;
      patterns[17464] = 29'b0_100010000111_000_0_100010000111;
      patterns[17465] = 29'b0_100010000111_001_0_000111100010;
      patterns[17466] = 29'b0_100010000111_010_1_000100001110;
      patterns[17467] = 29'b0_100010000111_011_0_001000011101;
      patterns[17468] = 29'b0_100010000111_100_1_010001000011;
      patterns[17469] = 29'b0_100010000111_101_1_101000100001;
      patterns[17470] = 29'b0_100010000111_110_0_100010000111;
      patterns[17471] = 29'b0_100010000111_111_0_100010000111;
      patterns[17472] = 29'b0_100010001000_000_0_100010001000;
      patterns[17473] = 29'b0_100010001000_001_0_001000100010;
      patterns[17474] = 29'b0_100010001000_010_1_000100010000;
      patterns[17475] = 29'b0_100010001000_011_0_001000100001;
      patterns[17476] = 29'b0_100010001000_100_0_010001000100;
      patterns[17477] = 29'b0_100010001000_101_0_001000100010;
      patterns[17478] = 29'b0_100010001000_110_0_100010001000;
      patterns[17479] = 29'b0_100010001000_111_0_100010001000;
      patterns[17480] = 29'b0_100010001001_000_0_100010001001;
      patterns[17481] = 29'b0_100010001001_001_0_001001100010;
      patterns[17482] = 29'b0_100010001001_010_1_000100010010;
      patterns[17483] = 29'b0_100010001001_011_0_001000100101;
      patterns[17484] = 29'b0_100010001001_100_1_010001000100;
      patterns[17485] = 29'b0_100010001001_101_0_101000100010;
      patterns[17486] = 29'b0_100010001001_110_0_100010001001;
      patterns[17487] = 29'b0_100010001001_111_0_100010001001;
      patterns[17488] = 29'b0_100010001010_000_0_100010001010;
      patterns[17489] = 29'b0_100010001010_001_0_001010100010;
      patterns[17490] = 29'b0_100010001010_010_1_000100010100;
      patterns[17491] = 29'b0_100010001010_011_0_001000101001;
      patterns[17492] = 29'b0_100010001010_100_0_010001000101;
      patterns[17493] = 29'b0_100010001010_101_1_001000100010;
      patterns[17494] = 29'b0_100010001010_110_0_100010001010;
      patterns[17495] = 29'b0_100010001010_111_0_100010001010;
      patterns[17496] = 29'b0_100010001011_000_0_100010001011;
      patterns[17497] = 29'b0_100010001011_001_0_001011100010;
      patterns[17498] = 29'b0_100010001011_010_1_000100010110;
      patterns[17499] = 29'b0_100010001011_011_0_001000101101;
      patterns[17500] = 29'b0_100010001011_100_1_010001000101;
      patterns[17501] = 29'b0_100010001011_101_1_101000100010;
      patterns[17502] = 29'b0_100010001011_110_0_100010001011;
      patterns[17503] = 29'b0_100010001011_111_0_100010001011;
      patterns[17504] = 29'b0_100010001100_000_0_100010001100;
      patterns[17505] = 29'b0_100010001100_001_0_001100100010;
      patterns[17506] = 29'b0_100010001100_010_1_000100011000;
      patterns[17507] = 29'b0_100010001100_011_0_001000110001;
      patterns[17508] = 29'b0_100010001100_100_0_010001000110;
      patterns[17509] = 29'b0_100010001100_101_0_001000100011;
      patterns[17510] = 29'b0_100010001100_110_0_100010001100;
      patterns[17511] = 29'b0_100010001100_111_0_100010001100;
      patterns[17512] = 29'b0_100010001101_000_0_100010001101;
      patterns[17513] = 29'b0_100010001101_001_0_001101100010;
      patterns[17514] = 29'b0_100010001101_010_1_000100011010;
      patterns[17515] = 29'b0_100010001101_011_0_001000110101;
      patterns[17516] = 29'b0_100010001101_100_1_010001000110;
      patterns[17517] = 29'b0_100010001101_101_0_101000100011;
      patterns[17518] = 29'b0_100010001101_110_0_100010001101;
      patterns[17519] = 29'b0_100010001101_111_0_100010001101;
      patterns[17520] = 29'b0_100010001110_000_0_100010001110;
      patterns[17521] = 29'b0_100010001110_001_0_001110100010;
      patterns[17522] = 29'b0_100010001110_010_1_000100011100;
      patterns[17523] = 29'b0_100010001110_011_0_001000111001;
      patterns[17524] = 29'b0_100010001110_100_0_010001000111;
      patterns[17525] = 29'b0_100010001110_101_1_001000100011;
      patterns[17526] = 29'b0_100010001110_110_0_100010001110;
      patterns[17527] = 29'b0_100010001110_111_0_100010001110;
      patterns[17528] = 29'b0_100010001111_000_0_100010001111;
      patterns[17529] = 29'b0_100010001111_001_0_001111100010;
      patterns[17530] = 29'b0_100010001111_010_1_000100011110;
      patterns[17531] = 29'b0_100010001111_011_0_001000111101;
      patterns[17532] = 29'b0_100010001111_100_1_010001000111;
      patterns[17533] = 29'b0_100010001111_101_1_101000100011;
      patterns[17534] = 29'b0_100010001111_110_0_100010001111;
      patterns[17535] = 29'b0_100010001111_111_0_100010001111;
      patterns[17536] = 29'b0_100010010000_000_0_100010010000;
      patterns[17537] = 29'b0_100010010000_001_0_010000100010;
      patterns[17538] = 29'b0_100010010000_010_1_000100100000;
      patterns[17539] = 29'b0_100010010000_011_0_001001000001;
      patterns[17540] = 29'b0_100010010000_100_0_010001001000;
      patterns[17541] = 29'b0_100010010000_101_0_001000100100;
      patterns[17542] = 29'b0_100010010000_110_0_100010010000;
      patterns[17543] = 29'b0_100010010000_111_0_100010010000;
      patterns[17544] = 29'b0_100010010001_000_0_100010010001;
      patterns[17545] = 29'b0_100010010001_001_0_010001100010;
      patterns[17546] = 29'b0_100010010001_010_1_000100100010;
      patterns[17547] = 29'b0_100010010001_011_0_001001000101;
      patterns[17548] = 29'b0_100010010001_100_1_010001001000;
      patterns[17549] = 29'b0_100010010001_101_0_101000100100;
      patterns[17550] = 29'b0_100010010001_110_0_100010010001;
      patterns[17551] = 29'b0_100010010001_111_0_100010010001;
      patterns[17552] = 29'b0_100010010010_000_0_100010010010;
      patterns[17553] = 29'b0_100010010010_001_0_010010100010;
      patterns[17554] = 29'b0_100010010010_010_1_000100100100;
      patterns[17555] = 29'b0_100010010010_011_0_001001001001;
      patterns[17556] = 29'b0_100010010010_100_0_010001001001;
      patterns[17557] = 29'b0_100010010010_101_1_001000100100;
      patterns[17558] = 29'b0_100010010010_110_0_100010010010;
      patterns[17559] = 29'b0_100010010010_111_0_100010010010;
      patterns[17560] = 29'b0_100010010011_000_0_100010010011;
      patterns[17561] = 29'b0_100010010011_001_0_010011100010;
      patterns[17562] = 29'b0_100010010011_010_1_000100100110;
      patterns[17563] = 29'b0_100010010011_011_0_001001001101;
      patterns[17564] = 29'b0_100010010011_100_1_010001001001;
      patterns[17565] = 29'b0_100010010011_101_1_101000100100;
      patterns[17566] = 29'b0_100010010011_110_0_100010010011;
      patterns[17567] = 29'b0_100010010011_111_0_100010010011;
      patterns[17568] = 29'b0_100010010100_000_0_100010010100;
      patterns[17569] = 29'b0_100010010100_001_0_010100100010;
      patterns[17570] = 29'b0_100010010100_010_1_000100101000;
      patterns[17571] = 29'b0_100010010100_011_0_001001010001;
      patterns[17572] = 29'b0_100010010100_100_0_010001001010;
      patterns[17573] = 29'b0_100010010100_101_0_001000100101;
      patterns[17574] = 29'b0_100010010100_110_0_100010010100;
      patterns[17575] = 29'b0_100010010100_111_0_100010010100;
      patterns[17576] = 29'b0_100010010101_000_0_100010010101;
      patterns[17577] = 29'b0_100010010101_001_0_010101100010;
      patterns[17578] = 29'b0_100010010101_010_1_000100101010;
      patterns[17579] = 29'b0_100010010101_011_0_001001010101;
      patterns[17580] = 29'b0_100010010101_100_1_010001001010;
      patterns[17581] = 29'b0_100010010101_101_0_101000100101;
      patterns[17582] = 29'b0_100010010101_110_0_100010010101;
      patterns[17583] = 29'b0_100010010101_111_0_100010010101;
      patterns[17584] = 29'b0_100010010110_000_0_100010010110;
      patterns[17585] = 29'b0_100010010110_001_0_010110100010;
      patterns[17586] = 29'b0_100010010110_010_1_000100101100;
      patterns[17587] = 29'b0_100010010110_011_0_001001011001;
      patterns[17588] = 29'b0_100010010110_100_0_010001001011;
      patterns[17589] = 29'b0_100010010110_101_1_001000100101;
      patterns[17590] = 29'b0_100010010110_110_0_100010010110;
      patterns[17591] = 29'b0_100010010110_111_0_100010010110;
      patterns[17592] = 29'b0_100010010111_000_0_100010010111;
      patterns[17593] = 29'b0_100010010111_001_0_010111100010;
      patterns[17594] = 29'b0_100010010111_010_1_000100101110;
      patterns[17595] = 29'b0_100010010111_011_0_001001011101;
      patterns[17596] = 29'b0_100010010111_100_1_010001001011;
      patterns[17597] = 29'b0_100010010111_101_1_101000100101;
      patterns[17598] = 29'b0_100010010111_110_0_100010010111;
      patterns[17599] = 29'b0_100010010111_111_0_100010010111;
      patterns[17600] = 29'b0_100010011000_000_0_100010011000;
      patterns[17601] = 29'b0_100010011000_001_0_011000100010;
      patterns[17602] = 29'b0_100010011000_010_1_000100110000;
      patterns[17603] = 29'b0_100010011000_011_0_001001100001;
      patterns[17604] = 29'b0_100010011000_100_0_010001001100;
      patterns[17605] = 29'b0_100010011000_101_0_001000100110;
      patterns[17606] = 29'b0_100010011000_110_0_100010011000;
      patterns[17607] = 29'b0_100010011000_111_0_100010011000;
      patterns[17608] = 29'b0_100010011001_000_0_100010011001;
      patterns[17609] = 29'b0_100010011001_001_0_011001100010;
      patterns[17610] = 29'b0_100010011001_010_1_000100110010;
      patterns[17611] = 29'b0_100010011001_011_0_001001100101;
      patterns[17612] = 29'b0_100010011001_100_1_010001001100;
      patterns[17613] = 29'b0_100010011001_101_0_101000100110;
      patterns[17614] = 29'b0_100010011001_110_0_100010011001;
      patterns[17615] = 29'b0_100010011001_111_0_100010011001;
      patterns[17616] = 29'b0_100010011010_000_0_100010011010;
      patterns[17617] = 29'b0_100010011010_001_0_011010100010;
      patterns[17618] = 29'b0_100010011010_010_1_000100110100;
      patterns[17619] = 29'b0_100010011010_011_0_001001101001;
      patterns[17620] = 29'b0_100010011010_100_0_010001001101;
      patterns[17621] = 29'b0_100010011010_101_1_001000100110;
      patterns[17622] = 29'b0_100010011010_110_0_100010011010;
      patterns[17623] = 29'b0_100010011010_111_0_100010011010;
      patterns[17624] = 29'b0_100010011011_000_0_100010011011;
      patterns[17625] = 29'b0_100010011011_001_0_011011100010;
      patterns[17626] = 29'b0_100010011011_010_1_000100110110;
      patterns[17627] = 29'b0_100010011011_011_0_001001101101;
      patterns[17628] = 29'b0_100010011011_100_1_010001001101;
      patterns[17629] = 29'b0_100010011011_101_1_101000100110;
      patterns[17630] = 29'b0_100010011011_110_0_100010011011;
      patterns[17631] = 29'b0_100010011011_111_0_100010011011;
      patterns[17632] = 29'b0_100010011100_000_0_100010011100;
      patterns[17633] = 29'b0_100010011100_001_0_011100100010;
      patterns[17634] = 29'b0_100010011100_010_1_000100111000;
      patterns[17635] = 29'b0_100010011100_011_0_001001110001;
      patterns[17636] = 29'b0_100010011100_100_0_010001001110;
      patterns[17637] = 29'b0_100010011100_101_0_001000100111;
      patterns[17638] = 29'b0_100010011100_110_0_100010011100;
      patterns[17639] = 29'b0_100010011100_111_0_100010011100;
      patterns[17640] = 29'b0_100010011101_000_0_100010011101;
      patterns[17641] = 29'b0_100010011101_001_0_011101100010;
      patterns[17642] = 29'b0_100010011101_010_1_000100111010;
      patterns[17643] = 29'b0_100010011101_011_0_001001110101;
      patterns[17644] = 29'b0_100010011101_100_1_010001001110;
      patterns[17645] = 29'b0_100010011101_101_0_101000100111;
      patterns[17646] = 29'b0_100010011101_110_0_100010011101;
      patterns[17647] = 29'b0_100010011101_111_0_100010011101;
      patterns[17648] = 29'b0_100010011110_000_0_100010011110;
      patterns[17649] = 29'b0_100010011110_001_0_011110100010;
      patterns[17650] = 29'b0_100010011110_010_1_000100111100;
      patterns[17651] = 29'b0_100010011110_011_0_001001111001;
      patterns[17652] = 29'b0_100010011110_100_0_010001001111;
      patterns[17653] = 29'b0_100010011110_101_1_001000100111;
      patterns[17654] = 29'b0_100010011110_110_0_100010011110;
      patterns[17655] = 29'b0_100010011110_111_0_100010011110;
      patterns[17656] = 29'b0_100010011111_000_0_100010011111;
      patterns[17657] = 29'b0_100010011111_001_0_011111100010;
      patterns[17658] = 29'b0_100010011111_010_1_000100111110;
      patterns[17659] = 29'b0_100010011111_011_0_001001111101;
      patterns[17660] = 29'b0_100010011111_100_1_010001001111;
      patterns[17661] = 29'b0_100010011111_101_1_101000100111;
      patterns[17662] = 29'b0_100010011111_110_0_100010011111;
      patterns[17663] = 29'b0_100010011111_111_0_100010011111;
      patterns[17664] = 29'b0_100010100000_000_0_100010100000;
      patterns[17665] = 29'b0_100010100000_001_0_100000100010;
      patterns[17666] = 29'b0_100010100000_010_1_000101000000;
      patterns[17667] = 29'b0_100010100000_011_0_001010000001;
      patterns[17668] = 29'b0_100010100000_100_0_010001010000;
      patterns[17669] = 29'b0_100010100000_101_0_001000101000;
      patterns[17670] = 29'b0_100010100000_110_0_100010100000;
      patterns[17671] = 29'b0_100010100000_111_0_100010100000;
      patterns[17672] = 29'b0_100010100001_000_0_100010100001;
      patterns[17673] = 29'b0_100010100001_001_0_100001100010;
      patterns[17674] = 29'b0_100010100001_010_1_000101000010;
      patterns[17675] = 29'b0_100010100001_011_0_001010000101;
      patterns[17676] = 29'b0_100010100001_100_1_010001010000;
      patterns[17677] = 29'b0_100010100001_101_0_101000101000;
      patterns[17678] = 29'b0_100010100001_110_0_100010100001;
      patterns[17679] = 29'b0_100010100001_111_0_100010100001;
      patterns[17680] = 29'b0_100010100010_000_0_100010100010;
      patterns[17681] = 29'b0_100010100010_001_0_100010100010;
      patterns[17682] = 29'b0_100010100010_010_1_000101000100;
      patterns[17683] = 29'b0_100010100010_011_0_001010001001;
      patterns[17684] = 29'b0_100010100010_100_0_010001010001;
      patterns[17685] = 29'b0_100010100010_101_1_001000101000;
      patterns[17686] = 29'b0_100010100010_110_0_100010100010;
      patterns[17687] = 29'b0_100010100010_111_0_100010100010;
      patterns[17688] = 29'b0_100010100011_000_0_100010100011;
      patterns[17689] = 29'b0_100010100011_001_0_100011100010;
      patterns[17690] = 29'b0_100010100011_010_1_000101000110;
      patterns[17691] = 29'b0_100010100011_011_0_001010001101;
      patterns[17692] = 29'b0_100010100011_100_1_010001010001;
      patterns[17693] = 29'b0_100010100011_101_1_101000101000;
      patterns[17694] = 29'b0_100010100011_110_0_100010100011;
      patterns[17695] = 29'b0_100010100011_111_0_100010100011;
      patterns[17696] = 29'b0_100010100100_000_0_100010100100;
      patterns[17697] = 29'b0_100010100100_001_0_100100100010;
      patterns[17698] = 29'b0_100010100100_010_1_000101001000;
      patterns[17699] = 29'b0_100010100100_011_0_001010010001;
      patterns[17700] = 29'b0_100010100100_100_0_010001010010;
      patterns[17701] = 29'b0_100010100100_101_0_001000101001;
      patterns[17702] = 29'b0_100010100100_110_0_100010100100;
      patterns[17703] = 29'b0_100010100100_111_0_100010100100;
      patterns[17704] = 29'b0_100010100101_000_0_100010100101;
      patterns[17705] = 29'b0_100010100101_001_0_100101100010;
      patterns[17706] = 29'b0_100010100101_010_1_000101001010;
      patterns[17707] = 29'b0_100010100101_011_0_001010010101;
      patterns[17708] = 29'b0_100010100101_100_1_010001010010;
      patterns[17709] = 29'b0_100010100101_101_0_101000101001;
      patterns[17710] = 29'b0_100010100101_110_0_100010100101;
      patterns[17711] = 29'b0_100010100101_111_0_100010100101;
      patterns[17712] = 29'b0_100010100110_000_0_100010100110;
      patterns[17713] = 29'b0_100010100110_001_0_100110100010;
      patterns[17714] = 29'b0_100010100110_010_1_000101001100;
      patterns[17715] = 29'b0_100010100110_011_0_001010011001;
      patterns[17716] = 29'b0_100010100110_100_0_010001010011;
      patterns[17717] = 29'b0_100010100110_101_1_001000101001;
      patterns[17718] = 29'b0_100010100110_110_0_100010100110;
      patterns[17719] = 29'b0_100010100110_111_0_100010100110;
      patterns[17720] = 29'b0_100010100111_000_0_100010100111;
      patterns[17721] = 29'b0_100010100111_001_0_100111100010;
      patterns[17722] = 29'b0_100010100111_010_1_000101001110;
      patterns[17723] = 29'b0_100010100111_011_0_001010011101;
      patterns[17724] = 29'b0_100010100111_100_1_010001010011;
      patterns[17725] = 29'b0_100010100111_101_1_101000101001;
      patterns[17726] = 29'b0_100010100111_110_0_100010100111;
      patterns[17727] = 29'b0_100010100111_111_0_100010100111;
      patterns[17728] = 29'b0_100010101000_000_0_100010101000;
      patterns[17729] = 29'b0_100010101000_001_0_101000100010;
      patterns[17730] = 29'b0_100010101000_010_1_000101010000;
      patterns[17731] = 29'b0_100010101000_011_0_001010100001;
      patterns[17732] = 29'b0_100010101000_100_0_010001010100;
      patterns[17733] = 29'b0_100010101000_101_0_001000101010;
      patterns[17734] = 29'b0_100010101000_110_0_100010101000;
      patterns[17735] = 29'b0_100010101000_111_0_100010101000;
      patterns[17736] = 29'b0_100010101001_000_0_100010101001;
      patterns[17737] = 29'b0_100010101001_001_0_101001100010;
      patterns[17738] = 29'b0_100010101001_010_1_000101010010;
      patterns[17739] = 29'b0_100010101001_011_0_001010100101;
      patterns[17740] = 29'b0_100010101001_100_1_010001010100;
      patterns[17741] = 29'b0_100010101001_101_0_101000101010;
      patterns[17742] = 29'b0_100010101001_110_0_100010101001;
      patterns[17743] = 29'b0_100010101001_111_0_100010101001;
      patterns[17744] = 29'b0_100010101010_000_0_100010101010;
      patterns[17745] = 29'b0_100010101010_001_0_101010100010;
      patterns[17746] = 29'b0_100010101010_010_1_000101010100;
      patterns[17747] = 29'b0_100010101010_011_0_001010101001;
      patterns[17748] = 29'b0_100010101010_100_0_010001010101;
      patterns[17749] = 29'b0_100010101010_101_1_001000101010;
      patterns[17750] = 29'b0_100010101010_110_0_100010101010;
      patterns[17751] = 29'b0_100010101010_111_0_100010101010;
      patterns[17752] = 29'b0_100010101011_000_0_100010101011;
      patterns[17753] = 29'b0_100010101011_001_0_101011100010;
      patterns[17754] = 29'b0_100010101011_010_1_000101010110;
      patterns[17755] = 29'b0_100010101011_011_0_001010101101;
      patterns[17756] = 29'b0_100010101011_100_1_010001010101;
      patterns[17757] = 29'b0_100010101011_101_1_101000101010;
      patterns[17758] = 29'b0_100010101011_110_0_100010101011;
      patterns[17759] = 29'b0_100010101011_111_0_100010101011;
      patterns[17760] = 29'b0_100010101100_000_0_100010101100;
      patterns[17761] = 29'b0_100010101100_001_0_101100100010;
      patterns[17762] = 29'b0_100010101100_010_1_000101011000;
      patterns[17763] = 29'b0_100010101100_011_0_001010110001;
      patterns[17764] = 29'b0_100010101100_100_0_010001010110;
      patterns[17765] = 29'b0_100010101100_101_0_001000101011;
      patterns[17766] = 29'b0_100010101100_110_0_100010101100;
      patterns[17767] = 29'b0_100010101100_111_0_100010101100;
      patterns[17768] = 29'b0_100010101101_000_0_100010101101;
      patterns[17769] = 29'b0_100010101101_001_0_101101100010;
      patterns[17770] = 29'b0_100010101101_010_1_000101011010;
      patterns[17771] = 29'b0_100010101101_011_0_001010110101;
      patterns[17772] = 29'b0_100010101101_100_1_010001010110;
      patterns[17773] = 29'b0_100010101101_101_0_101000101011;
      patterns[17774] = 29'b0_100010101101_110_0_100010101101;
      patterns[17775] = 29'b0_100010101101_111_0_100010101101;
      patterns[17776] = 29'b0_100010101110_000_0_100010101110;
      patterns[17777] = 29'b0_100010101110_001_0_101110100010;
      patterns[17778] = 29'b0_100010101110_010_1_000101011100;
      patterns[17779] = 29'b0_100010101110_011_0_001010111001;
      patterns[17780] = 29'b0_100010101110_100_0_010001010111;
      patterns[17781] = 29'b0_100010101110_101_1_001000101011;
      patterns[17782] = 29'b0_100010101110_110_0_100010101110;
      patterns[17783] = 29'b0_100010101110_111_0_100010101110;
      patterns[17784] = 29'b0_100010101111_000_0_100010101111;
      patterns[17785] = 29'b0_100010101111_001_0_101111100010;
      patterns[17786] = 29'b0_100010101111_010_1_000101011110;
      patterns[17787] = 29'b0_100010101111_011_0_001010111101;
      patterns[17788] = 29'b0_100010101111_100_1_010001010111;
      patterns[17789] = 29'b0_100010101111_101_1_101000101011;
      patterns[17790] = 29'b0_100010101111_110_0_100010101111;
      patterns[17791] = 29'b0_100010101111_111_0_100010101111;
      patterns[17792] = 29'b0_100010110000_000_0_100010110000;
      patterns[17793] = 29'b0_100010110000_001_0_110000100010;
      patterns[17794] = 29'b0_100010110000_010_1_000101100000;
      patterns[17795] = 29'b0_100010110000_011_0_001011000001;
      patterns[17796] = 29'b0_100010110000_100_0_010001011000;
      patterns[17797] = 29'b0_100010110000_101_0_001000101100;
      patterns[17798] = 29'b0_100010110000_110_0_100010110000;
      patterns[17799] = 29'b0_100010110000_111_0_100010110000;
      patterns[17800] = 29'b0_100010110001_000_0_100010110001;
      patterns[17801] = 29'b0_100010110001_001_0_110001100010;
      patterns[17802] = 29'b0_100010110001_010_1_000101100010;
      patterns[17803] = 29'b0_100010110001_011_0_001011000101;
      patterns[17804] = 29'b0_100010110001_100_1_010001011000;
      patterns[17805] = 29'b0_100010110001_101_0_101000101100;
      patterns[17806] = 29'b0_100010110001_110_0_100010110001;
      patterns[17807] = 29'b0_100010110001_111_0_100010110001;
      patterns[17808] = 29'b0_100010110010_000_0_100010110010;
      patterns[17809] = 29'b0_100010110010_001_0_110010100010;
      patterns[17810] = 29'b0_100010110010_010_1_000101100100;
      patterns[17811] = 29'b0_100010110010_011_0_001011001001;
      patterns[17812] = 29'b0_100010110010_100_0_010001011001;
      patterns[17813] = 29'b0_100010110010_101_1_001000101100;
      patterns[17814] = 29'b0_100010110010_110_0_100010110010;
      patterns[17815] = 29'b0_100010110010_111_0_100010110010;
      patterns[17816] = 29'b0_100010110011_000_0_100010110011;
      patterns[17817] = 29'b0_100010110011_001_0_110011100010;
      patterns[17818] = 29'b0_100010110011_010_1_000101100110;
      patterns[17819] = 29'b0_100010110011_011_0_001011001101;
      patterns[17820] = 29'b0_100010110011_100_1_010001011001;
      patterns[17821] = 29'b0_100010110011_101_1_101000101100;
      patterns[17822] = 29'b0_100010110011_110_0_100010110011;
      patterns[17823] = 29'b0_100010110011_111_0_100010110011;
      patterns[17824] = 29'b0_100010110100_000_0_100010110100;
      patterns[17825] = 29'b0_100010110100_001_0_110100100010;
      patterns[17826] = 29'b0_100010110100_010_1_000101101000;
      patterns[17827] = 29'b0_100010110100_011_0_001011010001;
      patterns[17828] = 29'b0_100010110100_100_0_010001011010;
      patterns[17829] = 29'b0_100010110100_101_0_001000101101;
      patterns[17830] = 29'b0_100010110100_110_0_100010110100;
      patterns[17831] = 29'b0_100010110100_111_0_100010110100;
      patterns[17832] = 29'b0_100010110101_000_0_100010110101;
      patterns[17833] = 29'b0_100010110101_001_0_110101100010;
      patterns[17834] = 29'b0_100010110101_010_1_000101101010;
      patterns[17835] = 29'b0_100010110101_011_0_001011010101;
      patterns[17836] = 29'b0_100010110101_100_1_010001011010;
      patterns[17837] = 29'b0_100010110101_101_0_101000101101;
      patterns[17838] = 29'b0_100010110101_110_0_100010110101;
      patterns[17839] = 29'b0_100010110101_111_0_100010110101;
      patterns[17840] = 29'b0_100010110110_000_0_100010110110;
      patterns[17841] = 29'b0_100010110110_001_0_110110100010;
      patterns[17842] = 29'b0_100010110110_010_1_000101101100;
      patterns[17843] = 29'b0_100010110110_011_0_001011011001;
      patterns[17844] = 29'b0_100010110110_100_0_010001011011;
      patterns[17845] = 29'b0_100010110110_101_1_001000101101;
      patterns[17846] = 29'b0_100010110110_110_0_100010110110;
      patterns[17847] = 29'b0_100010110110_111_0_100010110110;
      patterns[17848] = 29'b0_100010110111_000_0_100010110111;
      patterns[17849] = 29'b0_100010110111_001_0_110111100010;
      patterns[17850] = 29'b0_100010110111_010_1_000101101110;
      patterns[17851] = 29'b0_100010110111_011_0_001011011101;
      patterns[17852] = 29'b0_100010110111_100_1_010001011011;
      patterns[17853] = 29'b0_100010110111_101_1_101000101101;
      patterns[17854] = 29'b0_100010110111_110_0_100010110111;
      patterns[17855] = 29'b0_100010110111_111_0_100010110111;
      patterns[17856] = 29'b0_100010111000_000_0_100010111000;
      patterns[17857] = 29'b0_100010111000_001_0_111000100010;
      patterns[17858] = 29'b0_100010111000_010_1_000101110000;
      patterns[17859] = 29'b0_100010111000_011_0_001011100001;
      patterns[17860] = 29'b0_100010111000_100_0_010001011100;
      patterns[17861] = 29'b0_100010111000_101_0_001000101110;
      patterns[17862] = 29'b0_100010111000_110_0_100010111000;
      patterns[17863] = 29'b0_100010111000_111_0_100010111000;
      patterns[17864] = 29'b0_100010111001_000_0_100010111001;
      patterns[17865] = 29'b0_100010111001_001_0_111001100010;
      patterns[17866] = 29'b0_100010111001_010_1_000101110010;
      patterns[17867] = 29'b0_100010111001_011_0_001011100101;
      patterns[17868] = 29'b0_100010111001_100_1_010001011100;
      patterns[17869] = 29'b0_100010111001_101_0_101000101110;
      patterns[17870] = 29'b0_100010111001_110_0_100010111001;
      patterns[17871] = 29'b0_100010111001_111_0_100010111001;
      patterns[17872] = 29'b0_100010111010_000_0_100010111010;
      patterns[17873] = 29'b0_100010111010_001_0_111010100010;
      patterns[17874] = 29'b0_100010111010_010_1_000101110100;
      patterns[17875] = 29'b0_100010111010_011_0_001011101001;
      patterns[17876] = 29'b0_100010111010_100_0_010001011101;
      patterns[17877] = 29'b0_100010111010_101_1_001000101110;
      patterns[17878] = 29'b0_100010111010_110_0_100010111010;
      patterns[17879] = 29'b0_100010111010_111_0_100010111010;
      patterns[17880] = 29'b0_100010111011_000_0_100010111011;
      patterns[17881] = 29'b0_100010111011_001_0_111011100010;
      patterns[17882] = 29'b0_100010111011_010_1_000101110110;
      patterns[17883] = 29'b0_100010111011_011_0_001011101101;
      patterns[17884] = 29'b0_100010111011_100_1_010001011101;
      patterns[17885] = 29'b0_100010111011_101_1_101000101110;
      patterns[17886] = 29'b0_100010111011_110_0_100010111011;
      patterns[17887] = 29'b0_100010111011_111_0_100010111011;
      patterns[17888] = 29'b0_100010111100_000_0_100010111100;
      patterns[17889] = 29'b0_100010111100_001_0_111100100010;
      patterns[17890] = 29'b0_100010111100_010_1_000101111000;
      patterns[17891] = 29'b0_100010111100_011_0_001011110001;
      patterns[17892] = 29'b0_100010111100_100_0_010001011110;
      patterns[17893] = 29'b0_100010111100_101_0_001000101111;
      patterns[17894] = 29'b0_100010111100_110_0_100010111100;
      patterns[17895] = 29'b0_100010111100_111_0_100010111100;
      patterns[17896] = 29'b0_100010111101_000_0_100010111101;
      patterns[17897] = 29'b0_100010111101_001_0_111101100010;
      patterns[17898] = 29'b0_100010111101_010_1_000101111010;
      patterns[17899] = 29'b0_100010111101_011_0_001011110101;
      patterns[17900] = 29'b0_100010111101_100_1_010001011110;
      patterns[17901] = 29'b0_100010111101_101_0_101000101111;
      patterns[17902] = 29'b0_100010111101_110_0_100010111101;
      patterns[17903] = 29'b0_100010111101_111_0_100010111101;
      patterns[17904] = 29'b0_100010111110_000_0_100010111110;
      patterns[17905] = 29'b0_100010111110_001_0_111110100010;
      patterns[17906] = 29'b0_100010111110_010_1_000101111100;
      patterns[17907] = 29'b0_100010111110_011_0_001011111001;
      patterns[17908] = 29'b0_100010111110_100_0_010001011111;
      patterns[17909] = 29'b0_100010111110_101_1_001000101111;
      patterns[17910] = 29'b0_100010111110_110_0_100010111110;
      patterns[17911] = 29'b0_100010111110_111_0_100010111110;
      patterns[17912] = 29'b0_100010111111_000_0_100010111111;
      patterns[17913] = 29'b0_100010111111_001_0_111111100010;
      patterns[17914] = 29'b0_100010111111_010_1_000101111110;
      patterns[17915] = 29'b0_100010111111_011_0_001011111101;
      patterns[17916] = 29'b0_100010111111_100_1_010001011111;
      patterns[17917] = 29'b0_100010111111_101_1_101000101111;
      patterns[17918] = 29'b0_100010111111_110_0_100010111111;
      patterns[17919] = 29'b0_100010111111_111_0_100010111111;
      patterns[17920] = 29'b0_100011000000_000_0_100011000000;
      patterns[17921] = 29'b0_100011000000_001_0_000000100011;
      patterns[17922] = 29'b0_100011000000_010_1_000110000000;
      patterns[17923] = 29'b0_100011000000_011_0_001100000001;
      patterns[17924] = 29'b0_100011000000_100_0_010001100000;
      patterns[17925] = 29'b0_100011000000_101_0_001000110000;
      patterns[17926] = 29'b0_100011000000_110_0_100011000000;
      patterns[17927] = 29'b0_100011000000_111_0_100011000000;
      patterns[17928] = 29'b0_100011000001_000_0_100011000001;
      patterns[17929] = 29'b0_100011000001_001_0_000001100011;
      patterns[17930] = 29'b0_100011000001_010_1_000110000010;
      patterns[17931] = 29'b0_100011000001_011_0_001100000101;
      patterns[17932] = 29'b0_100011000001_100_1_010001100000;
      patterns[17933] = 29'b0_100011000001_101_0_101000110000;
      patterns[17934] = 29'b0_100011000001_110_0_100011000001;
      patterns[17935] = 29'b0_100011000001_111_0_100011000001;
      patterns[17936] = 29'b0_100011000010_000_0_100011000010;
      patterns[17937] = 29'b0_100011000010_001_0_000010100011;
      patterns[17938] = 29'b0_100011000010_010_1_000110000100;
      patterns[17939] = 29'b0_100011000010_011_0_001100001001;
      patterns[17940] = 29'b0_100011000010_100_0_010001100001;
      patterns[17941] = 29'b0_100011000010_101_1_001000110000;
      patterns[17942] = 29'b0_100011000010_110_0_100011000010;
      patterns[17943] = 29'b0_100011000010_111_0_100011000010;
      patterns[17944] = 29'b0_100011000011_000_0_100011000011;
      patterns[17945] = 29'b0_100011000011_001_0_000011100011;
      patterns[17946] = 29'b0_100011000011_010_1_000110000110;
      patterns[17947] = 29'b0_100011000011_011_0_001100001101;
      patterns[17948] = 29'b0_100011000011_100_1_010001100001;
      patterns[17949] = 29'b0_100011000011_101_1_101000110000;
      patterns[17950] = 29'b0_100011000011_110_0_100011000011;
      patterns[17951] = 29'b0_100011000011_111_0_100011000011;
      patterns[17952] = 29'b0_100011000100_000_0_100011000100;
      patterns[17953] = 29'b0_100011000100_001_0_000100100011;
      patterns[17954] = 29'b0_100011000100_010_1_000110001000;
      patterns[17955] = 29'b0_100011000100_011_0_001100010001;
      patterns[17956] = 29'b0_100011000100_100_0_010001100010;
      patterns[17957] = 29'b0_100011000100_101_0_001000110001;
      patterns[17958] = 29'b0_100011000100_110_0_100011000100;
      patterns[17959] = 29'b0_100011000100_111_0_100011000100;
      patterns[17960] = 29'b0_100011000101_000_0_100011000101;
      patterns[17961] = 29'b0_100011000101_001_0_000101100011;
      patterns[17962] = 29'b0_100011000101_010_1_000110001010;
      patterns[17963] = 29'b0_100011000101_011_0_001100010101;
      patterns[17964] = 29'b0_100011000101_100_1_010001100010;
      patterns[17965] = 29'b0_100011000101_101_0_101000110001;
      patterns[17966] = 29'b0_100011000101_110_0_100011000101;
      patterns[17967] = 29'b0_100011000101_111_0_100011000101;
      patterns[17968] = 29'b0_100011000110_000_0_100011000110;
      patterns[17969] = 29'b0_100011000110_001_0_000110100011;
      patterns[17970] = 29'b0_100011000110_010_1_000110001100;
      patterns[17971] = 29'b0_100011000110_011_0_001100011001;
      patterns[17972] = 29'b0_100011000110_100_0_010001100011;
      patterns[17973] = 29'b0_100011000110_101_1_001000110001;
      patterns[17974] = 29'b0_100011000110_110_0_100011000110;
      patterns[17975] = 29'b0_100011000110_111_0_100011000110;
      patterns[17976] = 29'b0_100011000111_000_0_100011000111;
      patterns[17977] = 29'b0_100011000111_001_0_000111100011;
      patterns[17978] = 29'b0_100011000111_010_1_000110001110;
      patterns[17979] = 29'b0_100011000111_011_0_001100011101;
      patterns[17980] = 29'b0_100011000111_100_1_010001100011;
      patterns[17981] = 29'b0_100011000111_101_1_101000110001;
      patterns[17982] = 29'b0_100011000111_110_0_100011000111;
      patterns[17983] = 29'b0_100011000111_111_0_100011000111;
      patterns[17984] = 29'b0_100011001000_000_0_100011001000;
      patterns[17985] = 29'b0_100011001000_001_0_001000100011;
      patterns[17986] = 29'b0_100011001000_010_1_000110010000;
      patterns[17987] = 29'b0_100011001000_011_0_001100100001;
      patterns[17988] = 29'b0_100011001000_100_0_010001100100;
      patterns[17989] = 29'b0_100011001000_101_0_001000110010;
      patterns[17990] = 29'b0_100011001000_110_0_100011001000;
      patterns[17991] = 29'b0_100011001000_111_0_100011001000;
      patterns[17992] = 29'b0_100011001001_000_0_100011001001;
      patterns[17993] = 29'b0_100011001001_001_0_001001100011;
      patterns[17994] = 29'b0_100011001001_010_1_000110010010;
      patterns[17995] = 29'b0_100011001001_011_0_001100100101;
      patterns[17996] = 29'b0_100011001001_100_1_010001100100;
      patterns[17997] = 29'b0_100011001001_101_0_101000110010;
      patterns[17998] = 29'b0_100011001001_110_0_100011001001;
      patterns[17999] = 29'b0_100011001001_111_0_100011001001;
      patterns[18000] = 29'b0_100011001010_000_0_100011001010;
      patterns[18001] = 29'b0_100011001010_001_0_001010100011;
      patterns[18002] = 29'b0_100011001010_010_1_000110010100;
      patterns[18003] = 29'b0_100011001010_011_0_001100101001;
      patterns[18004] = 29'b0_100011001010_100_0_010001100101;
      patterns[18005] = 29'b0_100011001010_101_1_001000110010;
      patterns[18006] = 29'b0_100011001010_110_0_100011001010;
      patterns[18007] = 29'b0_100011001010_111_0_100011001010;
      patterns[18008] = 29'b0_100011001011_000_0_100011001011;
      patterns[18009] = 29'b0_100011001011_001_0_001011100011;
      patterns[18010] = 29'b0_100011001011_010_1_000110010110;
      patterns[18011] = 29'b0_100011001011_011_0_001100101101;
      patterns[18012] = 29'b0_100011001011_100_1_010001100101;
      patterns[18013] = 29'b0_100011001011_101_1_101000110010;
      patterns[18014] = 29'b0_100011001011_110_0_100011001011;
      patterns[18015] = 29'b0_100011001011_111_0_100011001011;
      patterns[18016] = 29'b0_100011001100_000_0_100011001100;
      patterns[18017] = 29'b0_100011001100_001_0_001100100011;
      patterns[18018] = 29'b0_100011001100_010_1_000110011000;
      patterns[18019] = 29'b0_100011001100_011_0_001100110001;
      patterns[18020] = 29'b0_100011001100_100_0_010001100110;
      patterns[18021] = 29'b0_100011001100_101_0_001000110011;
      patterns[18022] = 29'b0_100011001100_110_0_100011001100;
      patterns[18023] = 29'b0_100011001100_111_0_100011001100;
      patterns[18024] = 29'b0_100011001101_000_0_100011001101;
      patterns[18025] = 29'b0_100011001101_001_0_001101100011;
      patterns[18026] = 29'b0_100011001101_010_1_000110011010;
      patterns[18027] = 29'b0_100011001101_011_0_001100110101;
      patterns[18028] = 29'b0_100011001101_100_1_010001100110;
      patterns[18029] = 29'b0_100011001101_101_0_101000110011;
      patterns[18030] = 29'b0_100011001101_110_0_100011001101;
      patterns[18031] = 29'b0_100011001101_111_0_100011001101;
      patterns[18032] = 29'b0_100011001110_000_0_100011001110;
      patterns[18033] = 29'b0_100011001110_001_0_001110100011;
      patterns[18034] = 29'b0_100011001110_010_1_000110011100;
      patterns[18035] = 29'b0_100011001110_011_0_001100111001;
      patterns[18036] = 29'b0_100011001110_100_0_010001100111;
      patterns[18037] = 29'b0_100011001110_101_1_001000110011;
      patterns[18038] = 29'b0_100011001110_110_0_100011001110;
      patterns[18039] = 29'b0_100011001110_111_0_100011001110;
      patterns[18040] = 29'b0_100011001111_000_0_100011001111;
      patterns[18041] = 29'b0_100011001111_001_0_001111100011;
      patterns[18042] = 29'b0_100011001111_010_1_000110011110;
      patterns[18043] = 29'b0_100011001111_011_0_001100111101;
      patterns[18044] = 29'b0_100011001111_100_1_010001100111;
      patterns[18045] = 29'b0_100011001111_101_1_101000110011;
      patterns[18046] = 29'b0_100011001111_110_0_100011001111;
      patterns[18047] = 29'b0_100011001111_111_0_100011001111;
      patterns[18048] = 29'b0_100011010000_000_0_100011010000;
      patterns[18049] = 29'b0_100011010000_001_0_010000100011;
      patterns[18050] = 29'b0_100011010000_010_1_000110100000;
      patterns[18051] = 29'b0_100011010000_011_0_001101000001;
      patterns[18052] = 29'b0_100011010000_100_0_010001101000;
      patterns[18053] = 29'b0_100011010000_101_0_001000110100;
      patterns[18054] = 29'b0_100011010000_110_0_100011010000;
      patterns[18055] = 29'b0_100011010000_111_0_100011010000;
      patterns[18056] = 29'b0_100011010001_000_0_100011010001;
      patterns[18057] = 29'b0_100011010001_001_0_010001100011;
      patterns[18058] = 29'b0_100011010001_010_1_000110100010;
      patterns[18059] = 29'b0_100011010001_011_0_001101000101;
      patterns[18060] = 29'b0_100011010001_100_1_010001101000;
      patterns[18061] = 29'b0_100011010001_101_0_101000110100;
      patterns[18062] = 29'b0_100011010001_110_0_100011010001;
      patterns[18063] = 29'b0_100011010001_111_0_100011010001;
      patterns[18064] = 29'b0_100011010010_000_0_100011010010;
      patterns[18065] = 29'b0_100011010010_001_0_010010100011;
      patterns[18066] = 29'b0_100011010010_010_1_000110100100;
      patterns[18067] = 29'b0_100011010010_011_0_001101001001;
      patterns[18068] = 29'b0_100011010010_100_0_010001101001;
      patterns[18069] = 29'b0_100011010010_101_1_001000110100;
      patterns[18070] = 29'b0_100011010010_110_0_100011010010;
      patterns[18071] = 29'b0_100011010010_111_0_100011010010;
      patterns[18072] = 29'b0_100011010011_000_0_100011010011;
      patterns[18073] = 29'b0_100011010011_001_0_010011100011;
      patterns[18074] = 29'b0_100011010011_010_1_000110100110;
      patterns[18075] = 29'b0_100011010011_011_0_001101001101;
      patterns[18076] = 29'b0_100011010011_100_1_010001101001;
      patterns[18077] = 29'b0_100011010011_101_1_101000110100;
      patterns[18078] = 29'b0_100011010011_110_0_100011010011;
      patterns[18079] = 29'b0_100011010011_111_0_100011010011;
      patterns[18080] = 29'b0_100011010100_000_0_100011010100;
      patterns[18081] = 29'b0_100011010100_001_0_010100100011;
      patterns[18082] = 29'b0_100011010100_010_1_000110101000;
      patterns[18083] = 29'b0_100011010100_011_0_001101010001;
      patterns[18084] = 29'b0_100011010100_100_0_010001101010;
      patterns[18085] = 29'b0_100011010100_101_0_001000110101;
      patterns[18086] = 29'b0_100011010100_110_0_100011010100;
      patterns[18087] = 29'b0_100011010100_111_0_100011010100;
      patterns[18088] = 29'b0_100011010101_000_0_100011010101;
      patterns[18089] = 29'b0_100011010101_001_0_010101100011;
      patterns[18090] = 29'b0_100011010101_010_1_000110101010;
      patterns[18091] = 29'b0_100011010101_011_0_001101010101;
      patterns[18092] = 29'b0_100011010101_100_1_010001101010;
      patterns[18093] = 29'b0_100011010101_101_0_101000110101;
      patterns[18094] = 29'b0_100011010101_110_0_100011010101;
      patterns[18095] = 29'b0_100011010101_111_0_100011010101;
      patterns[18096] = 29'b0_100011010110_000_0_100011010110;
      patterns[18097] = 29'b0_100011010110_001_0_010110100011;
      patterns[18098] = 29'b0_100011010110_010_1_000110101100;
      patterns[18099] = 29'b0_100011010110_011_0_001101011001;
      patterns[18100] = 29'b0_100011010110_100_0_010001101011;
      patterns[18101] = 29'b0_100011010110_101_1_001000110101;
      patterns[18102] = 29'b0_100011010110_110_0_100011010110;
      patterns[18103] = 29'b0_100011010110_111_0_100011010110;
      patterns[18104] = 29'b0_100011010111_000_0_100011010111;
      patterns[18105] = 29'b0_100011010111_001_0_010111100011;
      patterns[18106] = 29'b0_100011010111_010_1_000110101110;
      patterns[18107] = 29'b0_100011010111_011_0_001101011101;
      patterns[18108] = 29'b0_100011010111_100_1_010001101011;
      patterns[18109] = 29'b0_100011010111_101_1_101000110101;
      patterns[18110] = 29'b0_100011010111_110_0_100011010111;
      patterns[18111] = 29'b0_100011010111_111_0_100011010111;
      patterns[18112] = 29'b0_100011011000_000_0_100011011000;
      patterns[18113] = 29'b0_100011011000_001_0_011000100011;
      patterns[18114] = 29'b0_100011011000_010_1_000110110000;
      patterns[18115] = 29'b0_100011011000_011_0_001101100001;
      patterns[18116] = 29'b0_100011011000_100_0_010001101100;
      patterns[18117] = 29'b0_100011011000_101_0_001000110110;
      patterns[18118] = 29'b0_100011011000_110_0_100011011000;
      patterns[18119] = 29'b0_100011011000_111_0_100011011000;
      patterns[18120] = 29'b0_100011011001_000_0_100011011001;
      patterns[18121] = 29'b0_100011011001_001_0_011001100011;
      patterns[18122] = 29'b0_100011011001_010_1_000110110010;
      patterns[18123] = 29'b0_100011011001_011_0_001101100101;
      patterns[18124] = 29'b0_100011011001_100_1_010001101100;
      patterns[18125] = 29'b0_100011011001_101_0_101000110110;
      patterns[18126] = 29'b0_100011011001_110_0_100011011001;
      patterns[18127] = 29'b0_100011011001_111_0_100011011001;
      patterns[18128] = 29'b0_100011011010_000_0_100011011010;
      patterns[18129] = 29'b0_100011011010_001_0_011010100011;
      patterns[18130] = 29'b0_100011011010_010_1_000110110100;
      patterns[18131] = 29'b0_100011011010_011_0_001101101001;
      patterns[18132] = 29'b0_100011011010_100_0_010001101101;
      patterns[18133] = 29'b0_100011011010_101_1_001000110110;
      patterns[18134] = 29'b0_100011011010_110_0_100011011010;
      patterns[18135] = 29'b0_100011011010_111_0_100011011010;
      patterns[18136] = 29'b0_100011011011_000_0_100011011011;
      patterns[18137] = 29'b0_100011011011_001_0_011011100011;
      patterns[18138] = 29'b0_100011011011_010_1_000110110110;
      patterns[18139] = 29'b0_100011011011_011_0_001101101101;
      patterns[18140] = 29'b0_100011011011_100_1_010001101101;
      patterns[18141] = 29'b0_100011011011_101_1_101000110110;
      patterns[18142] = 29'b0_100011011011_110_0_100011011011;
      patterns[18143] = 29'b0_100011011011_111_0_100011011011;
      patterns[18144] = 29'b0_100011011100_000_0_100011011100;
      patterns[18145] = 29'b0_100011011100_001_0_011100100011;
      patterns[18146] = 29'b0_100011011100_010_1_000110111000;
      patterns[18147] = 29'b0_100011011100_011_0_001101110001;
      patterns[18148] = 29'b0_100011011100_100_0_010001101110;
      patterns[18149] = 29'b0_100011011100_101_0_001000110111;
      patterns[18150] = 29'b0_100011011100_110_0_100011011100;
      patterns[18151] = 29'b0_100011011100_111_0_100011011100;
      patterns[18152] = 29'b0_100011011101_000_0_100011011101;
      patterns[18153] = 29'b0_100011011101_001_0_011101100011;
      patterns[18154] = 29'b0_100011011101_010_1_000110111010;
      patterns[18155] = 29'b0_100011011101_011_0_001101110101;
      patterns[18156] = 29'b0_100011011101_100_1_010001101110;
      patterns[18157] = 29'b0_100011011101_101_0_101000110111;
      patterns[18158] = 29'b0_100011011101_110_0_100011011101;
      patterns[18159] = 29'b0_100011011101_111_0_100011011101;
      patterns[18160] = 29'b0_100011011110_000_0_100011011110;
      patterns[18161] = 29'b0_100011011110_001_0_011110100011;
      patterns[18162] = 29'b0_100011011110_010_1_000110111100;
      patterns[18163] = 29'b0_100011011110_011_0_001101111001;
      patterns[18164] = 29'b0_100011011110_100_0_010001101111;
      patterns[18165] = 29'b0_100011011110_101_1_001000110111;
      patterns[18166] = 29'b0_100011011110_110_0_100011011110;
      patterns[18167] = 29'b0_100011011110_111_0_100011011110;
      patterns[18168] = 29'b0_100011011111_000_0_100011011111;
      patterns[18169] = 29'b0_100011011111_001_0_011111100011;
      patterns[18170] = 29'b0_100011011111_010_1_000110111110;
      patterns[18171] = 29'b0_100011011111_011_0_001101111101;
      patterns[18172] = 29'b0_100011011111_100_1_010001101111;
      patterns[18173] = 29'b0_100011011111_101_1_101000110111;
      patterns[18174] = 29'b0_100011011111_110_0_100011011111;
      patterns[18175] = 29'b0_100011011111_111_0_100011011111;
      patterns[18176] = 29'b0_100011100000_000_0_100011100000;
      patterns[18177] = 29'b0_100011100000_001_0_100000100011;
      patterns[18178] = 29'b0_100011100000_010_1_000111000000;
      patterns[18179] = 29'b0_100011100000_011_0_001110000001;
      patterns[18180] = 29'b0_100011100000_100_0_010001110000;
      patterns[18181] = 29'b0_100011100000_101_0_001000111000;
      patterns[18182] = 29'b0_100011100000_110_0_100011100000;
      patterns[18183] = 29'b0_100011100000_111_0_100011100000;
      patterns[18184] = 29'b0_100011100001_000_0_100011100001;
      patterns[18185] = 29'b0_100011100001_001_0_100001100011;
      patterns[18186] = 29'b0_100011100001_010_1_000111000010;
      patterns[18187] = 29'b0_100011100001_011_0_001110000101;
      patterns[18188] = 29'b0_100011100001_100_1_010001110000;
      patterns[18189] = 29'b0_100011100001_101_0_101000111000;
      patterns[18190] = 29'b0_100011100001_110_0_100011100001;
      patterns[18191] = 29'b0_100011100001_111_0_100011100001;
      patterns[18192] = 29'b0_100011100010_000_0_100011100010;
      patterns[18193] = 29'b0_100011100010_001_0_100010100011;
      patterns[18194] = 29'b0_100011100010_010_1_000111000100;
      patterns[18195] = 29'b0_100011100010_011_0_001110001001;
      patterns[18196] = 29'b0_100011100010_100_0_010001110001;
      patterns[18197] = 29'b0_100011100010_101_1_001000111000;
      patterns[18198] = 29'b0_100011100010_110_0_100011100010;
      patterns[18199] = 29'b0_100011100010_111_0_100011100010;
      patterns[18200] = 29'b0_100011100011_000_0_100011100011;
      patterns[18201] = 29'b0_100011100011_001_0_100011100011;
      patterns[18202] = 29'b0_100011100011_010_1_000111000110;
      patterns[18203] = 29'b0_100011100011_011_0_001110001101;
      patterns[18204] = 29'b0_100011100011_100_1_010001110001;
      patterns[18205] = 29'b0_100011100011_101_1_101000111000;
      patterns[18206] = 29'b0_100011100011_110_0_100011100011;
      patterns[18207] = 29'b0_100011100011_111_0_100011100011;
      patterns[18208] = 29'b0_100011100100_000_0_100011100100;
      patterns[18209] = 29'b0_100011100100_001_0_100100100011;
      patterns[18210] = 29'b0_100011100100_010_1_000111001000;
      patterns[18211] = 29'b0_100011100100_011_0_001110010001;
      patterns[18212] = 29'b0_100011100100_100_0_010001110010;
      patterns[18213] = 29'b0_100011100100_101_0_001000111001;
      patterns[18214] = 29'b0_100011100100_110_0_100011100100;
      patterns[18215] = 29'b0_100011100100_111_0_100011100100;
      patterns[18216] = 29'b0_100011100101_000_0_100011100101;
      patterns[18217] = 29'b0_100011100101_001_0_100101100011;
      patterns[18218] = 29'b0_100011100101_010_1_000111001010;
      patterns[18219] = 29'b0_100011100101_011_0_001110010101;
      patterns[18220] = 29'b0_100011100101_100_1_010001110010;
      patterns[18221] = 29'b0_100011100101_101_0_101000111001;
      patterns[18222] = 29'b0_100011100101_110_0_100011100101;
      patterns[18223] = 29'b0_100011100101_111_0_100011100101;
      patterns[18224] = 29'b0_100011100110_000_0_100011100110;
      patterns[18225] = 29'b0_100011100110_001_0_100110100011;
      patterns[18226] = 29'b0_100011100110_010_1_000111001100;
      patterns[18227] = 29'b0_100011100110_011_0_001110011001;
      patterns[18228] = 29'b0_100011100110_100_0_010001110011;
      patterns[18229] = 29'b0_100011100110_101_1_001000111001;
      patterns[18230] = 29'b0_100011100110_110_0_100011100110;
      patterns[18231] = 29'b0_100011100110_111_0_100011100110;
      patterns[18232] = 29'b0_100011100111_000_0_100011100111;
      patterns[18233] = 29'b0_100011100111_001_0_100111100011;
      patterns[18234] = 29'b0_100011100111_010_1_000111001110;
      patterns[18235] = 29'b0_100011100111_011_0_001110011101;
      patterns[18236] = 29'b0_100011100111_100_1_010001110011;
      patterns[18237] = 29'b0_100011100111_101_1_101000111001;
      patterns[18238] = 29'b0_100011100111_110_0_100011100111;
      patterns[18239] = 29'b0_100011100111_111_0_100011100111;
      patterns[18240] = 29'b0_100011101000_000_0_100011101000;
      patterns[18241] = 29'b0_100011101000_001_0_101000100011;
      patterns[18242] = 29'b0_100011101000_010_1_000111010000;
      patterns[18243] = 29'b0_100011101000_011_0_001110100001;
      patterns[18244] = 29'b0_100011101000_100_0_010001110100;
      patterns[18245] = 29'b0_100011101000_101_0_001000111010;
      patterns[18246] = 29'b0_100011101000_110_0_100011101000;
      patterns[18247] = 29'b0_100011101000_111_0_100011101000;
      patterns[18248] = 29'b0_100011101001_000_0_100011101001;
      patterns[18249] = 29'b0_100011101001_001_0_101001100011;
      patterns[18250] = 29'b0_100011101001_010_1_000111010010;
      patterns[18251] = 29'b0_100011101001_011_0_001110100101;
      patterns[18252] = 29'b0_100011101001_100_1_010001110100;
      patterns[18253] = 29'b0_100011101001_101_0_101000111010;
      patterns[18254] = 29'b0_100011101001_110_0_100011101001;
      patterns[18255] = 29'b0_100011101001_111_0_100011101001;
      patterns[18256] = 29'b0_100011101010_000_0_100011101010;
      patterns[18257] = 29'b0_100011101010_001_0_101010100011;
      patterns[18258] = 29'b0_100011101010_010_1_000111010100;
      patterns[18259] = 29'b0_100011101010_011_0_001110101001;
      patterns[18260] = 29'b0_100011101010_100_0_010001110101;
      patterns[18261] = 29'b0_100011101010_101_1_001000111010;
      patterns[18262] = 29'b0_100011101010_110_0_100011101010;
      patterns[18263] = 29'b0_100011101010_111_0_100011101010;
      patterns[18264] = 29'b0_100011101011_000_0_100011101011;
      patterns[18265] = 29'b0_100011101011_001_0_101011100011;
      patterns[18266] = 29'b0_100011101011_010_1_000111010110;
      patterns[18267] = 29'b0_100011101011_011_0_001110101101;
      patterns[18268] = 29'b0_100011101011_100_1_010001110101;
      patterns[18269] = 29'b0_100011101011_101_1_101000111010;
      patterns[18270] = 29'b0_100011101011_110_0_100011101011;
      patterns[18271] = 29'b0_100011101011_111_0_100011101011;
      patterns[18272] = 29'b0_100011101100_000_0_100011101100;
      patterns[18273] = 29'b0_100011101100_001_0_101100100011;
      patterns[18274] = 29'b0_100011101100_010_1_000111011000;
      patterns[18275] = 29'b0_100011101100_011_0_001110110001;
      patterns[18276] = 29'b0_100011101100_100_0_010001110110;
      patterns[18277] = 29'b0_100011101100_101_0_001000111011;
      patterns[18278] = 29'b0_100011101100_110_0_100011101100;
      patterns[18279] = 29'b0_100011101100_111_0_100011101100;
      patterns[18280] = 29'b0_100011101101_000_0_100011101101;
      patterns[18281] = 29'b0_100011101101_001_0_101101100011;
      patterns[18282] = 29'b0_100011101101_010_1_000111011010;
      patterns[18283] = 29'b0_100011101101_011_0_001110110101;
      patterns[18284] = 29'b0_100011101101_100_1_010001110110;
      patterns[18285] = 29'b0_100011101101_101_0_101000111011;
      patterns[18286] = 29'b0_100011101101_110_0_100011101101;
      patterns[18287] = 29'b0_100011101101_111_0_100011101101;
      patterns[18288] = 29'b0_100011101110_000_0_100011101110;
      patterns[18289] = 29'b0_100011101110_001_0_101110100011;
      patterns[18290] = 29'b0_100011101110_010_1_000111011100;
      patterns[18291] = 29'b0_100011101110_011_0_001110111001;
      patterns[18292] = 29'b0_100011101110_100_0_010001110111;
      patterns[18293] = 29'b0_100011101110_101_1_001000111011;
      patterns[18294] = 29'b0_100011101110_110_0_100011101110;
      patterns[18295] = 29'b0_100011101110_111_0_100011101110;
      patterns[18296] = 29'b0_100011101111_000_0_100011101111;
      patterns[18297] = 29'b0_100011101111_001_0_101111100011;
      patterns[18298] = 29'b0_100011101111_010_1_000111011110;
      patterns[18299] = 29'b0_100011101111_011_0_001110111101;
      patterns[18300] = 29'b0_100011101111_100_1_010001110111;
      patterns[18301] = 29'b0_100011101111_101_1_101000111011;
      patterns[18302] = 29'b0_100011101111_110_0_100011101111;
      patterns[18303] = 29'b0_100011101111_111_0_100011101111;
      patterns[18304] = 29'b0_100011110000_000_0_100011110000;
      patterns[18305] = 29'b0_100011110000_001_0_110000100011;
      patterns[18306] = 29'b0_100011110000_010_1_000111100000;
      patterns[18307] = 29'b0_100011110000_011_0_001111000001;
      patterns[18308] = 29'b0_100011110000_100_0_010001111000;
      patterns[18309] = 29'b0_100011110000_101_0_001000111100;
      patterns[18310] = 29'b0_100011110000_110_0_100011110000;
      patterns[18311] = 29'b0_100011110000_111_0_100011110000;
      patterns[18312] = 29'b0_100011110001_000_0_100011110001;
      patterns[18313] = 29'b0_100011110001_001_0_110001100011;
      patterns[18314] = 29'b0_100011110001_010_1_000111100010;
      patterns[18315] = 29'b0_100011110001_011_0_001111000101;
      patterns[18316] = 29'b0_100011110001_100_1_010001111000;
      patterns[18317] = 29'b0_100011110001_101_0_101000111100;
      patterns[18318] = 29'b0_100011110001_110_0_100011110001;
      patterns[18319] = 29'b0_100011110001_111_0_100011110001;
      patterns[18320] = 29'b0_100011110010_000_0_100011110010;
      patterns[18321] = 29'b0_100011110010_001_0_110010100011;
      patterns[18322] = 29'b0_100011110010_010_1_000111100100;
      patterns[18323] = 29'b0_100011110010_011_0_001111001001;
      patterns[18324] = 29'b0_100011110010_100_0_010001111001;
      patterns[18325] = 29'b0_100011110010_101_1_001000111100;
      patterns[18326] = 29'b0_100011110010_110_0_100011110010;
      patterns[18327] = 29'b0_100011110010_111_0_100011110010;
      patterns[18328] = 29'b0_100011110011_000_0_100011110011;
      patterns[18329] = 29'b0_100011110011_001_0_110011100011;
      patterns[18330] = 29'b0_100011110011_010_1_000111100110;
      patterns[18331] = 29'b0_100011110011_011_0_001111001101;
      patterns[18332] = 29'b0_100011110011_100_1_010001111001;
      patterns[18333] = 29'b0_100011110011_101_1_101000111100;
      patterns[18334] = 29'b0_100011110011_110_0_100011110011;
      patterns[18335] = 29'b0_100011110011_111_0_100011110011;
      patterns[18336] = 29'b0_100011110100_000_0_100011110100;
      patterns[18337] = 29'b0_100011110100_001_0_110100100011;
      patterns[18338] = 29'b0_100011110100_010_1_000111101000;
      patterns[18339] = 29'b0_100011110100_011_0_001111010001;
      patterns[18340] = 29'b0_100011110100_100_0_010001111010;
      patterns[18341] = 29'b0_100011110100_101_0_001000111101;
      patterns[18342] = 29'b0_100011110100_110_0_100011110100;
      patterns[18343] = 29'b0_100011110100_111_0_100011110100;
      patterns[18344] = 29'b0_100011110101_000_0_100011110101;
      patterns[18345] = 29'b0_100011110101_001_0_110101100011;
      patterns[18346] = 29'b0_100011110101_010_1_000111101010;
      patterns[18347] = 29'b0_100011110101_011_0_001111010101;
      patterns[18348] = 29'b0_100011110101_100_1_010001111010;
      patterns[18349] = 29'b0_100011110101_101_0_101000111101;
      patterns[18350] = 29'b0_100011110101_110_0_100011110101;
      patterns[18351] = 29'b0_100011110101_111_0_100011110101;
      patterns[18352] = 29'b0_100011110110_000_0_100011110110;
      patterns[18353] = 29'b0_100011110110_001_0_110110100011;
      patterns[18354] = 29'b0_100011110110_010_1_000111101100;
      patterns[18355] = 29'b0_100011110110_011_0_001111011001;
      patterns[18356] = 29'b0_100011110110_100_0_010001111011;
      patterns[18357] = 29'b0_100011110110_101_1_001000111101;
      patterns[18358] = 29'b0_100011110110_110_0_100011110110;
      patterns[18359] = 29'b0_100011110110_111_0_100011110110;
      patterns[18360] = 29'b0_100011110111_000_0_100011110111;
      patterns[18361] = 29'b0_100011110111_001_0_110111100011;
      patterns[18362] = 29'b0_100011110111_010_1_000111101110;
      patterns[18363] = 29'b0_100011110111_011_0_001111011101;
      patterns[18364] = 29'b0_100011110111_100_1_010001111011;
      patterns[18365] = 29'b0_100011110111_101_1_101000111101;
      patterns[18366] = 29'b0_100011110111_110_0_100011110111;
      patterns[18367] = 29'b0_100011110111_111_0_100011110111;
      patterns[18368] = 29'b0_100011111000_000_0_100011111000;
      patterns[18369] = 29'b0_100011111000_001_0_111000100011;
      patterns[18370] = 29'b0_100011111000_010_1_000111110000;
      patterns[18371] = 29'b0_100011111000_011_0_001111100001;
      patterns[18372] = 29'b0_100011111000_100_0_010001111100;
      patterns[18373] = 29'b0_100011111000_101_0_001000111110;
      patterns[18374] = 29'b0_100011111000_110_0_100011111000;
      patterns[18375] = 29'b0_100011111000_111_0_100011111000;
      patterns[18376] = 29'b0_100011111001_000_0_100011111001;
      patterns[18377] = 29'b0_100011111001_001_0_111001100011;
      patterns[18378] = 29'b0_100011111001_010_1_000111110010;
      patterns[18379] = 29'b0_100011111001_011_0_001111100101;
      patterns[18380] = 29'b0_100011111001_100_1_010001111100;
      patterns[18381] = 29'b0_100011111001_101_0_101000111110;
      patterns[18382] = 29'b0_100011111001_110_0_100011111001;
      patterns[18383] = 29'b0_100011111001_111_0_100011111001;
      patterns[18384] = 29'b0_100011111010_000_0_100011111010;
      patterns[18385] = 29'b0_100011111010_001_0_111010100011;
      patterns[18386] = 29'b0_100011111010_010_1_000111110100;
      patterns[18387] = 29'b0_100011111010_011_0_001111101001;
      patterns[18388] = 29'b0_100011111010_100_0_010001111101;
      patterns[18389] = 29'b0_100011111010_101_1_001000111110;
      patterns[18390] = 29'b0_100011111010_110_0_100011111010;
      patterns[18391] = 29'b0_100011111010_111_0_100011111010;
      patterns[18392] = 29'b0_100011111011_000_0_100011111011;
      patterns[18393] = 29'b0_100011111011_001_0_111011100011;
      patterns[18394] = 29'b0_100011111011_010_1_000111110110;
      patterns[18395] = 29'b0_100011111011_011_0_001111101101;
      patterns[18396] = 29'b0_100011111011_100_1_010001111101;
      patterns[18397] = 29'b0_100011111011_101_1_101000111110;
      patterns[18398] = 29'b0_100011111011_110_0_100011111011;
      patterns[18399] = 29'b0_100011111011_111_0_100011111011;
      patterns[18400] = 29'b0_100011111100_000_0_100011111100;
      patterns[18401] = 29'b0_100011111100_001_0_111100100011;
      patterns[18402] = 29'b0_100011111100_010_1_000111111000;
      patterns[18403] = 29'b0_100011111100_011_0_001111110001;
      patterns[18404] = 29'b0_100011111100_100_0_010001111110;
      patterns[18405] = 29'b0_100011111100_101_0_001000111111;
      patterns[18406] = 29'b0_100011111100_110_0_100011111100;
      patterns[18407] = 29'b0_100011111100_111_0_100011111100;
      patterns[18408] = 29'b0_100011111101_000_0_100011111101;
      patterns[18409] = 29'b0_100011111101_001_0_111101100011;
      patterns[18410] = 29'b0_100011111101_010_1_000111111010;
      patterns[18411] = 29'b0_100011111101_011_0_001111110101;
      patterns[18412] = 29'b0_100011111101_100_1_010001111110;
      patterns[18413] = 29'b0_100011111101_101_0_101000111111;
      patterns[18414] = 29'b0_100011111101_110_0_100011111101;
      patterns[18415] = 29'b0_100011111101_111_0_100011111101;
      patterns[18416] = 29'b0_100011111110_000_0_100011111110;
      patterns[18417] = 29'b0_100011111110_001_0_111110100011;
      patterns[18418] = 29'b0_100011111110_010_1_000111111100;
      patterns[18419] = 29'b0_100011111110_011_0_001111111001;
      patterns[18420] = 29'b0_100011111110_100_0_010001111111;
      patterns[18421] = 29'b0_100011111110_101_1_001000111111;
      patterns[18422] = 29'b0_100011111110_110_0_100011111110;
      patterns[18423] = 29'b0_100011111110_111_0_100011111110;
      patterns[18424] = 29'b0_100011111111_000_0_100011111111;
      patterns[18425] = 29'b0_100011111111_001_0_111111100011;
      patterns[18426] = 29'b0_100011111111_010_1_000111111110;
      patterns[18427] = 29'b0_100011111111_011_0_001111111101;
      patterns[18428] = 29'b0_100011111111_100_1_010001111111;
      patterns[18429] = 29'b0_100011111111_101_1_101000111111;
      patterns[18430] = 29'b0_100011111111_110_0_100011111111;
      patterns[18431] = 29'b0_100011111111_111_0_100011111111;
      patterns[18432] = 29'b0_100100000000_000_0_100100000000;
      patterns[18433] = 29'b0_100100000000_001_0_000000100100;
      patterns[18434] = 29'b0_100100000000_010_1_001000000000;
      patterns[18435] = 29'b0_100100000000_011_0_010000000001;
      patterns[18436] = 29'b0_100100000000_100_0_010010000000;
      patterns[18437] = 29'b0_100100000000_101_0_001001000000;
      patterns[18438] = 29'b0_100100000000_110_0_100100000000;
      patterns[18439] = 29'b0_100100000000_111_0_100100000000;
      patterns[18440] = 29'b0_100100000001_000_0_100100000001;
      patterns[18441] = 29'b0_100100000001_001_0_000001100100;
      patterns[18442] = 29'b0_100100000001_010_1_001000000010;
      patterns[18443] = 29'b0_100100000001_011_0_010000000101;
      patterns[18444] = 29'b0_100100000001_100_1_010010000000;
      patterns[18445] = 29'b0_100100000001_101_0_101001000000;
      patterns[18446] = 29'b0_100100000001_110_0_100100000001;
      patterns[18447] = 29'b0_100100000001_111_0_100100000001;
      patterns[18448] = 29'b0_100100000010_000_0_100100000010;
      patterns[18449] = 29'b0_100100000010_001_0_000010100100;
      patterns[18450] = 29'b0_100100000010_010_1_001000000100;
      patterns[18451] = 29'b0_100100000010_011_0_010000001001;
      patterns[18452] = 29'b0_100100000010_100_0_010010000001;
      patterns[18453] = 29'b0_100100000010_101_1_001001000000;
      patterns[18454] = 29'b0_100100000010_110_0_100100000010;
      patterns[18455] = 29'b0_100100000010_111_0_100100000010;
      patterns[18456] = 29'b0_100100000011_000_0_100100000011;
      patterns[18457] = 29'b0_100100000011_001_0_000011100100;
      patterns[18458] = 29'b0_100100000011_010_1_001000000110;
      patterns[18459] = 29'b0_100100000011_011_0_010000001101;
      patterns[18460] = 29'b0_100100000011_100_1_010010000001;
      patterns[18461] = 29'b0_100100000011_101_1_101001000000;
      patterns[18462] = 29'b0_100100000011_110_0_100100000011;
      patterns[18463] = 29'b0_100100000011_111_0_100100000011;
      patterns[18464] = 29'b0_100100000100_000_0_100100000100;
      patterns[18465] = 29'b0_100100000100_001_0_000100100100;
      patterns[18466] = 29'b0_100100000100_010_1_001000001000;
      patterns[18467] = 29'b0_100100000100_011_0_010000010001;
      patterns[18468] = 29'b0_100100000100_100_0_010010000010;
      patterns[18469] = 29'b0_100100000100_101_0_001001000001;
      patterns[18470] = 29'b0_100100000100_110_0_100100000100;
      patterns[18471] = 29'b0_100100000100_111_0_100100000100;
      patterns[18472] = 29'b0_100100000101_000_0_100100000101;
      patterns[18473] = 29'b0_100100000101_001_0_000101100100;
      patterns[18474] = 29'b0_100100000101_010_1_001000001010;
      patterns[18475] = 29'b0_100100000101_011_0_010000010101;
      patterns[18476] = 29'b0_100100000101_100_1_010010000010;
      patterns[18477] = 29'b0_100100000101_101_0_101001000001;
      patterns[18478] = 29'b0_100100000101_110_0_100100000101;
      patterns[18479] = 29'b0_100100000101_111_0_100100000101;
      patterns[18480] = 29'b0_100100000110_000_0_100100000110;
      patterns[18481] = 29'b0_100100000110_001_0_000110100100;
      patterns[18482] = 29'b0_100100000110_010_1_001000001100;
      patterns[18483] = 29'b0_100100000110_011_0_010000011001;
      patterns[18484] = 29'b0_100100000110_100_0_010010000011;
      patterns[18485] = 29'b0_100100000110_101_1_001001000001;
      patterns[18486] = 29'b0_100100000110_110_0_100100000110;
      patterns[18487] = 29'b0_100100000110_111_0_100100000110;
      patterns[18488] = 29'b0_100100000111_000_0_100100000111;
      patterns[18489] = 29'b0_100100000111_001_0_000111100100;
      patterns[18490] = 29'b0_100100000111_010_1_001000001110;
      patterns[18491] = 29'b0_100100000111_011_0_010000011101;
      patterns[18492] = 29'b0_100100000111_100_1_010010000011;
      patterns[18493] = 29'b0_100100000111_101_1_101001000001;
      patterns[18494] = 29'b0_100100000111_110_0_100100000111;
      patterns[18495] = 29'b0_100100000111_111_0_100100000111;
      patterns[18496] = 29'b0_100100001000_000_0_100100001000;
      patterns[18497] = 29'b0_100100001000_001_0_001000100100;
      patterns[18498] = 29'b0_100100001000_010_1_001000010000;
      patterns[18499] = 29'b0_100100001000_011_0_010000100001;
      patterns[18500] = 29'b0_100100001000_100_0_010010000100;
      patterns[18501] = 29'b0_100100001000_101_0_001001000010;
      patterns[18502] = 29'b0_100100001000_110_0_100100001000;
      patterns[18503] = 29'b0_100100001000_111_0_100100001000;
      patterns[18504] = 29'b0_100100001001_000_0_100100001001;
      patterns[18505] = 29'b0_100100001001_001_0_001001100100;
      patterns[18506] = 29'b0_100100001001_010_1_001000010010;
      patterns[18507] = 29'b0_100100001001_011_0_010000100101;
      patterns[18508] = 29'b0_100100001001_100_1_010010000100;
      patterns[18509] = 29'b0_100100001001_101_0_101001000010;
      patterns[18510] = 29'b0_100100001001_110_0_100100001001;
      patterns[18511] = 29'b0_100100001001_111_0_100100001001;
      patterns[18512] = 29'b0_100100001010_000_0_100100001010;
      patterns[18513] = 29'b0_100100001010_001_0_001010100100;
      patterns[18514] = 29'b0_100100001010_010_1_001000010100;
      patterns[18515] = 29'b0_100100001010_011_0_010000101001;
      patterns[18516] = 29'b0_100100001010_100_0_010010000101;
      patterns[18517] = 29'b0_100100001010_101_1_001001000010;
      patterns[18518] = 29'b0_100100001010_110_0_100100001010;
      patterns[18519] = 29'b0_100100001010_111_0_100100001010;
      patterns[18520] = 29'b0_100100001011_000_0_100100001011;
      patterns[18521] = 29'b0_100100001011_001_0_001011100100;
      patterns[18522] = 29'b0_100100001011_010_1_001000010110;
      patterns[18523] = 29'b0_100100001011_011_0_010000101101;
      patterns[18524] = 29'b0_100100001011_100_1_010010000101;
      patterns[18525] = 29'b0_100100001011_101_1_101001000010;
      patterns[18526] = 29'b0_100100001011_110_0_100100001011;
      patterns[18527] = 29'b0_100100001011_111_0_100100001011;
      patterns[18528] = 29'b0_100100001100_000_0_100100001100;
      patterns[18529] = 29'b0_100100001100_001_0_001100100100;
      patterns[18530] = 29'b0_100100001100_010_1_001000011000;
      patterns[18531] = 29'b0_100100001100_011_0_010000110001;
      patterns[18532] = 29'b0_100100001100_100_0_010010000110;
      patterns[18533] = 29'b0_100100001100_101_0_001001000011;
      patterns[18534] = 29'b0_100100001100_110_0_100100001100;
      patterns[18535] = 29'b0_100100001100_111_0_100100001100;
      patterns[18536] = 29'b0_100100001101_000_0_100100001101;
      patterns[18537] = 29'b0_100100001101_001_0_001101100100;
      patterns[18538] = 29'b0_100100001101_010_1_001000011010;
      patterns[18539] = 29'b0_100100001101_011_0_010000110101;
      patterns[18540] = 29'b0_100100001101_100_1_010010000110;
      patterns[18541] = 29'b0_100100001101_101_0_101001000011;
      patterns[18542] = 29'b0_100100001101_110_0_100100001101;
      patterns[18543] = 29'b0_100100001101_111_0_100100001101;
      patterns[18544] = 29'b0_100100001110_000_0_100100001110;
      patterns[18545] = 29'b0_100100001110_001_0_001110100100;
      patterns[18546] = 29'b0_100100001110_010_1_001000011100;
      patterns[18547] = 29'b0_100100001110_011_0_010000111001;
      patterns[18548] = 29'b0_100100001110_100_0_010010000111;
      patterns[18549] = 29'b0_100100001110_101_1_001001000011;
      patterns[18550] = 29'b0_100100001110_110_0_100100001110;
      patterns[18551] = 29'b0_100100001110_111_0_100100001110;
      patterns[18552] = 29'b0_100100001111_000_0_100100001111;
      patterns[18553] = 29'b0_100100001111_001_0_001111100100;
      patterns[18554] = 29'b0_100100001111_010_1_001000011110;
      patterns[18555] = 29'b0_100100001111_011_0_010000111101;
      patterns[18556] = 29'b0_100100001111_100_1_010010000111;
      patterns[18557] = 29'b0_100100001111_101_1_101001000011;
      patterns[18558] = 29'b0_100100001111_110_0_100100001111;
      patterns[18559] = 29'b0_100100001111_111_0_100100001111;
      patterns[18560] = 29'b0_100100010000_000_0_100100010000;
      patterns[18561] = 29'b0_100100010000_001_0_010000100100;
      patterns[18562] = 29'b0_100100010000_010_1_001000100000;
      patterns[18563] = 29'b0_100100010000_011_0_010001000001;
      patterns[18564] = 29'b0_100100010000_100_0_010010001000;
      patterns[18565] = 29'b0_100100010000_101_0_001001000100;
      patterns[18566] = 29'b0_100100010000_110_0_100100010000;
      patterns[18567] = 29'b0_100100010000_111_0_100100010000;
      patterns[18568] = 29'b0_100100010001_000_0_100100010001;
      patterns[18569] = 29'b0_100100010001_001_0_010001100100;
      patterns[18570] = 29'b0_100100010001_010_1_001000100010;
      patterns[18571] = 29'b0_100100010001_011_0_010001000101;
      patterns[18572] = 29'b0_100100010001_100_1_010010001000;
      patterns[18573] = 29'b0_100100010001_101_0_101001000100;
      patterns[18574] = 29'b0_100100010001_110_0_100100010001;
      patterns[18575] = 29'b0_100100010001_111_0_100100010001;
      patterns[18576] = 29'b0_100100010010_000_0_100100010010;
      patterns[18577] = 29'b0_100100010010_001_0_010010100100;
      patterns[18578] = 29'b0_100100010010_010_1_001000100100;
      patterns[18579] = 29'b0_100100010010_011_0_010001001001;
      patterns[18580] = 29'b0_100100010010_100_0_010010001001;
      patterns[18581] = 29'b0_100100010010_101_1_001001000100;
      patterns[18582] = 29'b0_100100010010_110_0_100100010010;
      patterns[18583] = 29'b0_100100010010_111_0_100100010010;
      patterns[18584] = 29'b0_100100010011_000_0_100100010011;
      patterns[18585] = 29'b0_100100010011_001_0_010011100100;
      patterns[18586] = 29'b0_100100010011_010_1_001000100110;
      patterns[18587] = 29'b0_100100010011_011_0_010001001101;
      patterns[18588] = 29'b0_100100010011_100_1_010010001001;
      patterns[18589] = 29'b0_100100010011_101_1_101001000100;
      patterns[18590] = 29'b0_100100010011_110_0_100100010011;
      patterns[18591] = 29'b0_100100010011_111_0_100100010011;
      patterns[18592] = 29'b0_100100010100_000_0_100100010100;
      patterns[18593] = 29'b0_100100010100_001_0_010100100100;
      patterns[18594] = 29'b0_100100010100_010_1_001000101000;
      patterns[18595] = 29'b0_100100010100_011_0_010001010001;
      patterns[18596] = 29'b0_100100010100_100_0_010010001010;
      patterns[18597] = 29'b0_100100010100_101_0_001001000101;
      patterns[18598] = 29'b0_100100010100_110_0_100100010100;
      patterns[18599] = 29'b0_100100010100_111_0_100100010100;
      patterns[18600] = 29'b0_100100010101_000_0_100100010101;
      patterns[18601] = 29'b0_100100010101_001_0_010101100100;
      patterns[18602] = 29'b0_100100010101_010_1_001000101010;
      patterns[18603] = 29'b0_100100010101_011_0_010001010101;
      patterns[18604] = 29'b0_100100010101_100_1_010010001010;
      patterns[18605] = 29'b0_100100010101_101_0_101001000101;
      patterns[18606] = 29'b0_100100010101_110_0_100100010101;
      patterns[18607] = 29'b0_100100010101_111_0_100100010101;
      patterns[18608] = 29'b0_100100010110_000_0_100100010110;
      patterns[18609] = 29'b0_100100010110_001_0_010110100100;
      patterns[18610] = 29'b0_100100010110_010_1_001000101100;
      patterns[18611] = 29'b0_100100010110_011_0_010001011001;
      patterns[18612] = 29'b0_100100010110_100_0_010010001011;
      patterns[18613] = 29'b0_100100010110_101_1_001001000101;
      patterns[18614] = 29'b0_100100010110_110_0_100100010110;
      patterns[18615] = 29'b0_100100010110_111_0_100100010110;
      patterns[18616] = 29'b0_100100010111_000_0_100100010111;
      patterns[18617] = 29'b0_100100010111_001_0_010111100100;
      patterns[18618] = 29'b0_100100010111_010_1_001000101110;
      patterns[18619] = 29'b0_100100010111_011_0_010001011101;
      patterns[18620] = 29'b0_100100010111_100_1_010010001011;
      patterns[18621] = 29'b0_100100010111_101_1_101001000101;
      patterns[18622] = 29'b0_100100010111_110_0_100100010111;
      patterns[18623] = 29'b0_100100010111_111_0_100100010111;
      patterns[18624] = 29'b0_100100011000_000_0_100100011000;
      patterns[18625] = 29'b0_100100011000_001_0_011000100100;
      patterns[18626] = 29'b0_100100011000_010_1_001000110000;
      patterns[18627] = 29'b0_100100011000_011_0_010001100001;
      patterns[18628] = 29'b0_100100011000_100_0_010010001100;
      patterns[18629] = 29'b0_100100011000_101_0_001001000110;
      patterns[18630] = 29'b0_100100011000_110_0_100100011000;
      patterns[18631] = 29'b0_100100011000_111_0_100100011000;
      patterns[18632] = 29'b0_100100011001_000_0_100100011001;
      patterns[18633] = 29'b0_100100011001_001_0_011001100100;
      patterns[18634] = 29'b0_100100011001_010_1_001000110010;
      patterns[18635] = 29'b0_100100011001_011_0_010001100101;
      patterns[18636] = 29'b0_100100011001_100_1_010010001100;
      patterns[18637] = 29'b0_100100011001_101_0_101001000110;
      patterns[18638] = 29'b0_100100011001_110_0_100100011001;
      patterns[18639] = 29'b0_100100011001_111_0_100100011001;
      patterns[18640] = 29'b0_100100011010_000_0_100100011010;
      patterns[18641] = 29'b0_100100011010_001_0_011010100100;
      patterns[18642] = 29'b0_100100011010_010_1_001000110100;
      patterns[18643] = 29'b0_100100011010_011_0_010001101001;
      patterns[18644] = 29'b0_100100011010_100_0_010010001101;
      patterns[18645] = 29'b0_100100011010_101_1_001001000110;
      patterns[18646] = 29'b0_100100011010_110_0_100100011010;
      patterns[18647] = 29'b0_100100011010_111_0_100100011010;
      patterns[18648] = 29'b0_100100011011_000_0_100100011011;
      patterns[18649] = 29'b0_100100011011_001_0_011011100100;
      patterns[18650] = 29'b0_100100011011_010_1_001000110110;
      patterns[18651] = 29'b0_100100011011_011_0_010001101101;
      patterns[18652] = 29'b0_100100011011_100_1_010010001101;
      patterns[18653] = 29'b0_100100011011_101_1_101001000110;
      patterns[18654] = 29'b0_100100011011_110_0_100100011011;
      patterns[18655] = 29'b0_100100011011_111_0_100100011011;
      patterns[18656] = 29'b0_100100011100_000_0_100100011100;
      patterns[18657] = 29'b0_100100011100_001_0_011100100100;
      patterns[18658] = 29'b0_100100011100_010_1_001000111000;
      patterns[18659] = 29'b0_100100011100_011_0_010001110001;
      patterns[18660] = 29'b0_100100011100_100_0_010010001110;
      patterns[18661] = 29'b0_100100011100_101_0_001001000111;
      patterns[18662] = 29'b0_100100011100_110_0_100100011100;
      patterns[18663] = 29'b0_100100011100_111_0_100100011100;
      patterns[18664] = 29'b0_100100011101_000_0_100100011101;
      patterns[18665] = 29'b0_100100011101_001_0_011101100100;
      patterns[18666] = 29'b0_100100011101_010_1_001000111010;
      patterns[18667] = 29'b0_100100011101_011_0_010001110101;
      patterns[18668] = 29'b0_100100011101_100_1_010010001110;
      patterns[18669] = 29'b0_100100011101_101_0_101001000111;
      patterns[18670] = 29'b0_100100011101_110_0_100100011101;
      patterns[18671] = 29'b0_100100011101_111_0_100100011101;
      patterns[18672] = 29'b0_100100011110_000_0_100100011110;
      patterns[18673] = 29'b0_100100011110_001_0_011110100100;
      patterns[18674] = 29'b0_100100011110_010_1_001000111100;
      patterns[18675] = 29'b0_100100011110_011_0_010001111001;
      patterns[18676] = 29'b0_100100011110_100_0_010010001111;
      patterns[18677] = 29'b0_100100011110_101_1_001001000111;
      patterns[18678] = 29'b0_100100011110_110_0_100100011110;
      patterns[18679] = 29'b0_100100011110_111_0_100100011110;
      patterns[18680] = 29'b0_100100011111_000_0_100100011111;
      patterns[18681] = 29'b0_100100011111_001_0_011111100100;
      patterns[18682] = 29'b0_100100011111_010_1_001000111110;
      patterns[18683] = 29'b0_100100011111_011_0_010001111101;
      patterns[18684] = 29'b0_100100011111_100_1_010010001111;
      patterns[18685] = 29'b0_100100011111_101_1_101001000111;
      patterns[18686] = 29'b0_100100011111_110_0_100100011111;
      patterns[18687] = 29'b0_100100011111_111_0_100100011111;
      patterns[18688] = 29'b0_100100100000_000_0_100100100000;
      patterns[18689] = 29'b0_100100100000_001_0_100000100100;
      patterns[18690] = 29'b0_100100100000_010_1_001001000000;
      patterns[18691] = 29'b0_100100100000_011_0_010010000001;
      patterns[18692] = 29'b0_100100100000_100_0_010010010000;
      patterns[18693] = 29'b0_100100100000_101_0_001001001000;
      patterns[18694] = 29'b0_100100100000_110_0_100100100000;
      patterns[18695] = 29'b0_100100100000_111_0_100100100000;
      patterns[18696] = 29'b0_100100100001_000_0_100100100001;
      patterns[18697] = 29'b0_100100100001_001_0_100001100100;
      patterns[18698] = 29'b0_100100100001_010_1_001001000010;
      patterns[18699] = 29'b0_100100100001_011_0_010010000101;
      patterns[18700] = 29'b0_100100100001_100_1_010010010000;
      patterns[18701] = 29'b0_100100100001_101_0_101001001000;
      patterns[18702] = 29'b0_100100100001_110_0_100100100001;
      patterns[18703] = 29'b0_100100100001_111_0_100100100001;
      patterns[18704] = 29'b0_100100100010_000_0_100100100010;
      patterns[18705] = 29'b0_100100100010_001_0_100010100100;
      patterns[18706] = 29'b0_100100100010_010_1_001001000100;
      patterns[18707] = 29'b0_100100100010_011_0_010010001001;
      patterns[18708] = 29'b0_100100100010_100_0_010010010001;
      patterns[18709] = 29'b0_100100100010_101_1_001001001000;
      patterns[18710] = 29'b0_100100100010_110_0_100100100010;
      patterns[18711] = 29'b0_100100100010_111_0_100100100010;
      patterns[18712] = 29'b0_100100100011_000_0_100100100011;
      patterns[18713] = 29'b0_100100100011_001_0_100011100100;
      patterns[18714] = 29'b0_100100100011_010_1_001001000110;
      patterns[18715] = 29'b0_100100100011_011_0_010010001101;
      patterns[18716] = 29'b0_100100100011_100_1_010010010001;
      patterns[18717] = 29'b0_100100100011_101_1_101001001000;
      patterns[18718] = 29'b0_100100100011_110_0_100100100011;
      patterns[18719] = 29'b0_100100100011_111_0_100100100011;
      patterns[18720] = 29'b0_100100100100_000_0_100100100100;
      patterns[18721] = 29'b0_100100100100_001_0_100100100100;
      patterns[18722] = 29'b0_100100100100_010_1_001001001000;
      patterns[18723] = 29'b0_100100100100_011_0_010010010001;
      patterns[18724] = 29'b0_100100100100_100_0_010010010010;
      patterns[18725] = 29'b0_100100100100_101_0_001001001001;
      patterns[18726] = 29'b0_100100100100_110_0_100100100100;
      patterns[18727] = 29'b0_100100100100_111_0_100100100100;
      patterns[18728] = 29'b0_100100100101_000_0_100100100101;
      patterns[18729] = 29'b0_100100100101_001_0_100101100100;
      patterns[18730] = 29'b0_100100100101_010_1_001001001010;
      patterns[18731] = 29'b0_100100100101_011_0_010010010101;
      patterns[18732] = 29'b0_100100100101_100_1_010010010010;
      patterns[18733] = 29'b0_100100100101_101_0_101001001001;
      patterns[18734] = 29'b0_100100100101_110_0_100100100101;
      patterns[18735] = 29'b0_100100100101_111_0_100100100101;
      patterns[18736] = 29'b0_100100100110_000_0_100100100110;
      patterns[18737] = 29'b0_100100100110_001_0_100110100100;
      patterns[18738] = 29'b0_100100100110_010_1_001001001100;
      patterns[18739] = 29'b0_100100100110_011_0_010010011001;
      patterns[18740] = 29'b0_100100100110_100_0_010010010011;
      patterns[18741] = 29'b0_100100100110_101_1_001001001001;
      patterns[18742] = 29'b0_100100100110_110_0_100100100110;
      patterns[18743] = 29'b0_100100100110_111_0_100100100110;
      patterns[18744] = 29'b0_100100100111_000_0_100100100111;
      patterns[18745] = 29'b0_100100100111_001_0_100111100100;
      patterns[18746] = 29'b0_100100100111_010_1_001001001110;
      patterns[18747] = 29'b0_100100100111_011_0_010010011101;
      patterns[18748] = 29'b0_100100100111_100_1_010010010011;
      patterns[18749] = 29'b0_100100100111_101_1_101001001001;
      patterns[18750] = 29'b0_100100100111_110_0_100100100111;
      patterns[18751] = 29'b0_100100100111_111_0_100100100111;
      patterns[18752] = 29'b0_100100101000_000_0_100100101000;
      patterns[18753] = 29'b0_100100101000_001_0_101000100100;
      patterns[18754] = 29'b0_100100101000_010_1_001001010000;
      patterns[18755] = 29'b0_100100101000_011_0_010010100001;
      patterns[18756] = 29'b0_100100101000_100_0_010010010100;
      patterns[18757] = 29'b0_100100101000_101_0_001001001010;
      patterns[18758] = 29'b0_100100101000_110_0_100100101000;
      patterns[18759] = 29'b0_100100101000_111_0_100100101000;
      patterns[18760] = 29'b0_100100101001_000_0_100100101001;
      patterns[18761] = 29'b0_100100101001_001_0_101001100100;
      patterns[18762] = 29'b0_100100101001_010_1_001001010010;
      patterns[18763] = 29'b0_100100101001_011_0_010010100101;
      patterns[18764] = 29'b0_100100101001_100_1_010010010100;
      patterns[18765] = 29'b0_100100101001_101_0_101001001010;
      patterns[18766] = 29'b0_100100101001_110_0_100100101001;
      patterns[18767] = 29'b0_100100101001_111_0_100100101001;
      patterns[18768] = 29'b0_100100101010_000_0_100100101010;
      patterns[18769] = 29'b0_100100101010_001_0_101010100100;
      patterns[18770] = 29'b0_100100101010_010_1_001001010100;
      patterns[18771] = 29'b0_100100101010_011_0_010010101001;
      patterns[18772] = 29'b0_100100101010_100_0_010010010101;
      patterns[18773] = 29'b0_100100101010_101_1_001001001010;
      patterns[18774] = 29'b0_100100101010_110_0_100100101010;
      patterns[18775] = 29'b0_100100101010_111_0_100100101010;
      patterns[18776] = 29'b0_100100101011_000_0_100100101011;
      patterns[18777] = 29'b0_100100101011_001_0_101011100100;
      patterns[18778] = 29'b0_100100101011_010_1_001001010110;
      patterns[18779] = 29'b0_100100101011_011_0_010010101101;
      patterns[18780] = 29'b0_100100101011_100_1_010010010101;
      patterns[18781] = 29'b0_100100101011_101_1_101001001010;
      patterns[18782] = 29'b0_100100101011_110_0_100100101011;
      patterns[18783] = 29'b0_100100101011_111_0_100100101011;
      patterns[18784] = 29'b0_100100101100_000_0_100100101100;
      patterns[18785] = 29'b0_100100101100_001_0_101100100100;
      patterns[18786] = 29'b0_100100101100_010_1_001001011000;
      patterns[18787] = 29'b0_100100101100_011_0_010010110001;
      patterns[18788] = 29'b0_100100101100_100_0_010010010110;
      patterns[18789] = 29'b0_100100101100_101_0_001001001011;
      patterns[18790] = 29'b0_100100101100_110_0_100100101100;
      patterns[18791] = 29'b0_100100101100_111_0_100100101100;
      patterns[18792] = 29'b0_100100101101_000_0_100100101101;
      patterns[18793] = 29'b0_100100101101_001_0_101101100100;
      patterns[18794] = 29'b0_100100101101_010_1_001001011010;
      patterns[18795] = 29'b0_100100101101_011_0_010010110101;
      patterns[18796] = 29'b0_100100101101_100_1_010010010110;
      patterns[18797] = 29'b0_100100101101_101_0_101001001011;
      patterns[18798] = 29'b0_100100101101_110_0_100100101101;
      patterns[18799] = 29'b0_100100101101_111_0_100100101101;
      patterns[18800] = 29'b0_100100101110_000_0_100100101110;
      patterns[18801] = 29'b0_100100101110_001_0_101110100100;
      patterns[18802] = 29'b0_100100101110_010_1_001001011100;
      patterns[18803] = 29'b0_100100101110_011_0_010010111001;
      patterns[18804] = 29'b0_100100101110_100_0_010010010111;
      patterns[18805] = 29'b0_100100101110_101_1_001001001011;
      patterns[18806] = 29'b0_100100101110_110_0_100100101110;
      patterns[18807] = 29'b0_100100101110_111_0_100100101110;
      patterns[18808] = 29'b0_100100101111_000_0_100100101111;
      patterns[18809] = 29'b0_100100101111_001_0_101111100100;
      patterns[18810] = 29'b0_100100101111_010_1_001001011110;
      patterns[18811] = 29'b0_100100101111_011_0_010010111101;
      patterns[18812] = 29'b0_100100101111_100_1_010010010111;
      patterns[18813] = 29'b0_100100101111_101_1_101001001011;
      patterns[18814] = 29'b0_100100101111_110_0_100100101111;
      patterns[18815] = 29'b0_100100101111_111_0_100100101111;
      patterns[18816] = 29'b0_100100110000_000_0_100100110000;
      patterns[18817] = 29'b0_100100110000_001_0_110000100100;
      patterns[18818] = 29'b0_100100110000_010_1_001001100000;
      patterns[18819] = 29'b0_100100110000_011_0_010011000001;
      patterns[18820] = 29'b0_100100110000_100_0_010010011000;
      patterns[18821] = 29'b0_100100110000_101_0_001001001100;
      patterns[18822] = 29'b0_100100110000_110_0_100100110000;
      patterns[18823] = 29'b0_100100110000_111_0_100100110000;
      patterns[18824] = 29'b0_100100110001_000_0_100100110001;
      patterns[18825] = 29'b0_100100110001_001_0_110001100100;
      patterns[18826] = 29'b0_100100110001_010_1_001001100010;
      patterns[18827] = 29'b0_100100110001_011_0_010011000101;
      patterns[18828] = 29'b0_100100110001_100_1_010010011000;
      patterns[18829] = 29'b0_100100110001_101_0_101001001100;
      patterns[18830] = 29'b0_100100110001_110_0_100100110001;
      patterns[18831] = 29'b0_100100110001_111_0_100100110001;
      patterns[18832] = 29'b0_100100110010_000_0_100100110010;
      patterns[18833] = 29'b0_100100110010_001_0_110010100100;
      patterns[18834] = 29'b0_100100110010_010_1_001001100100;
      patterns[18835] = 29'b0_100100110010_011_0_010011001001;
      patterns[18836] = 29'b0_100100110010_100_0_010010011001;
      patterns[18837] = 29'b0_100100110010_101_1_001001001100;
      patterns[18838] = 29'b0_100100110010_110_0_100100110010;
      patterns[18839] = 29'b0_100100110010_111_0_100100110010;
      patterns[18840] = 29'b0_100100110011_000_0_100100110011;
      patterns[18841] = 29'b0_100100110011_001_0_110011100100;
      patterns[18842] = 29'b0_100100110011_010_1_001001100110;
      patterns[18843] = 29'b0_100100110011_011_0_010011001101;
      patterns[18844] = 29'b0_100100110011_100_1_010010011001;
      patterns[18845] = 29'b0_100100110011_101_1_101001001100;
      patterns[18846] = 29'b0_100100110011_110_0_100100110011;
      patterns[18847] = 29'b0_100100110011_111_0_100100110011;
      patterns[18848] = 29'b0_100100110100_000_0_100100110100;
      patterns[18849] = 29'b0_100100110100_001_0_110100100100;
      patterns[18850] = 29'b0_100100110100_010_1_001001101000;
      patterns[18851] = 29'b0_100100110100_011_0_010011010001;
      patterns[18852] = 29'b0_100100110100_100_0_010010011010;
      patterns[18853] = 29'b0_100100110100_101_0_001001001101;
      patterns[18854] = 29'b0_100100110100_110_0_100100110100;
      patterns[18855] = 29'b0_100100110100_111_0_100100110100;
      patterns[18856] = 29'b0_100100110101_000_0_100100110101;
      patterns[18857] = 29'b0_100100110101_001_0_110101100100;
      patterns[18858] = 29'b0_100100110101_010_1_001001101010;
      patterns[18859] = 29'b0_100100110101_011_0_010011010101;
      patterns[18860] = 29'b0_100100110101_100_1_010010011010;
      patterns[18861] = 29'b0_100100110101_101_0_101001001101;
      patterns[18862] = 29'b0_100100110101_110_0_100100110101;
      patterns[18863] = 29'b0_100100110101_111_0_100100110101;
      patterns[18864] = 29'b0_100100110110_000_0_100100110110;
      patterns[18865] = 29'b0_100100110110_001_0_110110100100;
      patterns[18866] = 29'b0_100100110110_010_1_001001101100;
      patterns[18867] = 29'b0_100100110110_011_0_010011011001;
      patterns[18868] = 29'b0_100100110110_100_0_010010011011;
      patterns[18869] = 29'b0_100100110110_101_1_001001001101;
      patterns[18870] = 29'b0_100100110110_110_0_100100110110;
      patterns[18871] = 29'b0_100100110110_111_0_100100110110;
      patterns[18872] = 29'b0_100100110111_000_0_100100110111;
      patterns[18873] = 29'b0_100100110111_001_0_110111100100;
      patterns[18874] = 29'b0_100100110111_010_1_001001101110;
      patterns[18875] = 29'b0_100100110111_011_0_010011011101;
      patterns[18876] = 29'b0_100100110111_100_1_010010011011;
      patterns[18877] = 29'b0_100100110111_101_1_101001001101;
      patterns[18878] = 29'b0_100100110111_110_0_100100110111;
      patterns[18879] = 29'b0_100100110111_111_0_100100110111;
      patterns[18880] = 29'b0_100100111000_000_0_100100111000;
      patterns[18881] = 29'b0_100100111000_001_0_111000100100;
      patterns[18882] = 29'b0_100100111000_010_1_001001110000;
      patterns[18883] = 29'b0_100100111000_011_0_010011100001;
      patterns[18884] = 29'b0_100100111000_100_0_010010011100;
      patterns[18885] = 29'b0_100100111000_101_0_001001001110;
      patterns[18886] = 29'b0_100100111000_110_0_100100111000;
      patterns[18887] = 29'b0_100100111000_111_0_100100111000;
      patterns[18888] = 29'b0_100100111001_000_0_100100111001;
      patterns[18889] = 29'b0_100100111001_001_0_111001100100;
      patterns[18890] = 29'b0_100100111001_010_1_001001110010;
      patterns[18891] = 29'b0_100100111001_011_0_010011100101;
      patterns[18892] = 29'b0_100100111001_100_1_010010011100;
      patterns[18893] = 29'b0_100100111001_101_0_101001001110;
      patterns[18894] = 29'b0_100100111001_110_0_100100111001;
      patterns[18895] = 29'b0_100100111001_111_0_100100111001;
      patterns[18896] = 29'b0_100100111010_000_0_100100111010;
      patterns[18897] = 29'b0_100100111010_001_0_111010100100;
      patterns[18898] = 29'b0_100100111010_010_1_001001110100;
      patterns[18899] = 29'b0_100100111010_011_0_010011101001;
      patterns[18900] = 29'b0_100100111010_100_0_010010011101;
      patterns[18901] = 29'b0_100100111010_101_1_001001001110;
      patterns[18902] = 29'b0_100100111010_110_0_100100111010;
      patterns[18903] = 29'b0_100100111010_111_0_100100111010;
      patterns[18904] = 29'b0_100100111011_000_0_100100111011;
      patterns[18905] = 29'b0_100100111011_001_0_111011100100;
      patterns[18906] = 29'b0_100100111011_010_1_001001110110;
      patterns[18907] = 29'b0_100100111011_011_0_010011101101;
      patterns[18908] = 29'b0_100100111011_100_1_010010011101;
      patterns[18909] = 29'b0_100100111011_101_1_101001001110;
      patterns[18910] = 29'b0_100100111011_110_0_100100111011;
      patterns[18911] = 29'b0_100100111011_111_0_100100111011;
      patterns[18912] = 29'b0_100100111100_000_0_100100111100;
      patterns[18913] = 29'b0_100100111100_001_0_111100100100;
      patterns[18914] = 29'b0_100100111100_010_1_001001111000;
      patterns[18915] = 29'b0_100100111100_011_0_010011110001;
      patterns[18916] = 29'b0_100100111100_100_0_010010011110;
      patterns[18917] = 29'b0_100100111100_101_0_001001001111;
      patterns[18918] = 29'b0_100100111100_110_0_100100111100;
      patterns[18919] = 29'b0_100100111100_111_0_100100111100;
      patterns[18920] = 29'b0_100100111101_000_0_100100111101;
      patterns[18921] = 29'b0_100100111101_001_0_111101100100;
      patterns[18922] = 29'b0_100100111101_010_1_001001111010;
      patterns[18923] = 29'b0_100100111101_011_0_010011110101;
      patterns[18924] = 29'b0_100100111101_100_1_010010011110;
      patterns[18925] = 29'b0_100100111101_101_0_101001001111;
      patterns[18926] = 29'b0_100100111101_110_0_100100111101;
      patterns[18927] = 29'b0_100100111101_111_0_100100111101;
      patterns[18928] = 29'b0_100100111110_000_0_100100111110;
      patterns[18929] = 29'b0_100100111110_001_0_111110100100;
      patterns[18930] = 29'b0_100100111110_010_1_001001111100;
      patterns[18931] = 29'b0_100100111110_011_0_010011111001;
      patterns[18932] = 29'b0_100100111110_100_0_010010011111;
      patterns[18933] = 29'b0_100100111110_101_1_001001001111;
      patterns[18934] = 29'b0_100100111110_110_0_100100111110;
      patterns[18935] = 29'b0_100100111110_111_0_100100111110;
      patterns[18936] = 29'b0_100100111111_000_0_100100111111;
      patterns[18937] = 29'b0_100100111111_001_0_111111100100;
      patterns[18938] = 29'b0_100100111111_010_1_001001111110;
      patterns[18939] = 29'b0_100100111111_011_0_010011111101;
      patterns[18940] = 29'b0_100100111111_100_1_010010011111;
      patterns[18941] = 29'b0_100100111111_101_1_101001001111;
      patterns[18942] = 29'b0_100100111111_110_0_100100111111;
      patterns[18943] = 29'b0_100100111111_111_0_100100111111;
      patterns[18944] = 29'b0_100101000000_000_0_100101000000;
      patterns[18945] = 29'b0_100101000000_001_0_000000100101;
      patterns[18946] = 29'b0_100101000000_010_1_001010000000;
      patterns[18947] = 29'b0_100101000000_011_0_010100000001;
      patterns[18948] = 29'b0_100101000000_100_0_010010100000;
      patterns[18949] = 29'b0_100101000000_101_0_001001010000;
      patterns[18950] = 29'b0_100101000000_110_0_100101000000;
      patterns[18951] = 29'b0_100101000000_111_0_100101000000;
      patterns[18952] = 29'b0_100101000001_000_0_100101000001;
      patterns[18953] = 29'b0_100101000001_001_0_000001100101;
      patterns[18954] = 29'b0_100101000001_010_1_001010000010;
      patterns[18955] = 29'b0_100101000001_011_0_010100000101;
      patterns[18956] = 29'b0_100101000001_100_1_010010100000;
      patterns[18957] = 29'b0_100101000001_101_0_101001010000;
      patterns[18958] = 29'b0_100101000001_110_0_100101000001;
      patterns[18959] = 29'b0_100101000001_111_0_100101000001;
      patterns[18960] = 29'b0_100101000010_000_0_100101000010;
      patterns[18961] = 29'b0_100101000010_001_0_000010100101;
      patterns[18962] = 29'b0_100101000010_010_1_001010000100;
      patterns[18963] = 29'b0_100101000010_011_0_010100001001;
      patterns[18964] = 29'b0_100101000010_100_0_010010100001;
      patterns[18965] = 29'b0_100101000010_101_1_001001010000;
      patterns[18966] = 29'b0_100101000010_110_0_100101000010;
      patterns[18967] = 29'b0_100101000010_111_0_100101000010;
      patterns[18968] = 29'b0_100101000011_000_0_100101000011;
      patterns[18969] = 29'b0_100101000011_001_0_000011100101;
      patterns[18970] = 29'b0_100101000011_010_1_001010000110;
      patterns[18971] = 29'b0_100101000011_011_0_010100001101;
      patterns[18972] = 29'b0_100101000011_100_1_010010100001;
      patterns[18973] = 29'b0_100101000011_101_1_101001010000;
      patterns[18974] = 29'b0_100101000011_110_0_100101000011;
      patterns[18975] = 29'b0_100101000011_111_0_100101000011;
      patterns[18976] = 29'b0_100101000100_000_0_100101000100;
      patterns[18977] = 29'b0_100101000100_001_0_000100100101;
      patterns[18978] = 29'b0_100101000100_010_1_001010001000;
      patterns[18979] = 29'b0_100101000100_011_0_010100010001;
      patterns[18980] = 29'b0_100101000100_100_0_010010100010;
      patterns[18981] = 29'b0_100101000100_101_0_001001010001;
      patterns[18982] = 29'b0_100101000100_110_0_100101000100;
      patterns[18983] = 29'b0_100101000100_111_0_100101000100;
      patterns[18984] = 29'b0_100101000101_000_0_100101000101;
      patterns[18985] = 29'b0_100101000101_001_0_000101100101;
      patterns[18986] = 29'b0_100101000101_010_1_001010001010;
      patterns[18987] = 29'b0_100101000101_011_0_010100010101;
      patterns[18988] = 29'b0_100101000101_100_1_010010100010;
      patterns[18989] = 29'b0_100101000101_101_0_101001010001;
      patterns[18990] = 29'b0_100101000101_110_0_100101000101;
      patterns[18991] = 29'b0_100101000101_111_0_100101000101;
      patterns[18992] = 29'b0_100101000110_000_0_100101000110;
      patterns[18993] = 29'b0_100101000110_001_0_000110100101;
      patterns[18994] = 29'b0_100101000110_010_1_001010001100;
      patterns[18995] = 29'b0_100101000110_011_0_010100011001;
      patterns[18996] = 29'b0_100101000110_100_0_010010100011;
      patterns[18997] = 29'b0_100101000110_101_1_001001010001;
      patterns[18998] = 29'b0_100101000110_110_0_100101000110;
      patterns[18999] = 29'b0_100101000110_111_0_100101000110;
      patterns[19000] = 29'b0_100101000111_000_0_100101000111;
      patterns[19001] = 29'b0_100101000111_001_0_000111100101;
      patterns[19002] = 29'b0_100101000111_010_1_001010001110;
      patterns[19003] = 29'b0_100101000111_011_0_010100011101;
      patterns[19004] = 29'b0_100101000111_100_1_010010100011;
      patterns[19005] = 29'b0_100101000111_101_1_101001010001;
      patterns[19006] = 29'b0_100101000111_110_0_100101000111;
      patterns[19007] = 29'b0_100101000111_111_0_100101000111;
      patterns[19008] = 29'b0_100101001000_000_0_100101001000;
      patterns[19009] = 29'b0_100101001000_001_0_001000100101;
      patterns[19010] = 29'b0_100101001000_010_1_001010010000;
      patterns[19011] = 29'b0_100101001000_011_0_010100100001;
      patterns[19012] = 29'b0_100101001000_100_0_010010100100;
      patterns[19013] = 29'b0_100101001000_101_0_001001010010;
      patterns[19014] = 29'b0_100101001000_110_0_100101001000;
      patterns[19015] = 29'b0_100101001000_111_0_100101001000;
      patterns[19016] = 29'b0_100101001001_000_0_100101001001;
      patterns[19017] = 29'b0_100101001001_001_0_001001100101;
      patterns[19018] = 29'b0_100101001001_010_1_001010010010;
      patterns[19019] = 29'b0_100101001001_011_0_010100100101;
      patterns[19020] = 29'b0_100101001001_100_1_010010100100;
      patterns[19021] = 29'b0_100101001001_101_0_101001010010;
      patterns[19022] = 29'b0_100101001001_110_0_100101001001;
      patterns[19023] = 29'b0_100101001001_111_0_100101001001;
      patterns[19024] = 29'b0_100101001010_000_0_100101001010;
      patterns[19025] = 29'b0_100101001010_001_0_001010100101;
      patterns[19026] = 29'b0_100101001010_010_1_001010010100;
      patterns[19027] = 29'b0_100101001010_011_0_010100101001;
      patterns[19028] = 29'b0_100101001010_100_0_010010100101;
      patterns[19029] = 29'b0_100101001010_101_1_001001010010;
      patterns[19030] = 29'b0_100101001010_110_0_100101001010;
      patterns[19031] = 29'b0_100101001010_111_0_100101001010;
      patterns[19032] = 29'b0_100101001011_000_0_100101001011;
      patterns[19033] = 29'b0_100101001011_001_0_001011100101;
      patterns[19034] = 29'b0_100101001011_010_1_001010010110;
      patterns[19035] = 29'b0_100101001011_011_0_010100101101;
      patterns[19036] = 29'b0_100101001011_100_1_010010100101;
      patterns[19037] = 29'b0_100101001011_101_1_101001010010;
      patterns[19038] = 29'b0_100101001011_110_0_100101001011;
      patterns[19039] = 29'b0_100101001011_111_0_100101001011;
      patterns[19040] = 29'b0_100101001100_000_0_100101001100;
      patterns[19041] = 29'b0_100101001100_001_0_001100100101;
      patterns[19042] = 29'b0_100101001100_010_1_001010011000;
      patterns[19043] = 29'b0_100101001100_011_0_010100110001;
      patterns[19044] = 29'b0_100101001100_100_0_010010100110;
      patterns[19045] = 29'b0_100101001100_101_0_001001010011;
      patterns[19046] = 29'b0_100101001100_110_0_100101001100;
      patterns[19047] = 29'b0_100101001100_111_0_100101001100;
      patterns[19048] = 29'b0_100101001101_000_0_100101001101;
      patterns[19049] = 29'b0_100101001101_001_0_001101100101;
      patterns[19050] = 29'b0_100101001101_010_1_001010011010;
      patterns[19051] = 29'b0_100101001101_011_0_010100110101;
      patterns[19052] = 29'b0_100101001101_100_1_010010100110;
      patterns[19053] = 29'b0_100101001101_101_0_101001010011;
      patterns[19054] = 29'b0_100101001101_110_0_100101001101;
      patterns[19055] = 29'b0_100101001101_111_0_100101001101;
      patterns[19056] = 29'b0_100101001110_000_0_100101001110;
      patterns[19057] = 29'b0_100101001110_001_0_001110100101;
      patterns[19058] = 29'b0_100101001110_010_1_001010011100;
      patterns[19059] = 29'b0_100101001110_011_0_010100111001;
      patterns[19060] = 29'b0_100101001110_100_0_010010100111;
      patterns[19061] = 29'b0_100101001110_101_1_001001010011;
      patterns[19062] = 29'b0_100101001110_110_0_100101001110;
      patterns[19063] = 29'b0_100101001110_111_0_100101001110;
      patterns[19064] = 29'b0_100101001111_000_0_100101001111;
      patterns[19065] = 29'b0_100101001111_001_0_001111100101;
      patterns[19066] = 29'b0_100101001111_010_1_001010011110;
      patterns[19067] = 29'b0_100101001111_011_0_010100111101;
      patterns[19068] = 29'b0_100101001111_100_1_010010100111;
      patterns[19069] = 29'b0_100101001111_101_1_101001010011;
      patterns[19070] = 29'b0_100101001111_110_0_100101001111;
      patterns[19071] = 29'b0_100101001111_111_0_100101001111;
      patterns[19072] = 29'b0_100101010000_000_0_100101010000;
      patterns[19073] = 29'b0_100101010000_001_0_010000100101;
      patterns[19074] = 29'b0_100101010000_010_1_001010100000;
      patterns[19075] = 29'b0_100101010000_011_0_010101000001;
      patterns[19076] = 29'b0_100101010000_100_0_010010101000;
      patterns[19077] = 29'b0_100101010000_101_0_001001010100;
      patterns[19078] = 29'b0_100101010000_110_0_100101010000;
      patterns[19079] = 29'b0_100101010000_111_0_100101010000;
      patterns[19080] = 29'b0_100101010001_000_0_100101010001;
      patterns[19081] = 29'b0_100101010001_001_0_010001100101;
      patterns[19082] = 29'b0_100101010001_010_1_001010100010;
      patterns[19083] = 29'b0_100101010001_011_0_010101000101;
      patterns[19084] = 29'b0_100101010001_100_1_010010101000;
      patterns[19085] = 29'b0_100101010001_101_0_101001010100;
      patterns[19086] = 29'b0_100101010001_110_0_100101010001;
      patterns[19087] = 29'b0_100101010001_111_0_100101010001;
      patterns[19088] = 29'b0_100101010010_000_0_100101010010;
      patterns[19089] = 29'b0_100101010010_001_0_010010100101;
      patterns[19090] = 29'b0_100101010010_010_1_001010100100;
      patterns[19091] = 29'b0_100101010010_011_0_010101001001;
      patterns[19092] = 29'b0_100101010010_100_0_010010101001;
      patterns[19093] = 29'b0_100101010010_101_1_001001010100;
      patterns[19094] = 29'b0_100101010010_110_0_100101010010;
      patterns[19095] = 29'b0_100101010010_111_0_100101010010;
      patterns[19096] = 29'b0_100101010011_000_0_100101010011;
      patterns[19097] = 29'b0_100101010011_001_0_010011100101;
      patterns[19098] = 29'b0_100101010011_010_1_001010100110;
      patterns[19099] = 29'b0_100101010011_011_0_010101001101;
      patterns[19100] = 29'b0_100101010011_100_1_010010101001;
      patterns[19101] = 29'b0_100101010011_101_1_101001010100;
      patterns[19102] = 29'b0_100101010011_110_0_100101010011;
      patterns[19103] = 29'b0_100101010011_111_0_100101010011;
      patterns[19104] = 29'b0_100101010100_000_0_100101010100;
      patterns[19105] = 29'b0_100101010100_001_0_010100100101;
      patterns[19106] = 29'b0_100101010100_010_1_001010101000;
      patterns[19107] = 29'b0_100101010100_011_0_010101010001;
      patterns[19108] = 29'b0_100101010100_100_0_010010101010;
      patterns[19109] = 29'b0_100101010100_101_0_001001010101;
      patterns[19110] = 29'b0_100101010100_110_0_100101010100;
      patterns[19111] = 29'b0_100101010100_111_0_100101010100;
      patterns[19112] = 29'b0_100101010101_000_0_100101010101;
      patterns[19113] = 29'b0_100101010101_001_0_010101100101;
      patterns[19114] = 29'b0_100101010101_010_1_001010101010;
      patterns[19115] = 29'b0_100101010101_011_0_010101010101;
      patterns[19116] = 29'b0_100101010101_100_1_010010101010;
      patterns[19117] = 29'b0_100101010101_101_0_101001010101;
      patterns[19118] = 29'b0_100101010101_110_0_100101010101;
      patterns[19119] = 29'b0_100101010101_111_0_100101010101;
      patterns[19120] = 29'b0_100101010110_000_0_100101010110;
      patterns[19121] = 29'b0_100101010110_001_0_010110100101;
      patterns[19122] = 29'b0_100101010110_010_1_001010101100;
      patterns[19123] = 29'b0_100101010110_011_0_010101011001;
      patterns[19124] = 29'b0_100101010110_100_0_010010101011;
      patterns[19125] = 29'b0_100101010110_101_1_001001010101;
      patterns[19126] = 29'b0_100101010110_110_0_100101010110;
      patterns[19127] = 29'b0_100101010110_111_0_100101010110;
      patterns[19128] = 29'b0_100101010111_000_0_100101010111;
      patterns[19129] = 29'b0_100101010111_001_0_010111100101;
      patterns[19130] = 29'b0_100101010111_010_1_001010101110;
      patterns[19131] = 29'b0_100101010111_011_0_010101011101;
      patterns[19132] = 29'b0_100101010111_100_1_010010101011;
      patterns[19133] = 29'b0_100101010111_101_1_101001010101;
      patterns[19134] = 29'b0_100101010111_110_0_100101010111;
      patterns[19135] = 29'b0_100101010111_111_0_100101010111;
      patterns[19136] = 29'b0_100101011000_000_0_100101011000;
      patterns[19137] = 29'b0_100101011000_001_0_011000100101;
      patterns[19138] = 29'b0_100101011000_010_1_001010110000;
      patterns[19139] = 29'b0_100101011000_011_0_010101100001;
      patterns[19140] = 29'b0_100101011000_100_0_010010101100;
      patterns[19141] = 29'b0_100101011000_101_0_001001010110;
      patterns[19142] = 29'b0_100101011000_110_0_100101011000;
      patterns[19143] = 29'b0_100101011000_111_0_100101011000;
      patterns[19144] = 29'b0_100101011001_000_0_100101011001;
      patterns[19145] = 29'b0_100101011001_001_0_011001100101;
      patterns[19146] = 29'b0_100101011001_010_1_001010110010;
      patterns[19147] = 29'b0_100101011001_011_0_010101100101;
      patterns[19148] = 29'b0_100101011001_100_1_010010101100;
      patterns[19149] = 29'b0_100101011001_101_0_101001010110;
      patterns[19150] = 29'b0_100101011001_110_0_100101011001;
      patterns[19151] = 29'b0_100101011001_111_0_100101011001;
      patterns[19152] = 29'b0_100101011010_000_0_100101011010;
      patterns[19153] = 29'b0_100101011010_001_0_011010100101;
      patterns[19154] = 29'b0_100101011010_010_1_001010110100;
      patterns[19155] = 29'b0_100101011010_011_0_010101101001;
      patterns[19156] = 29'b0_100101011010_100_0_010010101101;
      patterns[19157] = 29'b0_100101011010_101_1_001001010110;
      patterns[19158] = 29'b0_100101011010_110_0_100101011010;
      patterns[19159] = 29'b0_100101011010_111_0_100101011010;
      patterns[19160] = 29'b0_100101011011_000_0_100101011011;
      patterns[19161] = 29'b0_100101011011_001_0_011011100101;
      patterns[19162] = 29'b0_100101011011_010_1_001010110110;
      patterns[19163] = 29'b0_100101011011_011_0_010101101101;
      patterns[19164] = 29'b0_100101011011_100_1_010010101101;
      patterns[19165] = 29'b0_100101011011_101_1_101001010110;
      patterns[19166] = 29'b0_100101011011_110_0_100101011011;
      patterns[19167] = 29'b0_100101011011_111_0_100101011011;
      patterns[19168] = 29'b0_100101011100_000_0_100101011100;
      patterns[19169] = 29'b0_100101011100_001_0_011100100101;
      patterns[19170] = 29'b0_100101011100_010_1_001010111000;
      patterns[19171] = 29'b0_100101011100_011_0_010101110001;
      patterns[19172] = 29'b0_100101011100_100_0_010010101110;
      patterns[19173] = 29'b0_100101011100_101_0_001001010111;
      patterns[19174] = 29'b0_100101011100_110_0_100101011100;
      patterns[19175] = 29'b0_100101011100_111_0_100101011100;
      patterns[19176] = 29'b0_100101011101_000_0_100101011101;
      patterns[19177] = 29'b0_100101011101_001_0_011101100101;
      patterns[19178] = 29'b0_100101011101_010_1_001010111010;
      patterns[19179] = 29'b0_100101011101_011_0_010101110101;
      patterns[19180] = 29'b0_100101011101_100_1_010010101110;
      patterns[19181] = 29'b0_100101011101_101_0_101001010111;
      patterns[19182] = 29'b0_100101011101_110_0_100101011101;
      patterns[19183] = 29'b0_100101011101_111_0_100101011101;
      patterns[19184] = 29'b0_100101011110_000_0_100101011110;
      patterns[19185] = 29'b0_100101011110_001_0_011110100101;
      patterns[19186] = 29'b0_100101011110_010_1_001010111100;
      patterns[19187] = 29'b0_100101011110_011_0_010101111001;
      patterns[19188] = 29'b0_100101011110_100_0_010010101111;
      patterns[19189] = 29'b0_100101011110_101_1_001001010111;
      patterns[19190] = 29'b0_100101011110_110_0_100101011110;
      patterns[19191] = 29'b0_100101011110_111_0_100101011110;
      patterns[19192] = 29'b0_100101011111_000_0_100101011111;
      patterns[19193] = 29'b0_100101011111_001_0_011111100101;
      patterns[19194] = 29'b0_100101011111_010_1_001010111110;
      patterns[19195] = 29'b0_100101011111_011_0_010101111101;
      patterns[19196] = 29'b0_100101011111_100_1_010010101111;
      patterns[19197] = 29'b0_100101011111_101_1_101001010111;
      patterns[19198] = 29'b0_100101011111_110_0_100101011111;
      patterns[19199] = 29'b0_100101011111_111_0_100101011111;
      patterns[19200] = 29'b0_100101100000_000_0_100101100000;
      patterns[19201] = 29'b0_100101100000_001_0_100000100101;
      patterns[19202] = 29'b0_100101100000_010_1_001011000000;
      patterns[19203] = 29'b0_100101100000_011_0_010110000001;
      patterns[19204] = 29'b0_100101100000_100_0_010010110000;
      patterns[19205] = 29'b0_100101100000_101_0_001001011000;
      patterns[19206] = 29'b0_100101100000_110_0_100101100000;
      patterns[19207] = 29'b0_100101100000_111_0_100101100000;
      patterns[19208] = 29'b0_100101100001_000_0_100101100001;
      patterns[19209] = 29'b0_100101100001_001_0_100001100101;
      patterns[19210] = 29'b0_100101100001_010_1_001011000010;
      patterns[19211] = 29'b0_100101100001_011_0_010110000101;
      patterns[19212] = 29'b0_100101100001_100_1_010010110000;
      patterns[19213] = 29'b0_100101100001_101_0_101001011000;
      patterns[19214] = 29'b0_100101100001_110_0_100101100001;
      patterns[19215] = 29'b0_100101100001_111_0_100101100001;
      patterns[19216] = 29'b0_100101100010_000_0_100101100010;
      patterns[19217] = 29'b0_100101100010_001_0_100010100101;
      patterns[19218] = 29'b0_100101100010_010_1_001011000100;
      patterns[19219] = 29'b0_100101100010_011_0_010110001001;
      patterns[19220] = 29'b0_100101100010_100_0_010010110001;
      patterns[19221] = 29'b0_100101100010_101_1_001001011000;
      patterns[19222] = 29'b0_100101100010_110_0_100101100010;
      patterns[19223] = 29'b0_100101100010_111_0_100101100010;
      patterns[19224] = 29'b0_100101100011_000_0_100101100011;
      patterns[19225] = 29'b0_100101100011_001_0_100011100101;
      patterns[19226] = 29'b0_100101100011_010_1_001011000110;
      patterns[19227] = 29'b0_100101100011_011_0_010110001101;
      patterns[19228] = 29'b0_100101100011_100_1_010010110001;
      patterns[19229] = 29'b0_100101100011_101_1_101001011000;
      patterns[19230] = 29'b0_100101100011_110_0_100101100011;
      patterns[19231] = 29'b0_100101100011_111_0_100101100011;
      patterns[19232] = 29'b0_100101100100_000_0_100101100100;
      patterns[19233] = 29'b0_100101100100_001_0_100100100101;
      patterns[19234] = 29'b0_100101100100_010_1_001011001000;
      patterns[19235] = 29'b0_100101100100_011_0_010110010001;
      patterns[19236] = 29'b0_100101100100_100_0_010010110010;
      patterns[19237] = 29'b0_100101100100_101_0_001001011001;
      patterns[19238] = 29'b0_100101100100_110_0_100101100100;
      patterns[19239] = 29'b0_100101100100_111_0_100101100100;
      patterns[19240] = 29'b0_100101100101_000_0_100101100101;
      patterns[19241] = 29'b0_100101100101_001_0_100101100101;
      patterns[19242] = 29'b0_100101100101_010_1_001011001010;
      patterns[19243] = 29'b0_100101100101_011_0_010110010101;
      patterns[19244] = 29'b0_100101100101_100_1_010010110010;
      patterns[19245] = 29'b0_100101100101_101_0_101001011001;
      patterns[19246] = 29'b0_100101100101_110_0_100101100101;
      patterns[19247] = 29'b0_100101100101_111_0_100101100101;
      patterns[19248] = 29'b0_100101100110_000_0_100101100110;
      patterns[19249] = 29'b0_100101100110_001_0_100110100101;
      patterns[19250] = 29'b0_100101100110_010_1_001011001100;
      patterns[19251] = 29'b0_100101100110_011_0_010110011001;
      patterns[19252] = 29'b0_100101100110_100_0_010010110011;
      patterns[19253] = 29'b0_100101100110_101_1_001001011001;
      patterns[19254] = 29'b0_100101100110_110_0_100101100110;
      patterns[19255] = 29'b0_100101100110_111_0_100101100110;
      patterns[19256] = 29'b0_100101100111_000_0_100101100111;
      patterns[19257] = 29'b0_100101100111_001_0_100111100101;
      patterns[19258] = 29'b0_100101100111_010_1_001011001110;
      patterns[19259] = 29'b0_100101100111_011_0_010110011101;
      patterns[19260] = 29'b0_100101100111_100_1_010010110011;
      patterns[19261] = 29'b0_100101100111_101_1_101001011001;
      patterns[19262] = 29'b0_100101100111_110_0_100101100111;
      patterns[19263] = 29'b0_100101100111_111_0_100101100111;
      patterns[19264] = 29'b0_100101101000_000_0_100101101000;
      patterns[19265] = 29'b0_100101101000_001_0_101000100101;
      patterns[19266] = 29'b0_100101101000_010_1_001011010000;
      patterns[19267] = 29'b0_100101101000_011_0_010110100001;
      patterns[19268] = 29'b0_100101101000_100_0_010010110100;
      patterns[19269] = 29'b0_100101101000_101_0_001001011010;
      patterns[19270] = 29'b0_100101101000_110_0_100101101000;
      patterns[19271] = 29'b0_100101101000_111_0_100101101000;
      patterns[19272] = 29'b0_100101101001_000_0_100101101001;
      patterns[19273] = 29'b0_100101101001_001_0_101001100101;
      patterns[19274] = 29'b0_100101101001_010_1_001011010010;
      patterns[19275] = 29'b0_100101101001_011_0_010110100101;
      patterns[19276] = 29'b0_100101101001_100_1_010010110100;
      patterns[19277] = 29'b0_100101101001_101_0_101001011010;
      patterns[19278] = 29'b0_100101101001_110_0_100101101001;
      patterns[19279] = 29'b0_100101101001_111_0_100101101001;
      patterns[19280] = 29'b0_100101101010_000_0_100101101010;
      patterns[19281] = 29'b0_100101101010_001_0_101010100101;
      patterns[19282] = 29'b0_100101101010_010_1_001011010100;
      patterns[19283] = 29'b0_100101101010_011_0_010110101001;
      patterns[19284] = 29'b0_100101101010_100_0_010010110101;
      patterns[19285] = 29'b0_100101101010_101_1_001001011010;
      patterns[19286] = 29'b0_100101101010_110_0_100101101010;
      patterns[19287] = 29'b0_100101101010_111_0_100101101010;
      patterns[19288] = 29'b0_100101101011_000_0_100101101011;
      patterns[19289] = 29'b0_100101101011_001_0_101011100101;
      patterns[19290] = 29'b0_100101101011_010_1_001011010110;
      patterns[19291] = 29'b0_100101101011_011_0_010110101101;
      patterns[19292] = 29'b0_100101101011_100_1_010010110101;
      patterns[19293] = 29'b0_100101101011_101_1_101001011010;
      patterns[19294] = 29'b0_100101101011_110_0_100101101011;
      patterns[19295] = 29'b0_100101101011_111_0_100101101011;
      patterns[19296] = 29'b0_100101101100_000_0_100101101100;
      patterns[19297] = 29'b0_100101101100_001_0_101100100101;
      patterns[19298] = 29'b0_100101101100_010_1_001011011000;
      patterns[19299] = 29'b0_100101101100_011_0_010110110001;
      patterns[19300] = 29'b0_100101101100_100_0_010010110110;
      patterns[19301] = 29'b0_100101101100_101_0_001001011011;
      patterns[19302] = 29'b0_100101101100_110_0_100101101100;
      patterns[19303] = 29'b0_100101101100_111_0_100101101100;
      patterns[19304] = 29'b0_100101101101_000_0_100101101101;
      patterns[19305] = 29'b0_100101101101_001_0_101101100101;
      patterns[19306] = 29'b0_100101101101_010_1_001011011010;
      patterns[19307] = 29'b0_100101101101_011_0_010110110101;
      patterns[19308] = 29'b0_100101101101_100_1_010010110110;
      patterns[19309] = 29'b0_100101101101_101_0_101001011011;
      patterns[19310] = 29'b0_100101101101_110_0_100101101101;
      patterns[19311] = 29'b0_100101101101_111_0_100101101101;
      patterns[19312] = 29'b0_100101101110_000_0_100101101110;
      patterns[19313] = 29'b0_100101101110_001_0_101110100101;
      patterns[19314] = 29'b0_100101101110_010_1_001011011100;
      patterns[19315] = 29'b0_100101101110_011_0_010110111001;
      patterns[19316] = 29'b0_100101101110_100_0_010010110111;
      patterns[19317] = 29'b0_100101101110_101_1_001001011011;
      patterns[19318] = 29'b0_100101101110_110_0_100101101110;
      patterns[19319] = 29'b0_100101101110_111_0_100101101110;
      patterns[19320] = 29'b0_100101101111_000_0_100101101111;
      patterns[19321] = 29'b0_100101101111_001_0_101111100101;
      patterns[19322] = 29'b0_100101101111_010_1_001011011110;
      patterns[19323] = 29'b0_100101101111_011_0_010110111101;
      patterns[19324] = 29'b0_100101101111_100_1_010010110111;
      patterns[19325] = 29'b0_100101101111_101_1_101001011011;
      patterns[19326] = 29'b0_100101101111_110_0_100101101111;
      patterns[19327] = 29'b0_100101101111_111_0_100101101111;
      patterns[19328] = 29'b0_100101110000_000_0_100101110000;
      patterns[19329] = 29'b0_100101110000_001_0_110000100101;
      patterns[19330] = 29'b0_100101110000_010_1_001011100000;
      patterns[19331] = 29'b0_100101110000_011_0_010111000001;
      patterns[19332] = 29'b0_100101110000_100_0_010010111000;
      patterns[19333] = 29'b0_100101110000_101_0_001001011100;
      patterns[19334] = 29'b0_100101110000_110_0_100101110000;
      patterns[19335] = 29'b0_100101110000_111_0_100101110000;
      patterns[19336] = 29'b0_100101110001_000_0_100101110001;
      patterns[19337] = 29'b0_100101110001_001_0_110001100101;
      patterns[19338] = 29'b0_100101110001_010_1_001011100010;
      patterns[19339] = 29'b0_100101110001_011_0_010111000101;
      patterns[19340] = 29'b0_100101110001_100_1_010010111000;
      patterns[19341] = 29'b0_100101110001_101_0_101001011100;
      patterns[19342] = 29'b0_100101110001_110_0_100101110001;
      patterns[19343] = 29'b0_100101110001_111_0_100101110001;
      patterns[19344] = 29'b0_100101110010_000_0_100101110010;
      patterns[19345] = 29'b0_100101110010_001_0_110010100101;
      patterns[19346] = 29'b0_100101110010_010_1_001011100100;
      patterns[19347] = 29'b0_100101110010_011_0_010111001001;
      patterns[19348] = 29'b0_100101110010_100_0_010010111001;
      patterns[19349] = 29'b0_100101110010_101_1_001001011100;
      patterns[19350] = 29'b0_100101110010_110_0_100101110010;
      patterns[19351] = 29'b0_100101110010_111_0_100101110010;
      patterns[19352] = 29'b0_100101110011_000_0_100101110011;
      patterns[19353] = 29'b0_100101110011_001_0_110011100101;
      patterns[19354] = 29'b0_100101110011_010_1_001011100110;
      patterns[19355] = 29'b0_100101110011_011_0_010111001101;
      patterns[19356] = 29'b0_100101110011_100_1_010010111001;
      patterns[19357] = 29'b0_100101110011_101_1_101001011100;
      patterns[19358] = 29'b0_100101110011_110_0_100101110011;
      patterns[19359] = 29'b0_100101110011_111_0_100101110011;
      patterns[19360] = 29'b0_100101110100_000_0_100101110100;
      patterns[19361] = 29'b0_100101110100_001_0_110100100101;
      patterns[19362] = 29'b0_100101110100_010_1_001011101000;
      patterns[19363] = 29'b0_100101110100_011_0_010111010001;
      patterns[19364] = 29'b0_100101110100_100_0_010010111010;
      patterns[19365] = 29'b0_100101110100_101_0_001001011101;
      patterns[19366] = 29'b0_100101110100_110_0_100101110100;
      patterns[19367] = 29'b0_100101110100_111_0_100101110100;
      patterns[19368] = 29'b0_100101110101_000_0_100101110101;
      patterns[19369] = 29'b0_100101110101_001_0_110101100101;
      patterns[19370] = 29'b0_100101110101_010_1_001011101010;
      patterns[19371] = 29'b0_100101110101_011_0_010111010101;
      patterns[19372] = 29'b0_100101110101_100_1_010010111010;
      patterns[19373] = 29'b0_100101110101_101_0_101001011101;
      patterns[19374] = 29'b0_100101110101_110_0_100101110101;
      patterns[19375] = 29'b0_100101110101_111_0_100101110101;
      patterns[19376] = 29'b0_100101110110_000_0_100101110110;
      patterns[19377] = 29'b0_100101110110_001_0_110110100101;
      patterns[19378] = 29'b0_100101110110_010_1_001011101100;
      patterns[19379] = 29'b0_100101110110_011_0_010111011001;
      patterns[19380] = 29'b0_100101110110_100_0_010010111011;
      patterns[19381] = 29'b0_100101110110_101_1_001001011101;
      patterns[19382] = 29'b0_100101110110_110_0_100101110110;
      patterns[19383] = 29'b0_100101110110_111_0_100101110110;
      patterns[19384] = 29'b0_100101110111_000_0_100101110111;
      patterns[19385] = 29'b0_100101110111_001_0_110111100101;
      patterns[19386] = 29'b0_100101110111_010_1_001011101110;
      patterns[19387] = 29'b0_100101110111_011_0_010111011101;
      patterns[19388] = 29'b0_100101110111_100_1_010010111011;
      patterns[19389] = 29'b0_100101110111_101_1_101001011101;
      patterns[19390] = 29'b0_100101110111_110_0_100101110111;
      patterns[19391] = 29'b0_100101110111_111_0_100101110111;
      patterns[19392] = 29'b0_100101111000_000_0_100101111000;
      patterns[19393] = 29'b0_100101111000_001_0_111000100101;
      patterns[19394] = 29'b0_100101111000_010_1_001011110000;
      patterns[19395] = 29'b0_100101111000_011_0_010111100001;
      patterns[19396] = 29'b0_100101111000_100_0_010010111100;
      patterns[19397] = 29'b0_100101111000_101_0_001001011110;
      patterns[19398] = 29'b0_100101111000_110_0_100101111000;
      patterns[19399] = 29'b0_100101111000_111_0_100101111000;
      patterns[19400] = 29'b0_100101111001_000_0_100101111001;
      patterns[19401] = 29'b0_100101111001_001_0_111001100101;
      patterns[19402] = 29'b0_100101111001_010_1_001011110010;
      patterns[19403] = 29'b0_100101111001_011_0_010111100101;
      patterns[19404] = 29'b0_100101111001_100_1_010010111100;
      patterns[19405] = 29'b0_100101111001_101_0_101001011110;
      patterns[19406] = 29'b0_100101111001_110_0_100101111001;
      patterns[19407] = 29'b0_100101111001_111_0_100101111001;
      patterns[19408] = 29'b0_100101111010_000_0_100101111010;
      patterns[19409] = 29'b0_100101111010_001_0_111010100101;
      patterns[19410] = 29'b0_100101111010_010_1_001011110100;
      patterns[19411] = 29'b0_100101111010_011_0_010111101001;
      patterns[19412] = 29'b0_100101111010_100_0_010010111101;
      patterns[19413] = 29'b0_100101111010_101_1_001001011110;
      patterns[19414] = 29'b0_100101111010_110_0_100101111010;
      patterns[19415] = 29'b0_100101111010_111_0_100101111010;
      patterns[19416] = 29'b0_100101111011_000_0_100101111011;
      patterns[19417] = 29'b0_100101111011_001_0_111011100101;
      patterns[19418] = 29'b0_100101111011_010_1_001011110110;
      patterns[19419] = 29'b0_100101111011_011_0_010111101101;
      patterns[19420] = 29'b0_100101111011_100_1_010010111101;
      patterns[19421] = 29'b0_100101111011_101_1_101001011110;
      patterns[19422] = 29'b0_100101111011_110_0_100101111011;
      patterns[19423] = 29'b0_100101111011_111_0_100101111011;
      patterns[19424] = 29'b0_100101111100_000_0_100101111100;
      patterns[19425] = 29'b0_100101111100_001_0_111100100101;
      patterns[19426] = 29'b0_100101111100_010_1_001011111000;
      patterns[19427] = 29'b0_100101111100_011_0_010111110001;
      patterns[19428] = 29'b0_100101111100_100_0_010010111110;
      patterns[19429] = 29'b0_100101111100_101_0_001001011111;
      patterns[19430] = 29'b0_100101111100_110_0_100101111100;
      patterns[19431] = 29'b0_100101111100_111_0_100101111100;
      patterns[19432] = 29'b0_100101111101_000_0_100101111101;
      patterns[19433] = 29'b0_100101111101_001_0_111101100101;
      patterns[19434] = 29'b0_100101111101_010_1_001011111010;
      patterns[19435] = 29'b0_100101111101_011_0_010111110101;
      patterns[19436] = 29'b0_100101111101_100_1_010010111110;
      patterns[19437] = 29'b0_100101111101_101_0_101001011111;
      patterns[19438] = 29'b0_100101111101_110_0_100101111101;
      patterns[19439] = 29'b0_100101111101_111_0_100101111101;
      patterns[19440] = 29'b0_100101111110_000_0_100101111110;
      patterns[19441] = 29'b0_100101111110_001_0_111110100101;
      patterns[19442] = 29'b0_100101111110_010_1_001011111100;
      patterns[19443] = 29'b0_100101111110_011_0_010111111001;
      patterns[19444] = 29'b0_100101111110_100_0_010010111111;
      patterns[19445] = 29'b0_100101111110_101_1_001001011111;
      patterns[19446] = 29'b0_100101111110_110_0_100101111110;
      patterns[19447] = 29'b0_100101111110_111_0_100101111110;
      patterns[19448] = 29'b0_100101111111_000_0_100101111111;
      patterns[19449] = 29'b0_100101111111_001_0_111111100101;
      patterns[19450] = 29'b0_100101111111_010_1_001011111110;
      patterns[19451] = 29'b0_100101111111_011_0_010111111101;
      patterns[19452] = 29'b0_100101111111_100_1_010010111111;
      patterns[19453] = 29'b0_100101111111_101_1_101001011111;
      patterns[19454] = 29'b0_100101111111_110_0_100101111111;
      patterns[19455] = 29'b0_100101111111_111_0_100101111111;
      patterns[19456] = 29'b0_100110000000_000_0_100110000000;
      patterns[19457] = 29'b0_100110000000_001_0_000000100110;
      patterns[19458] = 29'b0_100110000000_010_1_001100000000;
      patterns[19459] = 29'b0_100110000000_011_0_011000000001;
      patterns[19460] = 29'b0_100110000000_100_0_010011000000;
      patterns[19461] = 29'b0_100110000000_101_0_001001100000;
      patterns[19462] = 29'b0_100110000000_110_0_100110000000;
      patterns[19463] = 29'b0_100110000000_111_0_100110000000;
      patterns[19464] = 29'b0_100110000001_000_0_100110000001;
      patterns[19465] = 29'b0_100110000001_001_0_000001100110;
      patterns[19466] = 29'b0_100110000001_010_1_001100000010;
      patterns[19467] = 29'b0_100110000001_011_0_011000000101;
      patterns[19468] = 29'b0_100110000001_100_1_010011000000;
      patterns[19469] = 29'b0_100110000001_101_0_101001100000;
      patterns[19470] = 29'b0_100110000001_110_0_100110000001;
      patterns[19471] = 29'b0_100110000001_111_0_100110000001;
      patterns[19472] = 29'b0_100110000010_000_0_100110000010;
      patterns[19473] = 29'b0_100110000010_001_0_000010100110;
      patterns[19474] = 29'b0_100110000010_010_1_001100000100;
      patterns[19475] = 29'b0_100110000010_011_0_011000001001;
      patterns[19476] = 29'b0_100110000010_100_0_010011000001;
      patterns[19477] = 29'b0_100110000010_101_1_001001100000;
      patterns[19478] = 29'b0_100110000010_110_0_100110000010;
      patterns[19479] = 29'b0_100110000010_111_0_100110000010;
      patterns[19480] = 29'b0_100110000011_000_0_100110000011;
      patterns[19481] = 29'b0_100110000011_001_0_000011100110;
      patterns[19482] = 29'b0_100110000011_010_1_001100000110;
      patterns[19483] = 29'b0_100110000011_011_0_011000001101;
      patterns[19484] = 29'b0_100110000011_100_1_010011000001;
      patterns[19485] = 29'b0_100110000011_101_1_101001100000;
      patterns[19486] = 29'b0_100110000011_110_0_100110000011;
      patterns[19487] = 29'b0_100110000011_111_0_100110000011;
      patterns[19488] = 29'b0_100110000100_000_0_100110000100;
      patterns[19489] = 29'b0_100110000100_001_0_000100100110;
      patterns[19490] = 29'b0_100110000100_010_1_001100001000;
      patterns[19491] = 29'b0_100110000100_011_0_011000010001;
      patterns[19492] = 29'b0_100110000100_100_0_010011000010;
      patterns[19493] = 29'b0_100110000100_101_0_001001100001;
      patterns[19494] = 29'b0_100110000100_110_0_100110000100;
      patterns[19495] = 29'b0_100110000100_111_0_100110000100;
      patterns[19496] = 29'b0_100110000101_000_0_100110000101;
      patterns[19497] = 29'b0_100110000101_001_0_000101100110;
      patterns[19498] = 29'b0_100110000101_010_1_001100001010;
      patterns[19499] = 29'b0_100110000101_011_0_011000010101;
      patterns[19500] = 29'b0_100110000101_100_1_010011000010;
      patterns[19501] = 29'b0_100110000101_101_0_101001100001;
      patterns[19502] = 29'b0_100110000101_110_0_100110000101;
      patterns[19503] = 29'b0_100110000101_111_0_100110000101;
      patterns[19504] = 29'b0_100110000110_000_0_100110000110;
      patterns[19505] = 29'b0_100110000110_001_0_000110100110;
      patterns[19506] = 29'b0_100110000110_010_1_001100001100;
      patterns[19507] = 29'b0_100110000110_011_0_011000011001;
      patterns[19508] = 29'b0_100110000110_100_0_010011000011;
      patterns[19509] = 29'b0_100110000110_101_1_001001100001;
      patterns[19510] = 29'b0_100110000110_110_0_100110000110;
      patterns[19511] = 29'b0_100110000110_111_0_100110000110;
      patterns[19512] = 29'b0_100110000111_000_0_100110000111;
      patterns[19513] = 29'b0_100110000111_001_0_000111100110;
      patterns[19514] = 29'b0_100110000111_010_1_001100001110;
      patterns[19515] = 29'b0_100110000111_011_0_011000011101;
      patterns[19516] = 29'b0_100110000111_100_1_010011000011;
      patterns[19517] = 29'b0_100110000111_101_1_101001100001;
      patterns[19518] = 29'b0_100110000111_110_0_100110000111;
      patterns[19519] = 29'b0_100110000111_111_0_100110000111;
      patterns[19520] = 29'b0_100110001000_000_0_100110001000;
      patterns[19521] = 29'b0_100110001000_001_0_001000100110;
      patterns[19522] = 29'b0_100110001000_010_1_001100010000;
      patterns[19523] = 29'b0_100110001000_011_0_011000100001;
      patterns[19524] = 29'b0_100110001000_100_0_010011000100;
      patterns[19525] = 29'b0_100110001000_101_0_001001100010;
      patterns[19526] = 29'b0_100110001000_110_0_100110001000;
      patterns[19527] = 29'b0_100110001000_111_0_100110001000;
      patterns[19528] = 29'b0_100110001001_000_0_100110001001;
      patterns[19529] = 29'b0_100110001001_001_0_001001100110;
      patterns[19530] = 29'b0_100110001001_010_1_001100010010;
      patterns[19531] = 29'b0_100110001001_011_0_011000100101;
      patterns[19532] = 29'b0_100110001001_100_1_010011000100;
      patterns[19533] = 29'b0_100110001001_101_0_101001100010;
      patterns[19534] = 29'b0_100110001001_110_0_100110001001;
      patterns[19535] = 29'b0_100110001001_111_0_100110001001;
      patterns[19536] = 29'b0_100110001010_000_0_100110001010;
      patterns[19537] = 29'b0_100110001010_001_0_001010100110;
      patterns[19538] = 29'b0_100110001010_010_1_001100010100;
      patterns[19539] = 29'b0_100110001010_011_0_011000101001;
      patterns[19540] = 29'b0_100110001010_100_0_010011000101;
      patterns[19541] = 29'b0_100110001010_101_1_001001100010;
      patterns[19542] = 29'b0_100110001010_110_0_100110001010;
      patterns[19543] = 29'b0_100110001010_111_0_100110001010;
      patterns[19544] = 29'b0_100110001011_000_0_100110001011;
      patterns[19545] = 29'b0_100110001011_001_0_001011100110;
      patterns[19546] = 29'b0_100110001011_010_1_001100010110;
      patterns[19547] = 29'b0_100110001011_011_0_011000101101;
      patterns[19548] = 29'b0_100110001011_100_1_010011000101;
      patterns[19549] = 29'b0_100110001011_101_1_101001100010;
      patterns[19550] = 29'b0_100110001011_110_0_100110001011;
      patterns[19551] = 29'b0_100110001011_111_0_100110001011;
      patterns[19552] = 29'b0_100110001100_000_0_100110001100;
      patterns[19553] = 29'b0_100110001100_001_0_001100100110;
      patterns[19554] = 29'b0_100110001100_010_1_001100011000;
      patterns[19555] = 29'b0_100110001100_011_0_011000110001;
      patterns[19556] = 29'b0_100110001100_100_0_010011000110;
      patterns[19557] = 29'b0_100110001100_101_0_001001100011;
      patterns[19558] = 29'b0_100110001100_110_0_100110001100;
      patterns[19559] = 29'b0_100110001100_111_0_100110001100;
      patterns[19560] = 29'b0_100110001101_000_0_100110001101;
      patterns[19561] = 29'b0_100110001101_001_0_001101100110;
      patterns[19562] = 29'b0_100110001101_010_1_001100011010;
      patterns[19563] = 29'b0_100110001101_011_0_011000110101;
      patterns[19564] = 29'b0_100110001101_100_1_010011000110;
      patterns[19565] = 29'b0_100110001101_101_0_101001100011;
      patterns[19566] = 29'b0_100110001101_110_0_100110001101;
      patterns[19567] = 29'b0_100110001101_111_0_100110001101;
      patterns[19568] = 29'b0_100110001110_000_0_100110001110;
      patterns[19569] = 29'b0_100110001110_001_0_001110100110;
      patterns[19570] = 29'b0_100110001110_010_1_001100011100;
      patterns[19571] = 29'b0_100110001110_011_0_011000111001;
      patterns[19572] = 29'b0_100110001110_100_0_010011000111;
      patterns[19573] = 29'b0_100110001110_101_1_001001100011;
      patterns[19574] = 29'b0_100110001110_110_0_100110001110;
      patterns[19575] = 29'b0_100110001110_111_0_100110001110;
      patterns[19576] = 29'b0_100110001111_000_0_100110001111;
      patterns[19577] = 29'b0_100110001111_001_0_001111100110;
      patterns[19578] = 29'b0_100110001111_010_1_001100011110;
      patterns[19579] = 29'b0_100110001111_011_0_011000111101;
      patterns[19580] = 29'b0_100110001111_100_1_010011000111;
      patterns[19581] = 29'b0_100110001111_101_1_101001100011;
      patterns[19582] = 29'b0_100110001111_110_0_100110001111;
      patterns[19583] = 29'b0_100110001111_111_0_100110001111;
      patterns[19584] = 29'b0_100110010000_000_0_100110010000;
      patterns[19585] = 29'b0_100110010000_001_0_010000100110;
      patterns[19586] = 29'b0_100110010000_010_1_001100100000;
      patterns[19587] = 29'b0_100110010000_011_0_011001000001;
      patterns[19588] = 29'b0_100110010000_100_0_010011001000;
      patterns[19589] = 29'b0_100110010000_101_0_001001100100;
      patterns[19590] = 29'b0_100110010000_110_0_100110010000;
      patterns[19591] = 29'b0_100110010000_111_0_100110010000;
      patterns[19592] = 29'b0_100110010001_000_0_100110010001;
      patterns[19593] = 29'b0_100110010001_001_0_010001100110;
      patterns[19594] = 29'b0_100110010001_010_1_001100100010;
      patterns[19595] = 29'b0_100110010001_011_0_011001000101;
      patterns[19596] = 29'b0_100110010001_100_1_010011001000;
      patterns[19597] = 29'b0_100110010001_101_0_101001100100;
      patterns[19598] = 29'b0_100110010001_110_0_100110010001;
      patterns[19599] = 29'b0_100110010001_111_0_100110010001;
      patterns[19600] = 29'b0_100110010010_000_0_100110010010;
      patterns[19601] = 29'b0_100110010010_001_0_010010100110;
      patterns[19602] = 29'b0_100110010010_010_1_001100100100;
      patterns[19603] = 29'b0_100110010010_011_0_011001001001;
      patterns[19604] = 29'b0_100110010010_100_0_010011001001;
      patterns[19605] = 29'b0_100110010010_101_1_001001100100;
      patterns[19606] = 29'b0_100110010010_110_0_100110010010;
      patterns[19607] = 29'b0_100110010010_111_0_100110010010;
      patterns[19608] = 29'b0_100110010011_000_0_100110010011;
      patterns[19609] = 29'b0_100110010011_001_0_010011100110;
      patterns[19610] = 29'b0_100110010011_010_1_001100100110;
      patterns[19611] = 29'b0_100110010011_011_0_011001001101;
      patterns[19612] = 29'b0_100110010011_100_1_010011001001;
      patterns[19613] = 29'b0_100110010011_101_1_101001100100;
      patterns[19614] = 29'b0_100110010011_110_0_100110010011;
      patterns[19615] = 29'b0_100110010011_111_0_100110010011;
      patterns[19616] = 29'b0_100110010100_000_0_100110010100;
      patterns[19617] = 29'b0_100110010100_001_0_010100100110;
      patterns[19618] = 29'b0_100110010100_010_1_001100101000;
      patterns[19619] = 29'b0_100110010100_011_0_011001010001;
      patterns[19620] = 29'b0_100110010100_100_0_010011001010;
      patterns[19621] = 29'b0_100110010100_101_0_001001100101;
      patterns[19622] = 29'b0_100110010100_110_0_100110010100;
      patterns[19623] = 29'b0_100110010100_111_0_100110010100;
      patterns[19624] = 29'b0_100110010101_000_0_100110010101;
      patterns[19625] = 29'b0_100110010101_001_0_010101100110;
      patterns[19626] = 29'b0_100110010101_010_1_001100101010;
      patterns[19627] = 29'b0_100110010101_011_0_011001010101;
      patterns[19628] = 29'b0_100110010101_100_1_010011001010;
      patterns[19629] = 29'b0_100110010101_101_0_101001100101;
      patterns[19630] = 29'b0_100110010101_110_0_100110010101;
      patterns[19631] = 29'b0_100110010101_111_0_100110010101;
      patterns[19632] = 29'b0_100110010110_000_0_100110010110;
      patterns[19633] = 29'b0_100110010110_001_0_010110100110;
      patterns[19634] = 29'b0_100110010110_010_1_001100101100;
      patterns[19635] = 29'b0_100110010110_011_0_011001011001;
      patterns[19636] = 29'b0_100110010110_100_0_010011001011;
      patterns[19637] = 29'b0_100110010110_101_1_001001100101;
      patterns[19638] = 29'b0_100110010110_110_0_100110010110;
      patterns[19639] = 29'b0_100110010110_111_0_100110010110;
      patterns[19640] = 29'b0_100110010111_000_0_100110010111;
      patterns[19641] = 29'b0_100110010111_001_0_010111100110;
      patterns[19642] = 29'b0_100110010111_010_1_001100101110;
      patterns[19643] = 29'b0_100110010111_011_0_011001011101;
      patterns[19644] = 29'b0_100110010111_100_1_010011001011;
      patterns[19645] = 29'b0_100110010111_101_1_101001100101;
      patterns[19646] = 29'b0_100110010111_110_0_100110010111;
      patterns[19647] = 29'b0_100110010111_111_0_100110010111;
      patterns[19648] = 29'b0_100110011000_000_0_100110011000;
      patterns[19649] = 29'b0_100110011000_001_0_011000100110;
      patterns[19650] = 29'b0_100110011000_010_1_001100110000;
      patterns[19651] = 29'b0_100110011000_011_0_011001100001;
      patterns[19652] = 29'b0_100110011000_100_0_010011001100;
      patterns[19653] = 29'b0_100110011000_101_0_001001100110;
      patterns[19654] = 29'b0_100110011000_110_0_100110011000;
      patterns[19655] = 29'b0_100110011000_111_0_100110011000;
      patterns[19656] = 29'b0_100110011001_000_0_100110011001;
      patterns[19657] = 29'b0_100110011001_001_0_011001100110;
      patterns[19658] = 29'b0_100110011001_010_1_001100110010;
      patterns[19659] = 29'b0_100110011001_011_0_011001100101;
      patterns[19660] = 29'b0_100110011001_100_1_010011001100;
      patterns[19661] = 29'b0_100110011001_101_0_101001100110;
      patterns[19662] = 29'b0_100110011001_110_0_100110011001;
      patterns[19663] = 29'b0_100110011001_111_0_100110011001;
      patterns[19664] = 29'b0_100110011010_000_0_100110011010;
      patterns[19665] = 29'b0_100110011010_001_0_011010100110;
      patterns[19666] = 29'b0_100110011010_010_1_001100110100;
      patterns[19667] = 29'b0_100110011010_011_0_011001101001;
      patterns[19668] = 29'b0_100110011010_100_0_010011001101;
      patterns[19669] = 29'b0_100110011010_101_1_001001100110;
      patterns[19670] = 29'b0_100110011010_110_0_100110011010;
      patterns[19671] = 29'b0_100110011010_111_0_100110011010;
      patterns[19672] = 29'b0_100110011011_000_0_100110011011;
      patterns[19673] = 29'b0_100110011011_001_0_011011100110;
      patterns[19674] = 29'b0_100110011011_010_1_001100110110;
      patterns[19675] = 29'b0_100110011011_011_0_011001101101;
      patterns[19676] = 29'b0_100110011011_100_1_010011001101;
      patterns[19677] = 29'b0_100110011011_101_1_101001100110;
      patterns[19678] = 29'b0_100110011011_110_0_100110011011;
      patterns[19679] = 29'b0_100110011011_111_0_100110011011;
      patterns[19680] = 29'b0_100110011100_000_0_100110011100;
      patterns[19681] = 29'b0_100110011100_001_0_011100100110;
      patterns[19682] = 29'b0_100110011100_010_1_001100111000;
      patterns[19683] = 29'b0_100110011100_011_0_011001110001;
      patterns[19684] = 29'b0_100110011100_100_0_010011001110;
      patterns[19685] = 29'b0_100110011100_101_0_001001100111;
      patterns[19686] = 29'b0_100110011100_110_0_100110011100;
      patterns[19687] = 29'b0_100110011100_111_0_100110011100;
      patterns[19688] = 29'b0_100110011101_000_0_100110011101;
      patterns[19689] = 29'b0_100110011101_001_0_011101100110;
      patterns[19690] = 29'b0_100110011101_010_1_001100111010;
      patterns[19691] = 29'b0_100110011101_011_0_011001110101;
      patterns[19692] = 29'b0_100110011101_100_1_010011001110;
      patterns[19693] = 29'b0_100110011101_101_0_101001100111;
      patterns[19694] = 29'b0_100110011101_110_0_100110011101;
      patterns[19695] = 29'b0_100110011101_111_0_100110011101;
      patterns[19696] = 29'b0_100110011110_000_0_100110011110;
      patterns[19697] = 29'b0_100110011110_001_0_011110100110;
      patterns[19698] = 29'b0_100110011110_010_1_001100111100;
      patterns[19699] = 29'b0_100110011110_011_0_011001111001;
      patterns[19700] = 29'b0_100110011110_100_0_010011001111;
      patterns[19701] = 29'b0_100110011110_101_1_001001100111;
      patterns[19702] = 29'b0_100110011110_110_0_100110011110;
      patterns[19703] = 29'b0_100110011110_111_0_100110011110;
      patterns[19704] = 29'b0_100110011111_000_0_100110011111;
      patterns[19705] = 29'b0_100110011111_001_0_011111100110;
      patterns[19706] = 29'b0_100110011111_010_1_001100111110;
      patterns[19707] = 29'b0_100110011111_011_0_011001111101;
      patterns[19708] = 29'b0_100110011111_100_1_010011001111;
      patterns[19709] = 29'b0_100110011111_101_1_101001100111;
      patterns[19710] = 29'b0_100110011111_110_0_100110011111;
      patterns[19711] = 29'b0_100110011111_111_0_100110011111;
      patterns[19712] = 29'b0_100110100000_000_0_100110100000;
      patterns[19713] = 29'b0_100110100000_001_0_100000100110;
      patterns[19714] = 29'b0_100110100000_010_1_001101000000;
      patterns[19715] = 29'b0_100110100000_011_0_011010000001;
      patterns[19716] = 29'b0_100110100000_100_0_010011010000;
      patterns[19717] = 29'b0_100110100000_101_0_001001101000;
      patterns[19718] = 29'b0_100110100000_110_0_100110100000;
      patterns[19719] = 29'b0_100110100000_111_0_100110100000;
      patterns[19720] = 29'b0_100110100001_000_0_100110100001;
      patterns[19721] = 29'b0_100110100001_001_0_100001100110;
      patterns[19722] = 29'b0_100110100001_010_1_001101000010;
      patterns[19723] = 29'b0_100110100001_011_0_011010000101;
      patterns[19724] = 29'b0_100110100001_100_1_010011010000;
      patterns[19725] = 29'b0_100110100001_101_0_101001101000;
      patterns[19726] = 29'b0_100110100001_110_0_100110100001;
      patterns[19727] = 29'b0_100110100001_111_0_100110100001;
      patterns[19728] = 29'b0_100110100010_000_0_100110100010;
      patterns[19729] = 29'b0_100110100010_001_0_100010100110;
      patterns[19730] = 29'b0_100110100010_010_1_001101000100;
      patterns[19731] = 29'b0_100110100010_011_0_011010001001;
      patterns[19732] = 29'b0_100110100010_100_0_010011010001;
      patterns[19733] = 29'b0_100110100010_101_1_001001101000;
      patterns[19734] = 29'b0_100110100010_110_0_100110100010;
      patterns[19735] = 29'b0_100110100010_111_0_100110100010;
      patterns[19736] = 29'b0_100110100011_000_0_100110100011;
      patterns[19737] = 29'b0_100110100011_001_0_100011100110;
      patterns[19738] = 29'b0_100110100011_010_1_001101000110;
      patterns[19739] = 29'b0_100110100011_011_0_011010001101;
      patterns[19740] = 29'b0_100110100011_100_1_010011010001;
      patterns[19741] = 29'b0_100110100011_101_1_101001101000;
      patterns[19742] = 29'b0_100110100011_110_0_100110100011;
      patterns[19743] = 29'b0_100110100011_111_0_100110100011;
      patterns[19744] = 29'b0_100110100100_000_0_100110100100;
      patterns[19745] = 29'b0_100110100100_001_0_100100100110;
      patterns[19746] = 29'b0_100110100100_010_1_001101001000;
      patterns[19747] = 29'b0_100110100100_011_0_011010010001;
      patterns[19748] = 29'b0_100110100100_100_0_010011010010;
      patterns[19749] = 29'b0_100110100100_101_0_001001101001;
      patterns[19750] = 29'b0_100110100100_110_0_100110100100;
      patterns[19751] = 29'b0_100110100100_111_0_100110100100;
      patterns[19752] = 29'b0_100110100101_000_0_100110100101;
      patterns[19753] = 29'b0_100110100101_001_0_100101100110;
      patterns[19754] = 29'b0_100110100101_010_1_001101001010;
      patterns[19755] = 29'b0_100110100101_011_0_011010010101;
      patterns[19756] = 29'b0_100110100101_100_1_010011010010;
      patterns[19757] = 29'b0_100110100101_101_0_101001101001;
      patterns[19758] = 29'b0_100110100101_110_0_100110100101;
      patterns[19759] = 29'b0_100110100101_111_0_100110100101;
      patterns[19760] = 29'b0_100110100110_000_0_100110100110;
      patterns[19761] = 29'b0_100110100110_001_0_100110100110;
      patterns[19762] = 29'b0_100110100110_010_1_001101001100;
      patterns[19763] = 29'b0_100110100110_011_0_011010011001;
      patterns[19764] = 29'b0_100110100110_100_0_010011010011;
      patterns[19765] = 29'b0_100110100110_101_1_001001101001;
      patterns[19766] = 29'b0_100110100110_110_0_100110100110;
      patterns[19767] = 29'b0_100110100110_111_0_100110100110;
      patterns[19768] = 29'b0_100110100111_000_0_100110100111;
      patterns[19769] = 29'b0_100110100111_001_0_100111100110;
      patterns[19770] = 29'b0_100110100111_010_1_001101001110;
      patterns[19771] = 29'b0_100110100111_011_0_011010011101;
      patterns[19772] = 29'b0_100110100111_100_1_010011010011;
      patterns[19773] = 29'b0_100110100111_101_1_101001101001;
      patterns[19774] = 29'b0_100110100111_110_0_100110100111;
      patterns[19775] = 29'b0_100110100111_111_0_100110100111;
      patterns[19776] = 29'b0_100110101000_000_0_100110101000;
      patterns[19777] = 29'b0_100110101000_001_0_101000100110;
      patterns[19778] = 29'b0_100110101000_010_1_001101010000;
      patterns[19779] = 29'b0_100110101000_011_0_011010100001;
      patterns[19780] = 29'b0_100110101000_100_0_010011010100;
      patterns[19781] = 29'b0_100110101000_101_0_001001101010;
      patterns[19782] = 29'b0_100110101000_110_0_100110101000;
      patterns[19783] = 29'b0_100110101000_111_0_100110101000;
      patterns[19784] = 29'b0_100110101001_000_0_100110101001;
      patterns[19785] = 29'b0_100110101001_001_0_101001100110;
      patterns[19786] = 29'b0_100110101001_010_1_001101010010;
      patterns[19787] = 29'b0_100110101001_011_0_011010100101;
      patterns[19788] = 29'b0_100110101001_100_1_010011010100;
      patterns[19789] = 29'b0_100110101001_101_0_101001101010;
      patterns[19790] = 29'b0_100110101001_110_0_100110101001;
      patterns[19791] = 29'b0_100110101001_111_0_100110101001;
      patterns[19792] = 29'b0_100110101010_000_0_100110101010;
      patterns[19793] = 29'b0_100110101010_001_0_101010100110;
      patterns[19794] = 29'b0_100110101010_010_1_001101010100;
      patterns[19795] = 29'b0_100110101010_011_0_011010101001;
      patterns[19796] = 29'b0_100110101010_100_0_010011010101;
      patterns[19797] = 29'b0_100110101010_101_1_001001101010;
      patterns[19798] = 29'b0_100110101010_110_0_100110101010;
      patterns[19799] = 29'b0_100110101010_111_0_100110101010;
      patterns[19800] = 29'b0_100110101011_000_0_100110101011;
      patterns[19801] = 29'b0_100110101011_001_0_101011100110;
      patterns[19802] = 29'b0_100110101011_010_1_001101010110;
      patterns[19803] = 29'b0_100110101011_011_0_011010101101;
      patterns[19804] = 29'b0_100110101011_100_1_010011010101;
      patterns[19805] = 29'b0_100110101011_101_1_101001101010;
      patterns[19806] = 29'b0_100110101011_110_0_100110101011;
      patterns[19807] = 29'b0_100110101011_111_0_100110101011;
      patterns[19808] = 29'b0_100110101100_000_0_100110101100;
      patterns[19809] = 29'b0_100110101100_001_0_101100100110;
      patterns[19810] = 29'b0_100110101100_010_1_001101011000;
      patterns[19811] = 29'b0_100110101100_011_0_011010110001;
      patterns[19812] = 29'b0_100110101100_100_0_010011010110;
      patterns[19813] = 29'b0_100110101100_101_0_001001101011;
      patterns[19814] = 29'b0_100110101100_110_0_100110101100;
      patterns[19815] = 29'b0_100110101100_111_0_100110101100;
      patterns[19816] = 29'b0_100110101101_000_0_100110101101;
      patterns[19817] = 29'b0_100110101101_001_0_101101100110;
      patterns[19818] = 29'b0_100110101101_010_1_001101011010;
      patterns[19819] = 29'b0_100110101101_011_0_011010110101;
      patterns[19820] = 29'b0_100110101101_100_1_010011010110;
      patterns[19821] = 29'b0_100110101101_101_0_101001101011;
      patterns[19822] = 29'b0_100110101101_110_0_100110101101;
      patterns[19823] = 29'b0_100110101101_111_0_100110101101;
      patterns[19824] = 29'b0_100110101110_000_0_100110101110;
      patterns[19825] = 29'b0_100110101110_001_0_101110100110;
      patterns[19826] = 29'b0_100110101110_010_1_001101011100;
      patterns[19827] = 29'b0_100110101110_011_0_011010111001;
      patterns[19828] = 29'b0_100110101110_100_0_010011010111;
      patterns[19829] = 29'b0_100110101110_101_1_001001101011;
      patterns[19830] = 29'b0_100110101110_110_0_100110101110;
      patterns[19831] = 29'b0_100110101110_111_0_100110101110;
      patterns[19832] = 29'b0_100110101111_000_0_100110101111;
      patterns[19833] = 29'b0_100110101111_001_0_101111100110;
      patterns[19834] = 29'b0_100110101111_010_1_001101011110;
      patterns[19835] = 29'b0_100110101111_011_0_011010111101;
      patterns[19836] = 29'b0_100110101111_100_1_010011010111;
      patterns[19837] = 29'b0_100110101111_101_1_101001101011;
      patterns[19838] = 29'b0_100110101111_110_0_100110101111;
      patterns[19839] = 29'b0_100110101111_111_0_100110101111;
      patterns[19840] = 29'b0_100110110000_000_0_100110110000;
      patterns[19841] = 29'b0_100110110000_001_0_110000100110;
      patterns[19842] = 29'b0_100110110000_010_1_001101100000;
      patterns[19843] = 29'b0_100110110000_011_0_011011000001;
      patterns[19844] = 29'b0_100110110000_100_0_010011011000;
      patterns[19845] = 29'b0_100110110000_101_0_001001101100;
      patterns[19846] = 29'b0_100110110000_110_0_100110110000;
      patterns[19847] = 29'b0_100110110000_111_0_100110110000;
      patterns[19848] = 29'b0_100110110001_000_0_100110110001;
      patterns[19849] = 29'b0_100110110001_001_0_110001100110;
      patterns[19850] = 29'b0_100110110001_010_1_001101100010;
      patterns[19851] = 29'b0_100110110001_011_0_011011000101;
      patterns[19852] = 29'b0_100110110001_100_1_010011011000;
      patterns[19853] = 29'b0_100110110001_101_0_101001101100;
      patterns[19854] = 29'b0_100110110001_110_0_100110110001;
      patterns[19855] = 29'b0_100110110001_111_0_100110110001;
      patterns[19856] = 29'b0_100110110010_000_0_100110110010;
      patterns[19857] = 29'b0_100110110010_001_0_110010100110;
      patterns[19858] = 29'b0_100110110010_010_1_001101100100;
      patterns[19859] = 29'b0_100110110010_011_0_011011001001;
      patterns[19860] = 29'b0_100110110010_100_0_010011011001;
      patterns[19861] = 29'b0_100110110010_101_1_001001101100;
      patterns[19862] = 29'b0_100110110010_110_0_100110110010;
      patterns[19863] = 29'b0_100110110010_111_0_100110110010;
      patterns[19864] = 29'b0_100110110011_000_0_100110110011;
      patterns[19865] = 29'b0_100110110011_001_0_110011100110;
      patterns[19866] = 29'b0_100110110011_010_1_001101100110;
      patterns[19867] = 29'b0_100110110011_011_0_011011001101;
      patterns[19868] = 29'b0_100110110011_100_1_010011011001;
      patterns[19869] = 29'b0_100110110011_101_1_101001101100;
      patterns[19870] = 29'b0_100110110011_110_0_100110110011;
      patterns[19871] = 29'b0_100110110011_111_0_100110110011;
      patterns[19872] = 29'b0_100110110100_000_0_100110110100;
      patterns[19873] = 29'b0_100110110100_001_0_110100100110;
      patterns[19874] = 29'b0_100110110100_010_1_001101101000;
      patterns[19875] = 29'b0_100110110100_011_0_011011010001;
      patterns[19876] = 29'b0_100110110100_100_0_010011011010;
      patterns[19877] = 29'b0_100110110100_101_0_001001101101;
      patterns[19878] = 29'b0_100110110100_110_0_100110110100;
      patterns[19879] = 29'b0_100110110100_111_0_100110110100;
      patterns[19880] = 29'b0_100110110101_000_0_100110110101;
      patterns[19881] = 29'b0_100110110101_001_0_110101100110;
      patterns[19882] = 29'b0_100110110101_010_1_001101101010;
      patterns[19883] = 29'b0_100110110101_011_0_011011010101;
      patterns[19884] = 29'b0_100110110101_100_1_010011011010;
      patterns[19885] = 29'b0_100110110101_101_0_101001101101;
      patterns[19886] = 29'b0_100110110101_110_0_100110110101;
      patterns[19887] = 29'b0_100110110101_111_0_100110110101;
      patterns[19888] = 29'b0_100110110110_000_0_100110110110;
      patterns[19889] = 29'b0_100110110110_001_0_110110100110;
      patterns[19890] = 29'b0_100110110110_010_1_001101101100;
      patterns[19891] = 29'b0_100110110110_011_0_011011011001;
      patterns[19892] = 29'b0_100110110110_100_0_010011011011;
      patterns[19893] = 29'b0_100110110110_101_1_001001101101;
      patterns[19894] = 29'b0_100110110110_110_0_100110110110;
      patterns[19895] = 29'b0_100110110110_111_0_100110110110;
      patterns[19896] = 29'b0_100110110111_000_0_100110110111;
      patterns[19897] = 29'b0_100110110111_001_0_110111100110;
      patterns[19898] = 29'b0_100110110111_010_1_001101101110;
      patterns[19899] = 29'b0_100110110111_011_0_011011011101;
      patterns[19900] = 29'b0_100110110111_100_1_010011011011;
      patterns[19901] = 29'b0_100110110111_101_1_101001101101;
      patterns[19902] = 29'b0_100110110111_110_0_100110110111;
      patterns[19903] = 29'b0_100110110111_111_0_100110110111;
      patterns[19904] = 29'b0_100110111000_000_0_100110111000;
      patterns[19905] = 29'b0_100110111000_001_0_111000100110;
      patterns[19906] = 29'b0_100110111000_010_1_001101110000;
      patterns[19907] = 29'b0_100110111000_011_0_011011100001;
      patterns[19908] = 29'b0_100110111000_100_0_010011011100;
      patterns[19909] = 29'b0_100110111000_101_0_001001101110;
      patterns[19910] = 29'b0_100110111000_110_0_100110111000;
      patterns[19911] = 29'b0_100110111000_111_0_100110111000;
      patterns[19912] = 29'b0_100110111001_000_0_100110111001;
      patterns[19913] = 29'b0_100110111001_001_0_111001100110;
      patterns[19914] = 29'b0_100110111001_010_1_001101110010;
      patterns[19915] = 29'b0_100110111001_011_0_011011100101;
      patterns[19916] = 29'b0_100110111001_100_1_010011011100;
      patterns[19917] = 29'b0_100110111001_101_0_101001101110;
      patterns[19918] = 29'b0_100110111001_110_0_100110111001;
      patterns[19919] = 29'b0_100110111001_111_0_100110111001;
      patterns[19920] = 29'b0_100110111010_000_0_100110111010;
      patterns[19921] = 29'b0_100110111010_001_0_111010100110;
      patterns[19922] = 29'b0_100110111010_010_1_001101110100;
      patterns[19923] = 29'b0_100110111010_011_0_011011101001;
      patterns[19924] = 29'b0_100110111010_100_0_010011011101;
      patterns[19925] = 29'b0_100110111010_101_1_001001101110;
      patterns[19926] = 29'b0_100110111010_110_0_100110111010;
      patterns[19927] = 29'b0_100110111010_111_0_100110111010;
      patterns[19928] = 29'b0_100110111011_000_0_100110111011;
      patterns[19929] = 29'b0_100110111011_001_0_111011100110;
      patterns[19930] = 29'b0_100110111011_010_1_001101110110;
      patterns[19931] = 29'b0_100110111011_011_0_011011101101;
      patterns[19932] = 29'b0_100110111011_100_1_010011011101;
      patterns[19933] = 29'b0_100110111011_101_1_101001101110;
      patterns[19934] = 29'b0_100110111011_110_0_100110111011;
      patterns[19935] = 29'b0_100110111011_111_0_100110111011;
      patterns[19936] = 29'b0_100110111100_000_0_100110111100;
      patterns[19937] = 29'b0_100110111100_001_0_111100100110;
      patterns[19938] = 29'b0_100110111100_010_1_001101111000;
      patterns[19939] = 29'b0_100110111100_011_0_011011110001;
      patterns[19940] = 29'b0_100110111100_100_0_010011011110;
      patterns[19941] = 29'b0_100110111100_101_0_001001101111;
      patterns[19942] = 29'b0_100110111100_110_0_100110111100;
      patterns[19943] = 29'b0_100110111100_111_0_100110111100;
      patterns[19944] = 29'b0_100110111101_000_0_100110111101;
      patterns[19945] = 29'b0_100110111101_001_0_111101100110;
      patterns[19946] = 29'b0_100110111101_010_1_001101111010;
      patterns[19947] = 29'b0_100110111101_011_0_011011110101;
      patterns[19948] = 29'b0_100110111101_100_1_010011011110;
      patterns[19949] = 29'b0_100110111101_101_0_101001101111;
      patterns[19950] = 29'b0_100110111101_110_0_100110111101;
      patterns[19951] = 29'b0_100110111101_111_0_100110111101;
      patterns[19952] = 29'b0_100110111110_000_0_100110111110;
      patterns[19953] = 29'b0_100110111110_001_0_111110100110;
      patterns[19954] = 29'b0_100110111110_010_1_001101111100;
      patterns[19955] = 29'b0_100110111110_011_0_011011111001;
      patterns[19956] = 29'b0_100110111110_100_0_010011011111;
      patterns[19957] = 29'b0_100110111110_101_1_001001101111;
      patterns[19958] = 29'b0_100110111110_110_0_100110111110;
      patterns[19959] = 29'b0_100110111110_111_0_100110111110;
      patterns[19960] = 29'b0_100110111111_000_0_100110111111;
      patterns[19961] = 29'b0_100110111111_001_0_111111100110;
      patterns[19962] = 29'b0_100110111111_010_1_001101111110;
      patterns[19963] = 29'b0_100110111111_011_0_011011111101;
      patterns[19964] = 29'b0_100110111111_100_1_010011011111;
      patterns[19965] = 29'b0_100110111111_101_1_101001101111;
      patterns[19966] = 29'b0_100110111111_110_0_100110111111;
      patterns[19967] = 29'b0_100110111111_111_0_100110111111;
      patterns[19968] = 29'b0_100111000000_000_0_100111000000;
      patterns[19969] = 29'b0_100111000000_001_0_000000100111;
      patterns[19970] = 29'b0_100111000000_010_1_001110000000;
      patterns[19971] = 29'b0_100111000000_011_0_011100000001;
      patterns[19972] = 29'b0_100111000000_100_0_010011100000;
      patterns[19973] = 29'b0_100111000000_101_0_001001110000;
      patterns[19974] = 29'b0_100111000000_110_0_100111000000;
      patterns[19975] = 29'b0_100111000000_111_0_100111000000;
      patterns[19976] = 29'b0_100111000001_000_0_100111000001;
      patterns[19977] = 29'b0_100111000001_001_0_000001100111;
      patterns[19978] = 29'b0_100111000001_010_1_001110000010;
      patterns[19979] = 29'b0_100111000001_011_0_011100000101;
      patterns[19980] = 29'b0_100111000001_100_1_010011100000;
      patterns[19981] = 29'b0_100111000001_101_0_101001110000;
      patterns[19982] = 29'b0_100111000001_110_0_100111000001;
      patterns[19983] = 29'b0_100111000001_111_0_100111000001;
      patterns[19984] = 29'b0_100111000010_000_0_100111000010;
      patterns[19985] = 29'b0_100111000010_001_0_000010100111;
      patterns[19986] = 29'b0_100111000010_010_1_001110000100;
      patterns[19987] = 29'b0_100111000010_011_0_011100001001;
      patterns[19988] = 29'b0_100111000010_100_0_010011100001;
      patterns[19989] = 29'b0_100111000010_101_1_001001110000;
      patterns[19990] = 29'b0_100111000010_110_0_100111000010;
      patterns[19991] = 29'b0_100111000010_111_0_100111000010;
      patterns[19992] = 29'b0_100111000011_000_0_100111000011;
      patterns[19993] = 29'b0_100111000011_001_0_000011100111;
      patterns[19994] = 29'b0_100111000011_010_1_001110000110;
      patterns[19995] = 29'b0_100111000011_011_0_011100001101;
      patterns[19996] = 29'b0_100111000011_100_1_010011100001;
      patterns[19997] = 29'b0_100111000011_101_1_101001110000;
      patterns[19998] = 29'b0_100111000011_110_0_100111000011;
      patterns[19999] = 29'b0_100111000011_111_0_100111000011;
      patterns[20000] = 29'b0_100111000100_000_0_100111000100;
      patterns[20001] = 29'b0_100111000100_001_0_000100100111;
      patterns[20002] = 29'b0_100111000100_010_1_001110001000;
      patterns[20003] = 29'b0_100111000100_011_0_011100010001;
      patterns[20004] = 29'b0_100111000100_100_0_010011100010;
      patterns[20005] = 29'b0_100111000100_101_0_001001110001;
      patterns[20006] = 29'b0_100111000100_110_0_100111000100;
      patterns[20007] = 29'b0_100111000100_111_0_100111000100;
      patterns[20008] = 29'b0_100111000101_000_0_100111000101;
      patterns[20009] = 29'b0_100111000101_001_0_000101100111;
      patterns[20010] = 29'b0_100111000101_010_1_001110001010;
      patterns[20011] = 29'b0_100111000101_011_0_011100010101;
      patterns[20012] = 29'b0_100111000101_100_1_010011100010;
      patterns[20013] = 29'b0_100111000101_101_0_101001110001;
      patterns[20014] = 29'b0_100111000101_110_0_100111000101;
      patterns[20015] = 29'b0_100111000101_111_0_100111000101;
      patterns[20016] = 29'b0_100111000110_000_0_100111000110;
      patterns[20017] = 29'b0_100111000110_001_0_000110100111;
      patterns[20018] = 29'b0_100111000110_010_1_001110001100;
      patterns[20019] = 29'b0_100111000110_011_0_011100011001;
      patterns[20020] = 29'b0_100111000110_100_0_010011100011;
      patterns[20021] = 29'b0_100111000110_101_1_001001110001;
      patterns[20022] = 29'b0_100111000110_110_0_100111000110;
      patterns[20023] = 29'b0_100111000110_111_0_100111000110;
      patterns[20024] = 29'b0_100111000111_000_0_100111000111;
      patterns[20025] = 29'b0_100111000111_001_0_000111100111;
      patterns[20026] = 29'b0_100111000111_010_1_001110001110;
      patterns[20027] = 29'b0_100111000111_011_0_011100011101;
      patterns[20028] = 29'b0_100111000111_100_1_010011100011;
      patterns[20029] = 29'b0_100111000111_101_1_101001110001;
      patterns[20030] = 29'b0_100111000111_110_0_100111000111;
      patterns[20031] = 29'b0_100111000111_111_0_100111000111;
      patterns[20032] = 29'b0_100111001000_000_0_100111001000;
      patterns[20033] = 29'b0_100111001000_001_0_001000100111;
      patterns[20034] = 29'b0_100111001000_010_1_001110010000;
      patterns[20035] = 29'b0_100111001000_011_0_011100100001;
      patterns[20036] = 29'b0_100111001000_100_0_010011100100;
      patterns[20037] = 29'b0_100111001000_101_0_001001110010;
      patterns[20038] = 29'b0_100111001000_110_0_100111001000;
      patterns[20039] = 29'b0_100111001000_111_0_100111001000;
      patterns[20040] = 29'b0_100111001001_000_0_100111001001;
      patterns[20041] = 29'b0_100111001001_001_0_001001100111;
      patterns[20042] = 29'b0_100111001001_010_1_001110010010;
      patterns[20043] = 29'b0_100111001001_011_0_011100100101;
      patterns[20044] = 29'b0_100111001001_100_1_010011100100;
      patterns[20045] = 29'b0_100111001001_101_0_101001110010;
      patterns[20046] = 29'b0_100111001001_110_0_100111001001;
      patterns[20047] = 29'b0_100111001001_111_0_100111001001;
      patterns[20048] = 29'b0_100111001010_000_0_100111001010;
      patterns[20049] = 29'b0_100111001010_001_0_001010100111;
      patterns[20050] = 29'b0_100111001010_010_1_001110010100;
      patterns[20051] = 29'b0_100111001010_011_0_011100101001;
      patterns[20052] = 29'b0_100111001010_100_0_010011100101;
      patterns[20053] = 29'b0_100111001010_101_1_001001110010;
      patterns[20054] = 29'b0_100111001010_110_0_100111001010;
      patterns[20055] = 29'b0_100111001010_111_0_100111001010;
      patterns[20056] = 29'b0_100111001011_000_0_100111001011;
      patterns[20057] = 29'b0_100111001011_001_0_001011100111;
      patterns[20058] = 29'b0_100111001011_010_1_001110010110;
      patterns[20059] = 29'b0_100111001011_011_0_011100101101;
      patterns[20060] = 29'b0_100111001011_100_1_010011100101;
      patterns[20061] = 29'b0_100111001011_101_1_101001110010;
      patterns[20062] = 29'b0_100111001011_110_0_100111001011;
      patterns[20063] = 29'b0_100111001011_111_0_100111001011;
      patterns[20064] = 29'b0_100111001100_000_0_100111001100;
      patterns[20065] = 29'b0_100111001100_001_0_001100100111;
      patterns[20066] = 29'b0_100111001100_010_1_001110011000;
      patterns[20067] = 29'b0_100111001100_011_0_011100110001;
      patterns[20068] = 29'b0_100111001100_100_0_010011100110;
      patterns[20069] = 29'b0_100111001100_101_0_001001110011;
      patterns[20070] = 29'b0_100111001100_110_0_100111001100;
      patterns[20071] = 29'b0_100111001100_111_0_100111001100;
      patterns[20072] = 29'b0_100111001101_000_0_100111001101;
      patterns[20073] = 29'b0_100111001101_001_0_001101100111;
      patterns[20074] = 29'b0_100111001101_010_1_001110011010;
      patterns[20075] = 29'b0_100111001101_011_0_011100110101;
      patterns[20076] = 29'b0_100111001101_100_1_010011100110;
      patterns[20077] = 29'b0_100111001101_101_0_101001110011;
      patterns[20078] = 29'b0_100111001101_110_0_100111001101;
      patterns[20079] = 29'b0_100111001101_111_0_100111001101;
      patterns[20080] = 29'b0_100111001110_000_0_100111001110;
      patterns[20081] = 29'b0_100111001110_001_0_001110100111;
      patterns[20082] = 29'b0_100111001110_010_1_001110011100;
      patterns[20083] = 29'b0_100111001110_011_0_011100111001;
      patterns[20084] = 29'b0_100111001110_100_0_010011100111;
      patterns[20085] = 29'b0_100111001110_101_1_001001110011;
      patterns[20086] = 29'b0_100111001110_110_0_100111001110;
      patterns[20087] = 29'b0_100111001110_111_0_100111001110;
      patterns[20088] = 29'b0_100111001111_000_0_100111001111;
      patterns[20089] = 29'b0_100111001111_001_0_001111100111;
      patterns[20090] = 29'b0_100111001111_010_1_001110011110;
      patterns[20091] = 29'b0_100111001111_011_0_011100111101;
      patterns[20092] = 29'b0_100111001111_100_1_010011100111;
      patterns[20093] = 29'b0_100111001111_101_1_101001110011;
      patterns[20094] = 29'b0_100111001111_110_0_100111001111;
      patterns[20095] = 29'b0_100111001111_111_0_100111001111;
      patterns[20096] = 29'b0_100111010000_000_0_100111010000;
      patterns[20097] = 29'b0_100111010000_001_0_010000100111;
      patterns[20098] = 29'b0_100111010000_010_1_001110100000;
      patterns[20099] = 29'b0_100111010000_011_0_011101000001;
      patterns[20100] = 29'b0_100111010000_100_0_010011101000;
      patterns[20101] = 29'b0_100111010000_101_0_001001110100;
      patterns[20102] = 29'b0_100111010000_110_0_100111010000;
      patterns[20103] = 29'b0_100111010000_111_0_100111010000;
      patterns[20104] = 29'b0_100111010001_000_0_100111010001;
      patterns[20105] = 29'b0_100111010001_001_0_010001100111;
      patterns[20106] = 29'b0_100111010001_010_1_001110100010;
      patterns[20107] = 29'b0_100111010001_011_0_011101000101;
      patterns[20108] = 29'b0_100111010001_100_1_010011101000;
      patterns[20109] = 29'b0_100111010001_101_0_101001110100;
      patterns[20110] = 29'b0_100111010001_110_0_100111010001;
      patterns[20111] = 29'b0_100111010001_111_0_100111010001;
      patterns[20112] = 29'b0_100111010010_000_0_100111010010;
      patterns[20113] = 29'b0_100111010010_001_0_010010100111;
      patterns[20114] = 29'b0_100111010010_010_1_001110100100;
      patterns[20115] = 29'b0_100111010010_011_0_011101001001;
      patterns[20116] = 29'b0_100111010010_100_0_010011101001;
      patterns[20117] = 29'b0_100111010010_101_1_001001110100;
      patterns[20118] = 29'b0_100111010010_110_0_100111010010;
      patterns[20119] = 29'b0_100111010010_111_0_100111010010;
      patterns[20120] = 29'b0_100111010011_000_0_100111010011;
      patterns[20121] = 29'b0_100111010011_001_0_010011100111;
      patterns[20122] = 29'b0_100111010011_010_1_001110100110;
      patterns[20123] = 29'b0_100111010011_011_0_011101001101;
      patterns[20124] = 29'b0_100111010011_100_1_010011101001;
      patterns[20125] = 29'b0_100111010011_101_1_101001110100;
      patterns[20126] = 29'b0_100111010011_110_0_100111010011;
      patterns[20127] = 29'b0_100111010011_111_0_100111010011;
      patterns[20128] = 29'b0_100111010100_000_0_100111010100;
      patterns[20129] = 29'b0_100111010100_001_0_010100100111;
      patterns[20130] = 29'b0_100111010100_010_1_001110101000;
      patterns[20131] = 29'b0_100111010100_011_0_011101010001;
      patterns[20132] = 29'b0_100111010100_100_0_010011101010;
      patterns[20133] = 29'b0_100111010100_101_0_001001110101;
      patterns[20134] = 29'b0_100111010100_110_0_100111010100;
      patterns[20135] = 29'b0_100111010100_111_0_100111010100;
      patterns[20136] = 29'b0_100111010101_000_0_100111010101;
      patterns[20137] = 29'b0_100111010101_001_0_010101100111;
      patterns[20138] = 29'b0_100111010101_010_1_001110101010;
      patterns[20139] = 29'b0_100111010101_011_0_011101010101;
      patterns[20140] = 29'b0_100111010101_100_1_010011101010;
      patterns[20141] = 29'b0_100111010101_101_0_101001110101;
      patterns[20142] = 29'b0_100111010101_110_0_100111010101;
      patterns[20143] = 29'b0_100111010101_111_0_100111010101;
      patterns[20144] = 29'b0_100111010110_000_0_100111010110;
      patterns[20145] = 29'b0_100111010110_001_0_010110100111;
      patterns[20146] = 29'b0_100111010110_010_1_001110101100;
      patterns[20147] = 29'b0_100111010110_011_0_011101011001;
      patterns[20148] = 29'b0_100111010110_100_0_010011101011;
      patterns[20149] = 29'b0_100111010110_101_1_001001110101;
      patterns[20150] = 29'b0_100111010110_110_0_100111010110;
      patterns[20151] = 29'b0_100111010110_111_0_100111010110;
      patterns[20152] = 29'b0_100111010111_000_0_100111010111;
      patterns[20153] = 29'b0_100111010111_001_0_010111100111;
      patterns[20154] = 29'b0_100111010111_010_1_001110101110;
      patterns[20155] = 29'b0_100111010111_011_0_011101011101;
      patterns[20156] = 29'b0_100111010111_100_1_010011101011;
      patterns[20157] = 29'b0_100111010111_101_1_101001110101;
      patterns[20158] = 29'b0_100111010111_110_0_100111010111;
      patterns[20159] = 29'b0_100111010111_111_0_100111010111;
      patterns[20160] = 29'b0_100111011000_000_0_100111011000;
      patterns[20161] = 29'b0_100111011000_001_0_011000100111;
      patterns[20162] = 29'b0_100111011000_010_1_001110110000;
      patterns[20163] = 29'b0_100111011000_011_0_011101100001;
      patterns[20164] = 29'b0_100111011000_100_0_010011101100;
      patterns[20165] = 29'b0_100111011000_101_0_001001110110;
      patterns[20166] = 29'b0_100111011000_110_0_100111011000;
      patterns[20167] = 29'b0_100111011000_111_0_100111011000;
      patterns[20168] = 29'b0_100111011001_000_0_100111011001;
      patterns[20169] = 29'b0_100111011001_001_0_011001100111;
      patterns[20170] = 29'b0_100111011001_010_1_001110110010;
      patterns[20171] = 29'b0_100111011001_011_0_011101100101;
      patterns[20172] = 29'b0_100111011001_100_1_010011101100;
      patterns[20173] = 29'b0_100111011001_101_0_101001110110;
      patterns[20174] = 29'b0_100111011001_110_0_100111011001;
      patterns[20175] = 29'b0_100111011001_111_0_100111011001;
      patterns[20176] = 29'b0_100111011010_000_0_100111011010;
      patterns[20177] = 29'b0_100111011010_001_0_011010100111;
      patterns[20178] = 29'b0_100111011010_010_1_001110110100;
      patterns[20179] = 29'b0_100111011010_011_0_011101101001;
      patterns[20180] = 29'b0_100111011010_100_0_010011101101;
      patterns[20181] = 29'b0_100111011010_101_1_001001110110;
      patterns[20182] = 29'b0_100111011010_110_0_100111011010;
      patterns[20183] = 29'b0_100111011010_111_0_100111011010;
      patterns[20184] = 29'b0_100111011011_000_0_100111011011;
      patterns[20185] = 29'b0_100111011011_001_0_011011100111;
      patterns[20186] = 29'b0_100111011011_010_1_001110110110;
      patterns[20187] = 29'b0_100111011011_011_0_011101101101;
      patterns[20188] = 29'b0_100111011011_100_1_010011101101;
      patterns[20189] = 29'b0_100111011011_101_1_101001110110;
      patterns[20190] = 29'b0_100111011011_110_0_100111011011;
      patterns[20191] = 29'b0_100111011011_111_0_100111011011;
      patterns[20192] = 29'b0_100111011100_000_0_100111011100;
      patterns[20193] = 29'b0_100111011100_001_0_011100100111;
      patterns[20194] = 29'b0_100111011100_010_1_001110111000;
      patterns[20195] = 29'b0_100111011100_011_0_011101110001;
      patterns[20196] = 29'b0_100111011100_100_0_010011101110;
      patterns[20197] = 29'b0_100111011100_101_0_001001110111;
      patterns[20198] = 29'b0_100111011100_110_0_100111011100;
      patterns[20199] = 29'b0_100111011100_111_0_100111011100;
      patterns[20200] = 29'b0_100111011101_000_0_100111011101;
      patterns[20201] = 29'b0_100111011101_001_0_011101100111;
      patterns[20202] = 29'b0_100111011101_010_1_001110111010;
      patterns[20203] = 29'b0_100111011101_011_0_011101110101;
      patterns[20204] = 29'b0_100111011101_100_1_010011101110;
      patterns[20205] = 29'b0_100111011101_101_0_101001110111;
      patterns[20206] = 29'b0_100111011101_110_0_100111011101;
      patterns[20207] = 29'b0_100111011101_111_0_100111011101;
      patterns[20208] = 29'b0_100111011110_000_0_100111011110;
      patterns[20209] = 29'b0_100111011110_001_0_011110100111;
      patterns[20210] = 29'b0_100111011110_010_1_001110111100;
      patterns[20211] = 29'b0_100111011110_011_0_011101111001;
      patterns[20212] = 29'b0_100111011110_100_0_010011101111;
      patterns[20213] = 29'b0_100111011110_101_1_001001110111;
      patterns[20214] = 29'b0_100111011110_110_0_100111011110;
      patterns[20215] = 29'b0_100111011110_111_0_100111011110;
      patterns[20216] = 29'b0_100111011111_000_0_100111011111;
      patterns[20217] = 29'b0_100111011111_001_0_011111100111;
      patterns[20218] = 29'b0_100111011111_010_1_001110111110;
      patterns[20219] = 29'b0_100111011111_011_0_011101111101;
      patterns[20220] = 29'b0_100111011111_100_1_010011101111;
      patterns[20221] = 29'b0_100111011111_101_1_101001110111;
      patterns[20222] = 29'b0_100111011111_110_0_100111011111;
      patterns[20223] = 29'b0_100111011111_111_0_100111011111;
      patterns[20224] = 29'b0_100111100000_000_0_100111100000;
      patterns[20225] = 29'b0_100111100000_001_0_100000100111;
      patterns[20226] = 29'b0_100111100000_010_1_001111000000;
      patterns[20227] = 29'b0_100111100000_011_0_011110000001;
      patterns[20228] = 29'b0_100111100000_100_0_010011110000;
      patterns[20229] = 29'b0_100111100000_101_0_001001111000;
      patterns[20230] = 29'b0_100111100000_110_0_100111100000;
      patterns[20231] = 29'b0_100111100000_111_0_100111100000;
      patterns[20232] = 29'b0_100111100001_000_0_100111100001;
      patterns[20233] = 29'b0_100111100001_001_0_100001100111;
      patterns[20234] = 29'b0_100111100001_010_1_001111000010;
      patterns[20235] = 29'b0_100111100001_011_0_011110000101;
      patterns[20236] = 29'b0_100111100001_100_1_010011110000;
      patterns[20237] = 29'b0_100111100001_101_0_101001111000;
      patterns[20238] = 29'b0_100111100001_110_0_100111100001;
      patterns[20239] = 29'b0_100111100001_111_0_100111100001;
      patterns[20240] = 29'b0_100111100010_000_0_100111100010;
      patterns[20241] = 29'b0_100111100010_001_0_100010100111;
      patterns[20242] = 29'b0_100111100010_010_1_001111000100;
      patterns[20243] = 29'b0_100111100010_011_0_011110001001;
      patterns[20244] = 29'b0_100111100010_100_0_010011110001;
      patterns[20245] = 29'b0_100111100010_101_1_001001111000;
      patterns[20246] = 29'b0_100111100010_110_0_100111100010;
      patterns[20247] = 29'b0_100111100010_111_0_100111100010;
      patterns[20248] = 29'b0_100111100011_000_0_100111100011;
      patterns[20249] = 29'b0_100111100011_001_0_100011100111;
      patterns[20250] = 29'b0_100111100011_010_1_001111000110;
      patterns[20251] = 29'b0_100111100011_011_0_011110001101;
      patterns[20252] = 29'b0_100111100011_100_1_010011110001;
      patterns[20253] = 29'b0_100111100011_101_1_101001111000;
      patterns[20254] = 29'b0_100111100011_110_0_100111100011;
      patterns[20255] = 29'b0_100111100011_111_0_100111100011;
      patterns[20256] = 29'b0_100111100100_000_0_100111100100;
      patterns[20257] = 29'b0_100111100100_001_0_100100100111;
      patterns[20258] = 29'b0_100111100100_010_1_001111001000;
      patterns[20259] = 29'b0_100111100100_011_0_011110010001;
      patterns[20260] = 29'b0_100111100100_100_0_010011110010;
      patterns[20261] = 29'b0_100111100100_101_0_001001111001;
      patterns[20262] = 29'b0_100111100100_110_0_100111100100;
      patterns[20263] = 29'b0_100111100100_111_0_100111100100;
      patterns[20264] = 29'b0_100111100101_000_0_100111100101;
      patterns[20265] = 29'b0_100111100101_001_0_100101100111;
      patterns[20266] = 29'b0_100111100101_010_1_001111001010;
      patterns[20267] = 29'b0_100111100101_011_0_011110010101;
      patterns[20268] = 29'b0_100111100101_100_1_010011110010;
      patterns[20269] = 29'b0_100111100101_101_0_101001111001;
      patterns[20270] = 29'b0_100111100101_110_0_100111100101;
      patterns[20271] = 29'b0_100111100101_111_0_100111100101;
      patterns[20272] = 29'b0_100111100110_000_0_100111100110;
      patterns[20273] = 29'b0_100111100110_001_0_100110100111;
      patterns[20274] = 29'b0_100111100110_010_1_001111001100;
      patterns[20275] = 29'b0_100111100110_011_0_011110011001;
      patterns[20276] = 29'b0_100111100110_100_0_010011110011;
      patterns[20277] = 29'b0_100111100110_101_1_001001111001;
      patterns[20278] = 29'b0_100111100110_110_0_100111100110;
      patterns[20279] = 29'b0_100111100110_111_0_100111100110;
      patterns[20280] = 29'b0_100111100111_000_0_100111100111;
      patterns[20281] = 29'b0_100111100111_001_0_100111100111;
      patterns[20282] = 29'b0_100111100111_010_1_001111001110;
      patterns[20283] = 29'b0_100111100111_011_0_011110011101;
      patterns[20284] = 29'b0_100111100111_100_1_010011110011;
      patterns[20285] = 29'b0_100111100111_101_1_101001111001;
      patterns[20286] = 29'b0_100111100111_110_0_100111100111;
      patterns[20287] = 29'b0_100111100111_111_0_100111100111;
      patterns[20288] = 29'b0_100111101000_000_0_100111101000;
      patterns[20289] = 29'b0_100111101000_001_0_101000100111;
      patterns[20290] = 29'b0_100111101000_010_1_001111010000;
      patterns[20291] = 29'b0_100111101000_011_0_011110100001;
      patterns[20292] = 29'b0_100111101000_100_0_010011110100;
      patterns[20293] = 29'b0_100111101000_101_0_001001111010;
      patterns[20294] = 29'b0_100111101000_110_0_100111101000;
      patterns[20295] = 29'b0_100111101000_111_0_100111101000;
      patterns[20296] = 29'b0_100111101001_000_0_100111101001;
      patterns[20297] = 29'b0_100111101001_001_0_101001100111;
      patterns[20298] = 29'b0_100111101001_010_1_001111010010;
      patterns[20299] = 29'b0_100111101001_011_0_011110100101;
      patterns[20300] = 29'b0_100111101001_100_1_010011110100;
      patterns[20301] = 29'b0_100111101001_101_0_101001111010;
      patterns[20302] = 29'b0_100111101001_110_0_100111101001;
      patterns[20303] = 29'b0_100111101001_111_0_100111101001;
      patterns[20304] = 29'b0_100111101010_000_0_100111101010;
      patterns[20305] = 29'b0_100111101010_001_0_101010100111;
      patterns[20306] = 29'b0_100111101010_010_1_001111010100;
      patterns[20307] = 29'b0_100111101010_011_0_011110101001;
      patterns[20308] = 29'b0_100111101010_100_0_010011110101;
      patterns[20309] = 29'b0_100111101010_101_1_001001111010;
      patterns[20310] = 29'b0_100111101010_110_0_100111101010;
      patterns[20311] = 29'b0_100111101010_111_0_100111101010;
      patterns[20312] = 29'b0_100111101011_000_0_100111101011;
      patterns[20313] = 29'b0_100111101011_001_0_101011100111;
      patterns[20314] = 29'b0_100111101011_010_1_001111010110;
      patterns[20315] = 29'b0_100111101011_011_0_011110101101;
      patterns[20316] = 29'b0_100111101011_100_1_010011110101;
      patterns[20317] = 29'b0_100111101011_101_1_101001111010;
      patterns[20318] = 29'b0_100111101011_110_0_100111101011;
      patterns[20319] = 29'b0_100111101011_111_0_100111101011;
      patterns[20320] = 29'b0_100111101100_000_0_100111101100;
      patterns[20321] = 29'b0_100111101100_001_0_101100100111;
      patterns[20322] = 29'b0_100111101100_010_1_001111011000;
      patterns[20323] = 29'b0_100111101100_011_0_011110110001;
      patterns[20324] = 29'b0_100111101100_100_0_010011110110;
      patterns[20325] = 29'b0_100111101100_101_0_001001111011;
      patterns[20326] = 29'b0_100111101100_110_0_100111101100;
      patterns[20327] = 29'b0_100111101100_111_0_100111101100;
      patterns[20328] = 29'b0_100111101101_000_0_100111101101;
      patterns[20329] = 29'b0_100111101101_001_0_101101100111;
      patterns[20330] = 29'b0_100111101101_010_1_001111011010;
      patterns[20331] = 29'b0_100111101101_011_0_011110110101;
      patterns[20332] = 29'b0_100111101101_100_1_010011110110;
      patterns[20333] = 29'b0_100111101101_101_0_101001111011;
      patterns[20334] = 29'b0_100111101101_110_0_100111101101;
      patterns[20335] = 29'b0_100111101101_111_0_100111101101;
      patterns[20336] = 29'b0_100111101110_000_0_100111101110;
      patterns[20337] = 29'b0_100111101110_001_0_101110100111;
      patterns[20338] = 29'b0_100111101110_010_1_001111011100;
      patterns[20339] = 29'b0_100111101110_011_0_011110111001;
      patterns[20340] = 29'b0_100111101110_100_0_010011110111;
      patterns[20341] = 29'b0_100111101110_101_1_001001111011;
      patterns[20342] = 29'b0_100111101110_110_0_100111101110;
      patterns[20343] = 29'b0_100111101110_111_0_100111101110;
      patterns[20344] = 29'b0_100111101111_000_0_100111101111;
      patterns[20345] = 29'b0_100111101111_001_0_101111100111;
      patterns[20346] = 29'b0_100111101111_010_1_001111011110;
      patterns[20347] = 29'b0_100111101111_011_0_011110111101;
      patterns[20348] = 29'b0_100111101111_100_1_010011110111;
      patterns[20349] = 29'b0_100111101111_101_1_101001111011;
      patterns[20350] = 29'b0_100111101111_110_0_100111101111;
      patterns[20351] = 29'b0_100111101111_111_0_100111101111;
      patterns[20352] = 29'b0_100111110000_000_0_100111110000;
      patterns[20353] = 29'b0_100111110000_001_0_110000100111;
      patterns[20354] = 29'b0_100111110000_010_1_001111100000;
      patterns[20355] = 29'b0_100111110000_011_0_011111000001;
      patterns[20356] = 29'b0_100111110000_100_0_010011111000;
      patterns[20357] = 29'b0_100111110000_101_0_001001111100;
      patterns[20358] = 29'b0_100111110000_110_0_100111110000;
      patterns[20359] = 29'b0_100111110000_111_0_100111110000;
      patterns[20360] = 29'b0_100111110001_000_0_100111110001;
      patterns[20361] = 29'b0_100111110001_001_0_110001100111;
      patterns[20362] = 29'b0_100111110001_010_1_001111100010;
      patterns[20363] = 29'b0_100111110001_011_0_011111000101;
      patterns[20364] = 29'b0_100111110001_100_1_010011111000;
      patterns[20365] = 29'b0_100111110001_101_0_101001111100;
      patterns[20366] = 29'b0_100111110001_110_0_100111110001;
      patterns[20367] = 29'b0_100111110001_111_0_100111110001;
      patterns[20368] = 29'b0_100111110010_000_0_100111110010;
      patterns[20369] = 29'b0_100111110010_001_0_110010100111;
      patterns[20370] = 29'b0_100111110010_010_1_001111100100;
      patterns[20371] = 29'b0_100111110010_011_0_011111001001;
      patterns[20372] = 29'b0_100111110010_100_0_010011111001;
      patterns[20373] = 29'b0_100111110010_101_1_001001111100;
      patterns[20374] = 29'b0_100111110010_110_0_100111110010;
      patterns[20375] = 29'b0_100111110010_111_0_100111110010;
      patterns[20376] = 29'b0_100111110011_000_0_100111110011;
      patterns[20377] = 29'b0_100111110011_001_0_110011100111;
      patterns[20378] = 29'b0_100111110011_010_1_001111100110;
      patterns[20379] = 29'b0_100111110011_011_0_011111001101;
      patterns[20380] = 29'b0_100111110011_100_1_010011111001;
      patterns[20381] = 29'b0_100111110011_101_1_101001111100;
      patterns[20382] = 29'b0_100111110011_110_0_100111110011;
      patterns[20383] = 29'b0_100111110011_111_0_100111110011;
      patterns[20384] = 29'b0_100111110100_000_0_100111110100;
      patterns[20385] = 29'b0_100111110100_001_0_110100100111;
      patterns[20386] = 29'b0_100111110100_010_1_001111101000;
      patterns[20387] = 29'b0_100111110100_011_0_011111010001;
      patterns[20388] = 29'b0_100111110100_100_0_010011111010;
      patterns[20389] = 29'b0_100111110100_101_0_001001111101;
      patterns[20390] = 29'b0_100111110100_110_0_100111110100;
      patterns[20391] = 29'b0_100111110100_111_0_100111110100;
      patterns[20392] = 29'b0_100111110101_000_0_100111110101;
      patterns[20393] = 29'b0_100111110101_001_0_110101100111;
      patterns[20394] = 29'b0_100111110101_010_1_001111101010;
      patterns[20395] = 29'b0_100111110101_011_0_011111010101;
      patterns[20396] = 29'b0_100111110101_100_1_010011111010;
      patterns[20397] = 29'b0_100111110101_101_0_101001111101;
      patterns[20398] = 29'b0_100111110101_110_0_100111110101;
      patterns[20399] = 29'b0_100111110101_111_0_100111110101;
      patterns[20400] = 29'b0_100111110110_000_0_100111110110;
      patterns[20401] = 29'b0_100111110110_001_0_110110100111;
      patterns[20402] = 29'b0_100111110110_010_1_001111101100;
      patterns[20403] = 29'b0_100111110110_011_0_011111011001;
      patterns[20404] = 29'b0_100111110110_100_0_010011111011;
      patterns[20405] = 29'b0_100111110110_101_1_001001111101;
      patterns[20406] = 29'b0_100111110110_110_0_100111110110;
      patterns[20407] = 29'b0_100111110110_111_0_100111110110;
      patterns[20408] = 29'b0_100111110111_000_0_100111110111;
      patterns[20409] = 29'b0_100111110111_001_0_110111100111;
      patterns[20410] = 29'b0_100111110111_010_1_001111101110;
      patterns[20411] = 29'b0_100111110111_011_0_011111011101;
      patterns[20412] = 29'b0_100111110111_100_1_010011111011;
      patterns[20413] = 29'b0_100111110111_101_1_101001111101;
      patterns[20414] = 29'b0_100111110111_110_0_100111110111;
      patterns[20415] = 29'b0_100111110111_111_0_100111110111;
      patterns[20416] = 29'b0_100111111000_000_0_100111111000;
      patterns[20417] = 29'b0_100111111000_001_0_111000100111;
      patterns[20418] = 29'b0_100111111000_010_1_001111110000;
      patterns[20419] = 29'b0_100111111000_011_0_011111100001;
      patterns[20420] = 29'b0_100111111000_100_0_010011111100;
      patterns[20421] = 29'b0_100111111000_101_0_001001111110;
      patterns[20422] = 29'b0_100111111000_110_0_100111111000;
      patterns[20423] = 29'b0_100111111000_111_0_100111111000;
      patterns[20424] = 29'b0_100111111001_000_0_100111111001;
      patterns[20425] = 29'b0_100111111001_001_0_111001100111;
      patterns[20426] = 29'b0_100111111001_010_1_001111110010;
      patterns[20427] = 29'b0_100111111001_011_0_011111100101;
      patterns[20428] = 29'b0_100111111001_100_1_010011111100;
      patterns[20429] = 29'b0_100111111001_101_0_101001111110;
      patterns[20430] = 29'b0_100111111001_110_0_100111111001;
      patterns[20431] = 29'b0_100111111001_111_0_100111111001;
      patterns[20432] = 29'b0_100111111010_000_0_100111111010;
      patterns[20433] = 29'b0_100111111010_001_0_111010100111;
      patterns[20434] = 29'b0_100111111010_010_1_001111110100;
      patterns[20435] = 29'b0_100111111010_011_0_011111101001;
      patterns[20436] = 29'b0_100111111010_100_0_010011111101;
      patterns[20437] = 29'b0_100111111010_101_1_001001111110;
      patterns[20438] = 29'b0_100111111010_110_0_100111111010;
      patterns[20439] = 29'b0_100111111010_111_0_100111111010;
      patterns[20440] = 29'b0_100111111011_000_0_100111111011;
      patterns[20441] = 29'b0_100111111011_001_0_111011100111;
      patterns[20442] = 29'b0_100111111011_010_1_001111110110;
      patterns[20443] = 29'b0_100111111011_011_0_011111101101;
      patterns[20444] = 29'b0_100111111011_100_1_010011111101;
      patterns[20445] = 29'b0_100111111011_101_1_101001111110;
      patterns[20446] = 29'b0_100111111011_110_0_100111111011;
      patterns[20447] = 29'b0_100111111011_111_0_100111111011;
      patterns[20448] = 29'b0_100111111100_000_0_100111111100;
      patterns[20449] = 29'b0_100111111100_001_0_111100100111;
      patterns[20450] = 29'b0_100111111100_010_1_001111111000;
      patterns[20451] = 29'b0_100111111100_011_0_011111110001;
      patterns[20452] = 29'b0_100111111100_100_0_010011111110;
      patterns[20453] = 29'b0_100111111100_101_0_001001111111;
      patterns[20454] = 29'b0_100111111100_110_0_100111111100;
      patterns[20455] = 29'b0_100111111100_111_0_100111111100;
      patterns[20456] = 29'b0_100111111101_000_0_100111111101;
      patterns[20457] = 29'b0_100111111101_001_0_111101100111;
      patterns[20458] = 29'b0_100111111101_010_1_001111111010;
      patterns[20459] = 29'b0_100111111101_011_0_011111110101;
      patterns[20460] = 29'b0_100111111101_100_1_010011111110;
      patterns[20461] = 29'b0_100111111101_101_0_101001111111;
      patterns[20462] = 29'b0_100111111101_110_0_100111111101;
      patterns[20463] = 29'b0_100111111101_111_0_100111111101;
      patterns[20464] = 29'b0_100111111110_000_0_100111111110;
      patterns[20465] = 29'b0_100111111110_001_0_111110100111;
      patterns[20466] = 29'b0_100111111110_010_1_001111111100;
      patterns[20467] = 29'b0_100111111110_011_0_011111111001;
      patterns[20468] = 29'b0_100111111110_100_0_010011111111;
      patterns[20469] = 29'b0_100111111110_101_1_001001111111;
      patterns[20470] = 29'b0_100111111110_110_0_100111111110;
      patterns[20471] = 29'b0_100111111110_111_0_100111111110;
      patterns[20472] = 29'b0_100111111111_000_0_100111111111;
      patterns[20473] = 29'b0_100111111111_001_0_111111100111;
      patterns[20474] = 29'b0_100111111111_010_1_001111111110;
      patterns[20475] = 29'b0_100111111111_011_0_011111111101;
      patterns[20476] = 29'b0_100111111111_100_1_010011111111;
      patterns[20477] = 29'b0_100111111111_101_1_101001111111;
      patterns[20478] = 29'b0_100111111111_110_0_100111111111;
      patterns[20479] = 29'b0_100111111111_111_0_100111111111;
      patterns[20480] = 29'b0_101000000000_000_0_101000000000;
      patterns[20481] = 29'b0_101000000000_001_0_000000101000;
      patterns[20482] = 29'b0_101000000000_010_1_010000000000;
      patterns[20483] = 29'b0_101000000000_011_0_100000000001;
      patterns[20484] = 29'b0_101000000000_100_0_010100000000;
      patterns[20485] = 29'b0_101000000000_101_0_001010000000;
      patterns[20486] = 29'b0_101000000000_110_0_101000000000;
      patterns[20487] = 29'b0_101000000000_111_0_101000000000;
      patterns[20488] = 29'b0_101000000001_000_0_101000000001;
      patterns[20489] = 29'b0_101000000001_001_0_000001101000;
      patterns[20490] = 29'b0_101000000001_010_1_010000000010;
      patterns[20491] = 29'b0_101000000001_011_0_100000000101;
      patterns[20492] = 29'b0_101000000001_100_1_010100000000;
      patterns[20493] = 29'b0_101000000001_101_0_101010000000;
      patterns[20494] = 29'b0_101000000001_110_0_101000000001;
      patterns[20495] = 29'b0_101000000001_111_0_101000000001;
      patterns[20496] = 29'b0_101000000010_000_0_101000000010;
      patterns[20497] = 29'b0_101000000010_001_0_000010101000;
      patterns[20498] = 29'b0_101000000010_010_1_010000000100;
      patterns[20499] = 29'b0_101000000010_011_0_100000001001;
      patterns[20500] = 29'b0_101000000010_100_0_010100000001;
      patterns[20501] = 29'b0_101000000010_101_1_001010000000;
      patterns[20502] = 29'b0_101000000010_110_0_101000000010;
      patterns[20503] = 29'b0_101000000010_111_0_101000000010;
      patterns[20504] = 29'b0_101000000011_000_0_101000000011;
      patterns[20505] = 29'b0_101000000011_001_0_000011101000;
      patterns[20506] = 29'b0_101000000011_010_1_010000000110;
      patterns[20507] = 29'b0_101000000011_011_0_100000001101;
      patterns[20508] = 29'b0_101000000011_100_1_010100000001;
      patterns[20509] = 29'b0_101000000011_101_1_101010000000;
      patterns[20510] = 29'b0_101000000011_110_0_101000000011;
      patterns[20511] = 29'b0_101000000011_111_0_101000000011;
      patterns[20512] = 29'b0_101000000100_000_0_101000000100;
      patterns[20513] = 29'b0_101000000100_001_0_000100101000;
      patterns[20514] = 29'b0_101000000100_010_1_010000001000;
      patterns[20515] = 29'b0_101000000100_011_0_100000010001;
      patterns[20516] = 29'b0_101000000100_100_0_010100000010;
      patterns[20517] = 29'b0_101000000100_101_0_001010000001;
      patterns[20518] = 29'b0_101000000100_110_0_101000000100;
      patterns[20519] = 29'b0_101000000100_111_0_101000000100;
      patterns[20520] = 29'b0_101000000101_000_0_101000000101;
      patterns[20521] = 29'b0_101000000101_001_0_000101101000;
      patterns[20522] = 29'b0_101000000101_010_1_010000001010;
      patterns[20523] = 29'b0_101000000101_011_0_100000010101;
      patterns[20524] = 29'b0_101000000101_100_1_010100000010;
      patterns[20525] = 29'b0_101000000101_101_0_101010000001;
      patterns[20526] = 29'b0_101000000101_110_0_101000000101;
      patterns[20527] = 29'b0_101000000101_111_0_101000000101;
      patterns[20528] = 29'b0_101000000110_000_0_101000000110;
      patterns[20529] = 29'b0_101000000110_001_0_000110101000;
      patterns[20530] = 29'b0_101000000110_010_1_010000001100;
      patterns[20531] = 29'b0_101000000110_011_0_100000011001;
      patterns[20532] = 29'b0_101000000110_100_0_010100000011;
      patterns[20533] = 29'b0_101000000110_101_1_001010000001;
      patterns[20534] = 29'b0_101000000110_110_0_101000000110;
      patterns[20535] = 29'b0_101000000110_111_0_101000000110;
      patterns[20536] = 29'b0_101000000111_000_0_101000000111;
      patterns[20537] = 29'b0_101000000111_001_0_000111101000;
      patterns[20538] = 29'b0_101000000111_010_1_010000001110;
      patterns[20539] = 29'b0_101000000111_011_0_100000011101;
      patterns[20540] = 29'b0_101000000111_100_1_010100000011;
      patterns[20541] = 29'b0_101000000111_101_1_101010000001;
      patterns[20542] = 29'b0_101000000111_110_0_101000000111;
      patterns[20543] = 29'b0_101000000111_111_0_101000000111;
      patterns[20544] = 29'b0_101000001000_000_0_101000001000;
      patterns[20545] = 29'b0_101000001000_001_0_001000101000;
      patterns[20546] = 29'b0_101000001000_010_1_010000010000;
      patterns[20547] = 29'b0_101000001000_011_0_100000100001;
      patterns[20548] = 29'b0_101000001000_100_0_010100000100;
      patterns[20549] = 29'b0_101000001000_101_0_001010000010;
      patterns[20550] = 29'b0_101000001000_110_0_101000001000;
      patterns[20551] = 29'b0_101000001000_111_0_101000001000;
      patterns[20552] = 29'b0_101000001001_000_0_101000001001;
      patterns[20553] = 29'b0_101000001001_001_0_001001101000;
      patterns[20554] = 29'b0_101000001001_010_1_010000010010;
      patterns[20555] = 29'b0_101000001001_011_0_100000100101;
      patterns[20556] = 29'b0_101000001001_100_1_010100000100;
      patterns[20557] = 29'b0_101000001001_101_0_101010000010;
      patterns[20558] = 29'b0_101000001001_110_0_101000001001;
      patterns[20559] = 29'b0_101000001001_111_0_101000001001;
      patterns[20560] = 29'b0_101000001010_000_0_101000001010;
      patterns[20561] = 29'b0_101000001010_001_0_001010101000;
      patterns[20562] = 29'b0_101000001010_010_1_010000010100;
      patterns[20563] = 29'b0_101000001010_011_0_100000101001;
      patterns[20564] = 29'b0_101000001010_100_0_010100000101;
      patterns[20565] = 29'b0_101000001010_101_1_001010000010;
      patterns[20566] = 29'b0_101000001010_110_0_101000001010;
      patterns[20567] = 29'b0_101000001010_111_0_101000001010;
      patterns[20568] = 29'b0_101000001011_000_0_101000001011;
      patterns[20569] = 29'b0_101000001011_001_0_001011101000;
      patterns[20570] = 29'b0_101000001011_010_1_010000010110;
      patterns[20571] = 29'b0_101000001011_011_0_100000101101;
      patterns[20572] = 29'b0_101000001011_100_1_010100000101;
      patterns[20573] = 29'b0_101000001011_101_1_101010000010;
      patterns[20574] = 29'b0_101000001011_110_0_101000001011;
      patterns[20575] = 29'b0_101000001011_111_0_101000001011;
      patterns[20576] = 29'b0_101000001100_000_0_101000001100;
      patterns[20577] = 29'b0_101000001100_001_0_001100101000;
      patterns[20578] = 29'b0_101000001100_010_1_010000011000;
      patterns[20579] = 29'b0_101000001100_011_0_100000110001;
      patterns[20580] = 29'b0_101000001100_100_0_010100000110;
      patterns[20581] = 29'b0_101000001100_101_0_001010000011;
      patterns[20582] = 29'b0_101000001100_110_0_101000001100;
      patterns[20583] = 29'b0_101000001100_111_0_101000001100;
      patterns[20584] = 29'b0_101000001101_000_0_101000001101;
      patterns[20585] = 29'b0_101000001101_001_0_001101101000;
      patterns[20586] = 29'b0_101000001101_010_1_010000011010;
      patterns[20587] = 29'b0_101000001101_011_0_100000110101;
      patterns[20588] = 29'b0_101000001101_100_1_010100000110;
      patterns[20589] = 29'b0_101000001101_101_0_101010000011;
      patterns[20590] = 29'b0_101000001101_110_0_101000001101;
      patterns[20591] = 29'b0_101000001101_111_0_101000001101;
      patterns[20592] = 29'b0_101000001110_000_0_101000001110;
      patterns[20593] = 29'b0_101000001110_001_0_001110101000;
      patterns[20594] = 29'b0_101000001110_010_1_010000011100;
      patterns[20595] = 29'b0_101000001110_011_0_100000111001;
      patterns[20596] = 29'b0_101000001110_100_0_010100000111;
      patterns[20597] = 29'b0_101000001110_101_1_001010000011;
      patterns[20598] = 29'b0_101000001110_110_0_101000001110;
      patterns[20599] = 29'b0_101000001110_111_0_101000001110;
      patterns[20600] = 29'b0_101000001111_000_0_101000001111;
      patterns[20601] = 29'b0_101000001111_001_0_001111101000;
      patterns[20602] = 29'b0_101000001111_010_1_010000011110;
      patterns[20603] = 29'b0_101000001111_011_0_100000111101;
      patterns[20604] = 29'b0_101000001111_100_1_010100000111;
      patterns[20605] = 29'b0_101000001111_101_1_101010000011;
      patterns[20606] = 29'b0_101000001111_110_0_101000001111;
      patterns[20607] = 29'b0_101000001111_111_0_101000001111;
      patterns[20608] = 29'b0_101000010000_000_0_101000010000;
      patterns[20609] = 29'b0_101000010000_001_0_010000101000;
      patterns[20610] = 29'b0_101000010000_010_1_010000100000;
      patterns[20611] = 29'b0_101000010000_011_0_100001000001;
      patterns[20612] = 29'b0_101000010000_100_0_010100001000;
      patterns[20613] = 29'b0_101000010000_101_0_001010000100;
      patterns[20614] = 29'b0_101000010000_110_0_101000010000;
      patterns[20615] = 29'b0_101000010000_111_0_101000010000;
      patterns[20616] = 29'b0_101000010001_000_0_101000010001;
      patterns[20617] = 29'b0_101000010001_001_0_010001101000;
      patterns[20618] = 29'b0_101000010001_010_1_010000100010;
      patterns[20619] = 29'b0_101000010001_011_0_100001000101;
      patterns[20620] = 29'b0_101000010001_100_1_010100001000;
      patterns[20621] = 29'b0_101000010001_101_0_101010000100;
      patterns[20622] = 29'b0_101000010001_110_0_101000010001;
      patterns[20623] = 29'b0_101000010001_111_0_101000010001;
      patterns[20624] = 29'b0_101000010010_000_0_101000010010;
      patterns[20625] = 29'b0_101000010010_001_0_010010101000;
      patterns[20626] = 29'b0_101000010010_010_1_010000100100;
      patterns[20627] = 29'b0_101000010010_011_0_100001001001;
      patterns[20628] = 29'b0_101000010010_100_0_010100001001;
      patterns[20629] = 29'b0_101000010010_101_1_001010000100;
      patterns[20630] = 29'b0_101000010010_110_0_101000010010;
      patterns[20631] = 29'b0_101000010010_111_0_101000010010;
      patterns[20632] = 29'b0_101000010011_000_0_101000010011;
      patterns[20633] = 29'b0_101000010011_001_0_010011101000;
      patterns[20634] = 29'b0_101000010011_010_1_010000100110;
      patterns[20635] = 29'b0_101000010011_011_0_100001001101;
      patterns[20636] = 29'b0_101000010011_100_1_010100001001;
      patterns[20637] = 29'b0_101000010011_101_1_101010000100;
      patterns[20638] = 29'b0_101000010011_110_0_101000010011;
      patterns[20639] = 29'b0_101000010011_111_0_101000010011;
      patterns[20640] = 29'b0_101000010100_000_0_101000010100;
      patterns[20641] = 29'b0_101000010100_001_0_010100101000;
      patterns[20642] = 29'b0_101000010100_010_1_010000101000;
      patterns[20643] = 29'b0_101000010100_011_0_100001010001;
      patterns[20644] = 29'b0_101000010100_100_0_010100001010;
      patterns[20645] = 29'b0_101000010100_101_0_001010000101;
      patterns[20646] = 29'b0_101000010100_110_0_101000010100;
      patterns[20647] = 29'b0_101000010100_111_0_101000010100;
      patterns[20648] = 29'b0_101000010101_000_0_101000010101;
      patterns[20649] = 29'b0_101000010101_001_0_010101101000;
      patterns[20650] = 29'b0_101000010101_010_1_010000101010;
      patterns[20651] = 29'b0_101000010101_011_0_100001010101;
      patterns[20652] = 29'b0_101000010101_100_1_010100001010;
      patterns[20653] = 29'b0_101000010101_101_0_101010000101;
      patterns[20654] = 29'b0_101000010101_110_0_101000010101;
      patterns[20655] = 29'b0_101000010101_111_0_101000010101;
      patterns[20656] = 29'b0_101000010110_000_0_101000010110;
      patterns[20657] = 29'b0_101000010110_001_0_010110101000;
      patterns[20658] = 29'b0_101000010110_010_1_010000101100;
      patterns[20659] = 29'b0_101000010110_011_0_100001011001;
      patterns[20660] = 29'b0_101000010110_100_0_010100001011;
      patterns[20661] = 29'b0_101000010110_101_1_001010000101;
      patterns[20662] = 29'b0_101000010110_110_0_101000010110;
      patterns[20663] = 29'b0_101000010110_111_0_101000010110;
      patterns[20664] = 29'b0_101000010111_000_0_101000010111;
      patterns[20665] = 29'b0_101000010111_001_0_010111101000;
      patterns[20666] = 29'b0_101000010111_010_1_010000101110;
      patterns[20667] = 29'b0_101000010111_011_0_100001011101;
      patterns[20668] = 29'b0_101000010111_100_1_010100001011;
      patterns[20669] = 29'b0_101000010111_101_1_101010000101;
      patterns[20670] = 29'b0_101000010111_110_0_101000010111;
      patterns[20671] = 29'b0_101000010111_111_0_101000010111;
      patterns[20672] = 29'b0_101000011000_000_0_101000011000;
      patterns[20673] = 29'b0_101000011000_001_0_011000101000;
      patterns[20674] = 29'b0_101000011000_010_1_010000110000;
      patterns[20675] = 29'b0_101000011000_011_0_100001100001;
      patterns[20676] = 29'b0_101000011000_100_0_010100001100;
      patterns[20677] = 29'b0_101000011000_101_0_001010000110;
      patterns[20678] = 29'b0_101000011000_110_0_101000011000;
      patterns[20679] = 29'b0_101000011000_111_0_101000011000;
      patterns[20680] = 29'b0_101000011001_000_0_101000011001;
      patterns[20681] = 29'b0_101000011001_001_0_011001101000;
      patterns[20682] = 29'b0_101000011001_010_1_010000110010;
      patterns[20683] = 29'b0_101000011001_011_0_100001100101;
      patterns[20684] = 29'b0_101000011001_100_1_010100001100;
      patterns[20685] = 29'b0_101000011001_101_0_101010000110;
      patterns[20686] = 29'b0_101000011001_110_0_101000011001;
      patterns[20687] = 29'b0_101000011001_111_0_101000011001;
      patterns[20688] = 29'b0_101000011010_000_0_101000011010;
      patterns[20689] = 29'b0_101000011010_001_0_011010101000;
      patterns[20690] = 29'b0_101000011010_010_1_010000110100;
      patterns[20691] = 29'b0_101000011010_011_0_100001101001;
      patterns[20692] = 29'b0_101000011010_100_0_010100001101;
      patterns[20693] = 29'b0_101000011010_101_1_001010000110;
      patterns[20694] = 29'b0_101000011010_110_0_101000011010;
      patterns[20695] = 29'b0_101000011010_111_0_101000011010;
      patterns[20696] = 29'b0_101000011011_000_0_101000011011;
      patterns[20697] = 29'b0_101000011011_001_0_011011101000;
      patterns[20698] = 29'b0_101000011011_010_1_010000110110;
      patterns[20699] = 29'b0_101000011011_011_0_100001101101;
      patterns[20700] = 29'b0_101000011011_100_1_010100001101;
      patterns[20701] = 29'b0_101000011011_101_1_101010000110;
      patterns[20702] = 29'b0_101000011011_110_0_101000011011;
      patterns[20703] = 29'b0_101000011011_111_0_101000011011;
      patterns[20704] = 29'b0_101000011100_000_0_101000011100;
      patterns[20705] = 29'b0_101000011100_001_0_011100101000;
      patterns[20706] = 29'b0_101000011100_010_1_010000111000;
      patterns[20707] = 29'b0_101000011100_011_0_100001110001;
      patterns[20708] = 29'b0_101000011100_100_0_010100001110;
      patterns[20709] = 29'b0_101000011100_101_0_001010000111;
      patterns[20710] = 29'b0_101000011100_110_0_101000011100;
      patterns[20711] = 29'b0_101000011100_111_0_101000011100;
      patterns[20712] = 29'b0_101000011101_000_0_101000011101;
      patterns[20713] = 29'b0_101000011101_001_0_011101101000;
      patterns[20714] = 29'b0_101000011101_010_1_010000111010;
      patterns[20715] = 29'b0_101000011101_011_0_100001110101;
      patterns[20716] = 29'b0_101000011101_100_1_010100001110;
      patterns[20717] = 29'b0_101000011101_101_0_101010000111;
      patterns[20718] = 29'b0_101000011101_110_0_101000011101;
      patterns[20719] = 29'b0_101000011101_111_0_101000011101;
      patterns[20720] = 29'b0_101000011110_000_0_101000011110;
      patterns[20721] = 29'b0_101000011110_001_0_011110101000;
      patterns[20722] = 29'b0_101000011110_010_1_010000111100;
      patterns[20723] = 29'b0_101000011110_011_0_100001111001;
      patterns[20724] = 29'b0_101000011110_100_0_010100001111;
      patterns[20725] = 29'b0_101000011110_101_1_001010000111;
      patterns[20726] = 29'b0_101000011110_110_0_101000011110;
      patterns[20727] = 29'b0_101000011110_111_0_101000011110;
      patterns[20728] = 29'b0_101000011111_000_0_101000011111;
      patterns[20729] = 29'b0_101000011111_001_0_011111101000;
      patterns[20730] = 29'b0_101000011111_010_1_010000111110;
      patterns[20731] = 29'b0_101000011111_011_0_100001111101;
      patterns[20732] = 29'b0_101000011111_100_1_010100001111;
      patterns[20733] = 29'b0_101000011111_101_1_101010000111;
      patterns[20734] = 29'b0_101000011111_110_0_101000011111;
      patterns[20735] = 29'b0_101000011111_111_0_101000011111;
      patterns[20736] = 29'b0_101000100000_000_0_101000100000;
      patterns[20737] = 29'b0_101000100000_001_0_100000101000;
      patterns[20738] = 29'b0_101000100000_010_1_010001000000;
      patterns[20739] = 29'b0_101000100000_011_0_100010000001;
      patterns[20740] = 29'b0_101000100000_100_0_010100010000;
      patterns[20741] = 29'b0_101000100000_101_0_001010001000;
      patterns[20742] = 29'b0_101000100000_110_0_101000100000;
      patterns[20743] = 29'b0_101000100000_111_0_101000100000;
      patterns[20744] = 29'b0_101000100001_000_0_101000100001;
      patterns[20745] = 29'b0_101000100001_001_0_100001101000;
      patterns[20746] = 29'b0_101000100001_010_1_010001000010;
      patterns[20747] = 29'b0_101000100001_011_0_100010000101;
      patterns[20748] = 29'b0_101000100001_100_1_010100010000;
      patterns[20749] = 29'b0_101000100001_101_0_101010001000;
      patterns[20750] = 29'b0_101000100001_110_0_101000100001;
      patterns[20751] = 29'b0_101000100001_111_0_101000100001;
      patterns[20752] = 29'b0_101000100010_000_0_101000100010;
      patterns[20753] = 29'b0_101000100010_001_0_100010101000;
      patterns[20754] = 29'b0_101000100010_010_1_010001000100;
      patterns[20755] = 29'b0_101000100010_011_0_100010001001;
      patterns[20756] = 29'b0_101000100010_100_0_010100010001;
      patterns[20757] = 29'b0_101000100010_101_1_001010001000;
      patterns[20758] = 29'b0_101000100010_110_0_101000100010;
      patterns[20759] = 29'b0_101000100010_111_0_101000100010;
      patterns[20760] = 29'b0_101000100011_000_0_101000100011;
      patterns[20761] = 29'b0_101000100011_001_0_100011101000;
      patterns[20762] = 29'b0_101000100011_010_1_010001000110;
      patterns[20763] = 29'b0_101000100011_011_0_100010001101;
      patterns[20764] = 29'b0_101000100011_100_1_010100010001;
      patterns[20765] = 29'b0_101000100011_101_1_101010001000;
      patterns[20766] = 29'b0_101000100011_110_0_101000100011;
      patterns[20767] = 29'b0_101000100011_111_0_101000100011;
      patterns[20768] = 29'b0_101000100100_000_0_101000100100;
      patterns[20769] = 29'b0_101000100100_001_0_100100101000;
      patterns[20770] = 29'b0_101000100100_010_1_010001001000;
      patterns[20771] = 29'b0_101000100100_011_0_100010010001;
      patterns[20772] = 29'b0_101000100100_100_0_010100010010;
      patterns[20773] = 29'b0_101000100100_101_0_001010001001;
      patterns[20774] = 29'b0_101000100100_110_0_101000100100;
      patterns[20775] = 29'b0_101000100100_111_0_101000100100;
      patterns[20776] = 29'b0_101000100101_000_0_101000100101;
      patterns[20777] = 29'b0_101000100101_001_0_100101101000;
      patterns[20778] = 29'b0_101000100101_010_1_010001001010;
      patterns[20779] = 29'b0_101000100101_011_0_100010010101;
      patterns[20780] = 29'b0_101000100101_100_1_010100010010;
      patterns[20781] = 29'b0_101000100101_101_0_101010001001;
      patterns[20782] = 29'b0_101000100101_110_0_101000100101;
      patterns[20783] = 29'b0_101000100101_111_0_101000100101;
      patterns[20784] = 29'b0_101000100110_000_0_101000100110;
      patterns[20785] = 29'b0_101000100110_001_0_100110101000;
      patterns[20786] = 29'b0_101000100110_010_1_010001001100;
      patterns[20787] = 29'b0_101000100110_011_0_100010011001;
      patterns[20788] = 29'b0_101000100110_100_0_010100010011;
      patterns[20789] = 29'b0_101000100110_101_1_001010001001;
      patterns[20790] = 29'b0_101000100110_110_0_101000100110;
      patterns[20791] = 29'b0_101000100110_111_0_101000100110;
      patterns[20792] = 29'b0_101000100111_000_0_101000100111;
      patterns[20793] = 29'b0_101000100111_001_0_100111101000;
      patterns[20794] = 29'b0_101000100111_010_1_010001001110;
      patterns[20795] = 29'b0_101000100111_011_0_100010011101;
      patterns[20796] = 29'b0_101000100111_100_1_010100010011;
      patterns[20797] = 29'b0_101000100111_101_1_101010001001;
      patterns[20798] = 29'b0_101000100111_110_0_101000100111;
      patterns[20799] = 29'b0_101000100111_111_0_101000100111;
      patterns[20800] = 29'b0_101000101000_000_0_101000101000;
      patterns[20801] = 29'b0_101000101000_001_0_101000101000;
      patterns[20802] = 29'b0_101000101000_010_1_010001010000;
      patterns[20803] = 29'b0_101000101000_011_0_100010100001;
      patterns[20804] = 29'b0_101000101000_100_0_010100010100;
      patterns[20805] = 29'b0_101000101000_101_0_001010001010;
      patterns[20806] = 29'b0_101000101000_110_0_101000101000;
      patterns[20807] = 29'b0_101000101000_111_0_101000101000;
      patterns[20808] = 29'b0_101000101001_000_0_101000101001;
      patterns[20809] = 29'b0_101000101001_001_0_101001101000;
      patterns[20810] = 29'b0_101000101001_010_1_010001010010;
      patterns[20811] = 29'b0_101000101001_011_0_100010100101;
      patterns[20812] = 29'b0_101000101001_100_1_010100010100;
      patterns[20813] = 29'b0_101000101001_101_0_101010001010;
      patterns[20814] = 29'b0_101000101001_110_0_101000101001;
      patterns[20815] = 29'b0_101000101001_111_0_101000101001;
      patterns[20816] = 29'b0_101000101010_000_0_101000101010;
      patterns[20817] = 29'b0_101000101010_001_0_101010101000;
      patterns[20818] = 29'b0_101000101010_010_1_010001010100;
      patterns[20819] = 29'b0_101000101010_011_0_100010101001;
      patterns[20820] = 29'b0_101000101010_100_0_010100010101;
      patterns[20821] = 29'b0_101000101010_101_1_001010001010;
      patterns[20822] = 29'b0_101000101010_110_0_101000101010;
      patterns[20823] = 29'b0_101000101010_111_0_101000101010;
      patterns[20824] = 29'b0_101000101011_000_0_101000101011;
      patterns[20825] = 29'b0_101000101011_001_0_101011101000;
      patterns[20826] = 29'b0_101000101011_010_1_010001010110;
      patterns[20827] = 29'b0_101000101011_011_0_100010101101;
      patterns[20828] = 29'b0_101000101011_100_1_010100010101;
      patterns[20829] = 29'b0_101000101011_101_1_101010001010;
      patterns[20830] = 29'b0_101000101011_110_0_101000101011;
      patterns[20831] = 29'b0_101000101011_111_0_101000101011;
      patterns[20832] = 29'b0_101000101100_000_0_101000101100;
      patterns[20833] = 29'b0_101000101100_001_0_101100101000;
      patterns[20834] = 29'b0_101000101100_010_1_010001011000;
      patterns[20835] = 29'b0_101000101100_011_0_100010110001;
      patterns[20836] = 29'b0_101000101100_100_0_010100010110;
      patterns[20837] = 29'b0_101000101100_101_0_001010001011;
      patterns[20838] = 29'b0_101000101100_110_0_101000101100;
      patterns[20839] = 29'b0_101000101100_111_0_101000101100;
      patterns[20840] = 29'b0_101000101101_000_0_101000101101;
      patterns[20841] = 29'b0_101000101101_001_0_101101101000;
      patterns[20842] = 29'b0_101000101101_010_1_010001011010;
      patterns[20843] = 29'b0_101000101101_011_0_100010110101;
      patterns[20844] = 29'b0_101000101101_100_1_010100010110;
      patterns[20845] = 29'b0_101000101101_101_0_101010001011;
      patterns[20846] = 29'b0_101000101101_110_0_101000101101;
      patterns[20847] = 29'b0_101000101101_111_0_101000101101;
      patterns[20848] = 29'b0_101000101110_000_0_101000101110;
      patterns[20849] = 29'b0_101000101110_001_0_101110101000;
      patterns[20850] = 29'b0_101000101110_010_1_010001011100;
      patterns[20851] = 29'b0_101000101110_011_0_100010111001;
      patterns[20852] = 29'b0_101000101110_100_0_010100010111;
      patterns[20853] = 29'b0_101000101110_101_1_001010001011;
      patterns[20854] = 29'b0_101000101110_110_0_101000101110;
      patterns[20855] = 29'b0_101000101110_111_0_101000101110;
      patterns[20856] = 29'b0_101000101111_000_0_101000101111;
      patterns[20857] = 29'b0_101000101111_001_0_101111101000;
      patterns[20858] = 29'b0_101000101111_010_1_010001011110;
      patterns[20859] = 29'b0_101000101111_011_0_100010111101;
      patterns[20860] = 29'b0_101000101111_100_1_010100010111;
      patterns[20861] = 29'b0_101000101111_101_1_101010001011;
      patterns[20862] = 29'b0_101000101111_110_0_101000101111;
      patterns[20863] = 29'b0_101000101111_111_0_101000101111;
      patterns[20864] = 29'b0_101000110000_000_0_101000110000;
      patterns[20865] = 29'b0_101000110000_001_0_110000101000;
      patterns[20866] = 29'b0_101000110000_010_1_010001100000;
      patterns[20867] = 29'b0_101000110000_011_0_100011000001;
      patterns[20868] = 29'b0_101000110000_100_0_010100011000;
      patterns[20869] = 29'b0_101000110000_101_0_001010001100;
      patterns[20870] = 29'b0_101000110000_110_0_101000110000;
      patterns[20871] = 29'b0_101000110000_111_0_101000110000;
      patterns[20872] = 29'b0_101000110001_000_0_101000110001;
      patterns[20873] = 29'b0_101000110001_001_0_110001101000;
      patterns[20874] = 29'b0_101000110001_010_1_010001100010;
      patterns[20875] = 29'b0_101000110001_011_0_100011000101;
      patterns[20876] = 29'b0_101000110001_100_1_010100011000;
      patterns[20877] = 29'b0_101000110001_101_0_101010001100;
      patterns[20878] = 29'b0_101000110001_110_0_101000110001;
      patterns[20879] = 29'b0_101000110001_111_0_101000110001;
      patterns[20880] = 29'b0_101000110010_000_0_101000110010;
      patterns[20881] = 29'b0_101000110010_001_0_110010101000;
      patterns[20882] = 29'b0_101000110010_010_1_010001100100;
      patterns[20883] = 29'b0_101000110010_011_0_100011001001;
      patterns[20884] = 29'b0_101000110010_100_0_010100011001;
      patterns[20885] = 29'b0_101000110010_101_1_001010001100;
      patterns[20886] = 29'b0_101000110010_110_0_101000110010;
      patterns[20887] = 29'b0_101000110010_111_0_101000110010;
      patterns[20888] = 29'b0_101000110011_000_0_101000110011;
      patterns[20889] = 29'b0_101000110011_001_0_110011101000;
      patterns[20890] = 29'b0_101000110011_010_1_010001100110;
      patterns[20891] = 29'b0_101000110011_011_0_100011001101;
      patterns[20892] = 29'b0_101000110011_100_1_010100011001;
      patterns[20893] = 29'b0_101000110011_101_1_101010001100;
      patterns[20894] = 29'b0_101000110011_110_0_101000110011;
      patterns[20895] = 29'b0_101000110011_111_0_101000110011;
      patterns[20896] = 29'b0_101000110100_000_0_101000110100;
      patterns[20897] = 29'b0_101000110100_001_0_110100101000;
      patterns[20898] = 29'b0_101000110100_010_1_010001101000;
      patterns[20899] = 29'b0_101000110100_011_0_100011010001;
      patterns[20900] = 29'b0_101000110100_100_0_010100011010;
      patterns[20901] = 29'b0_101000110100_101_0_001010001101;
      patterns[20902] = 29'b0_101000110100_110_0_101000110100;
      patterns[20903] = 29'b0_101000110100_111_0_101000110100;
      patterns[20904] = 29'b0_101000110101_000_0_101000110101;
      patterns[20905] = 29'b0_101000110101_001_0_110101101000;
      patterns[20906] = 29'b0_101000110101_010_1_010001101010;
      patterns[20907] = 29'b0_101000110101_011_0_100011010101;
      patterns[20908] = 29'b0_101000110101_100_1_010100011010;
      patterns[20909] = 29'b0_101000110101_101_0_101010001101;
      patterns[20910] = 29'b0_101000110101_110_0_101000110101;
      patterns[20911] = 29'b0_101000110101_111_0_101000110101;
      patterns[20912] = 29'b0_101000110110_000_0_101000110110;
      patterns[20913] = 29'b0_101000110110_001_0_110110101000;
      patterns[20914] = 29'b0_101000110110_010_1_010001101100;
      patterns[20915] = 29'b0_101000110110_011_0_100011011001;
      patterns[20916] = 29'b0_101000110110_100_0_010100011011;
      patterns[20917] = 29'b0_101000110110_101_1_001010001101;
      patterns[20918] = 29'b0_101000110110_110_0_101000110110;
      patterns[20919] = 29'b0_101000110110_111_0_101000110110;
      patterns[20920] = 29'b0_101000110111_000_0_101000110111;
      patterns[20921] = 29'b0_101000110111_001_0_110111101000;
      patterns[20922] = 29'b0_101000110111_010_1_010001101110;
      patterns[20923] = 29'b0_101000110111_011_0_100011011101;
      patterns[20924] = 29'b0_101000110111_100_1_010100011011;
      patterns[20925] = 29'b0_101000110111_101_1_101010001101;
      patterns[20926] = 29'b0_101000110111_110_0_101000110111;
      patterns[20927] = 29'b0_101000110111_111_0_101000110111;
      patterns[20928] = 29'b0_101000111000_000_0_101000111000;
      patterns[20929] = 29'b0_101000111000_001_0_111000101000;
      patterns[20930] = 29'b0_101000111000_010_1_010001110000;
      patterns[20931] = 29'b0_101000111000_011_0_100011100001;
      patterns[20932] = 29'b0_101000111000_100_0_010100011100;
      patterns[20933] = 29'b0_101000111000_101_0_001010001110;
      patterns[20934] = 29'b0_101000111000_110_0_101000111000;
      patterns[20935] = 29'b0_101000111000_111_0_101000111000;
      patterns[20936] = 29'b0_101000111001_000_0_101000111001;
      patterns[20937] = 29'b0_101000111001_001_0_111001101000;
      patterns[20938] = 29'b0_101000111001_010_1_010001110010;
      patterns[20939] = 29'b0_101000111001_011_0_100011100101;
      patterns[20940] = 29'b0_101000111001_100_1_010100011100;
      patterns[20941] = 29'b0_101000111001_101_0_101010001110;
      patterns[20942] = 29'b0_101000111001_110_0_101000111001;
      patterns[20943] = 29'b0_101000111001_111_0_101000111001;
      patterns[20944] = 29'b0_101000111010_000_0_101000111010;
      patterns[20945] = 29'b0_101000111010_001_0_111010101000;
      patterns[20946] = 29'b0_101000111010_010_1_010001110100;
      patterns[20947] = 29'b0_101000111010_011_0_100011101001;
      patterns[20948] = 29'b0_101000111010_100_0_010100011101;
      patterns[20949] = 29'b0_101000111010_101_1_001010001110;
      patterns[20950] = 29'b0_101000111010_110_0_101000111010;
      patterns[20951] = 29'b0_101000111010_111_0_101000111010;
      patterns[20952] = 29'b0_101000111011_000_0_101000111011;
      patterns[20953] = 29'b0_101000111011_001_0_111011101000;
      patterns[20954] = 29'b0_101000111011_010_1_010001110110;
      patterns[20955] = 29'b0_101000111011_011_0_100011101101;
      patterns[20956] = 29'b0_101000111011_100_1_010100011101;
      patterns[20957] = 29'b0_101000111011_101_1_101010001110;
      patterns[20958] = 29'b0_101000111011_110_0_101000111011;
      patterns[20959] = 29'b0_101000111011_111_0_101000111011;
      patterns[20960] = 29'b0_101000111100_000_0_101000111100;
      patterns[20961] = 29'b0_101000111100_001_0_111100101000;
      patterns[20962] = 29'b0_101000111100_010_1_010001111000;
      patterns[20963] = 29'b0_101000111100_011_0_100011110001;
      patterns[20964] = 29'b0_101000111100_100_0_010100011110;
      patterns[20965] = 29'b0_101000111100_101_0_001010001111;
      patterns[20966] = 29'b0_101000111100_110_0_101000111100;
      patterns[20967] = 29'b0_101000111100_111_0_101000111100;
      patterns[20968] = 29'b0_101000111101_000_0_101000111101;
      patterns[20969] = 29'b0_101000111101_001_0_111101101000;
      patterns[20970] = 29'b0_101000111101_010_1_010001111010;
      patterns[20971] = 29'b0_101000111101_011_0_100011110101;
      patterns[20972] = 29'b0_101000111101_100_1_010100011110;
      patterns[20973] = 29'b0_101000111101_101_0_101010001111;
      patterns[20974] = 29'b0_101000111101_110_0_101000111101;
      patterns[20975] = 29'b0_101000111101_111_0_101000111101;
      patterns[20976] = 29'b0_101000111110_000_0_101000111110;
      patterns[20977] = 29'b0_101000111110_001_0_111110101000;
      patterns[20978] = 29'b0_101000111110_010_1_010001111100;
      patterns[20979] = 29'b0_101000111110_011_0_100011111001;
      patterns[20980] = 29'b0_101000111110_100_0_010100011111;
      patterns[20981] = 29'b0_101000111110_101_1_001010001111;
      patterns[20982] = 29'b0_101000111110_110_0_101000111110;
      patterns[20983] = 29'b0_101000111110_111_0_101000111110;
      patterns[20984] = 29'b0_101000111111_000_0_101000111111;
      patterns[20985] = 29'b0_101000111111_001_0_111111101000;
      patterns[20986] = 29'b0_101000111111_010_1_010001111110;
      patterns[20987] = 29'b0_101000111111_011_0_100011111101;
      patterns[20988] = 29'b0_101000111111_100_1_010100011111;
      patterns[20989] = 29'b0_101000111111_101_1_101010001111;
      patterns[20990] = 29'b0_101000111111_110_0_101000111111;
      patterns[20991] = 29'b0_101000111111_111_0_101000111111;
      patterns[20992] = 29'b0_101001000000_000_0_101001000000;
      patterns[20993] = 29'b0_101001000000_001_0_000000101001;
      patterns[20994] = 29'b0_101001000000_010_1_010010000000;
      patterns[20995] = 29'b0_101001000000_011_0_100100000001;
      patterns[20996] = 29'b0_101001000000_100_0_010100100000;
      patterns[20997] = 29'b0_101001000000_101_0_001010010000;
      patterns[20998] = 29'b0_101001000000_110_0_101001000000;
      patterns[20999] = 29'b0_101001000000_111_0_101001000000;
      patterns[21000] = 29'b0_101001000001_000_0_101001000001;
      patterns[21001] = 29'b0_101001000001_001_0_000001101001;
      patterns[21002] = 29'b0_101001000001_010_1_010010000010;
      patterns[21003] = 29'b0_101001000001_011_0_100100000101;
      patterns[21004] = 29'b0_101001000001_100_1_010100100000;
      patterns[21005] = 29'b0_101001000001_101_0_101010010000;
      patterns[21006] = 29'b0_101001000001_110_0_101001000001;
      patterns[21007] = 29'b0_101001000001_111_0_101001000001;
      patterns[21008] = 29'b0_101001000010_000_0_101001000010;
      patterns[21009] = 29'b0_101001000010_001_0_000010101001;
      patterns[21010] = 29'b0_101001000010_010_1_010010000100;
      patterns[21011] = 29'b0_101001000010_011_0_100100001001;
      patterns[21012] = 29'b0_101001000010_100_0_010100100001;
      patterns[21013] = 29'b0_101001000010_101_1_001010010000;
      patterns[21014] = 29'b0_101001000010_110_0_101001000010;
      patterns[21015] = 29'b0_101001000010_111_0_101001000010;
      patterns[21016] = 29'b0_101001000011_000_0_101001000011;
      patterns[21017] = 29'b0_101001000011_001_0_000011101001;
      patterns[21018] = 29'b0_101001000011_010_1_010010000110;
      patterns[21019] = 29'b0_101001000011_011_0_100100001101;
      patterns[21020] = 29'b0_101001000011_100_1_010100100001;
      patterns[21021] = 29'b0_101001000011_101_1_101010010000;
      patterns[21022] = 29'b0_101001000011_110_0_101001000011;
      patterns[21023] = 29'b0_101001000011_111_0_101001000011;
      patterns[21024] = 29'b0_101001000100_000_0_101001000100;
      patterns[21025] = 29'b0_101001000100_001_0_000100101001;
      patterns[21026] = 29'b0_101001000100_010_1_010010001000;
      patterns[21027] = 29'b0_101001000100_011_0_100100010001;
      patterns[21028] = 29'b0_101001000100_100_0_010100100010;
      patterns[21029] = 29'b0_101001000100_101_0_001010010001;
      patterns[21030] = 29'b0_101001000100_110_0_101001000100;
      patterns[21031] = 29'b0_101001000100_111_0_101001000100;
      patterns[21032] = 29'b0_101001000101_000_0_101001000101;
      patterns[21033] = 29'b0_101001000101_001_0_000101101001;
      patterns[21034] = 29'b0_101001000101_010_1_010010001010;
      patterns[21035] = 29'b0_101001000101_011_0_100100010101;
      patterns[21036] = 29'b0_101001000101_100_1_010100100010;
      patterns[21037] = 29'b0_101001000101_101_0_101010010001;
      patterns[21038] = 29'b0_101001000101_110_0_101001000101;
      patterns[21039] = 29'b0_101001000101_111_0_101001000101;
      patterns[21040] = 29'b0_101001000110_000_0_101001000110;
      patterns[21041] = 29'b0_101001000110_001_0_000110101001;
      patterns[21042] = 29'b0_101001000110_010_1_010010001100;
      patterns[21043] = 29'b0_101001000110_011_0_100100011001;
      patterns[21044] = 29'b0_101001000110_100_0_010100100011;
      patterns[21045] = 29'b0_101001000110_101_1_001010010001;
      patterns[21046] = 29'b0_101001000110_110_0_101001000110;
      patterns[21047] = 29'b0_101001000110_111_0_101001000110;
      patterns[21048] = 29'b0_101001000111_000_0_101001000111;
      patterns[21049] = 29'b0_101001000111_001_0_000111101001;
      patterns[21050] = 29'b0_101001000111_010_1_010010001110;
      patterns[21051] = 29'b0_101001000111_011_0_100100011101;
      patterns[21052] = 29'b0_101001000111_100_1_010100100011;
      patterns[21053] = 29'b0_101001000111_101_1_101010010001;
      patterns[21054] = 29'b0_101001000111_110_0_101001000111;
      patterns[21055] = 29'b0_101001000111_111_0_101001000111;
      patterns[21056] = 29'b0_101001001000_000_0_101001001000;
      patterns[21057] = 29'b0_101001001000_001_0_001000101001;
      patterns[21058] = 29'b0_101001001000_010_1_010010010000;
      patterns[21059] = 29'b0_101001001000_011_0_100100100001;
      patterns[21060] = 29'b0_101001001000_100_0_010100100100;
      patterns[21061] = 29'b0_101001001000_101_0_001010010010;
      patterns[21062] = 29'b0_101001001000_110_0_101001001000;
      patterns[21063] = 29'b0_101001001000_111_0_101001001000;
      patterns[21064] = 29'b0_101001001001_000_0_101001001001;
      patterns[21065] = 29'b0_101001001001_001_0_001001101001;
      patterns[21066] = 29'b0_101001001001_010_1_010010010010;
      patterns[21067] = 29'b0_101001001001_011_0_100100100101;
      patterns[21068] = 29'b0_101001001001_100_1_010100100100;
      patterns[21069] = 29'b0_101001001001_101_0_101010010010;
      patterns[21070] = 29'b0_101001001001_110_0_101001001001;
      patterns[21071] = 29'b0_101001001001_111_0_101001001001;
      patterns[21072] = 29'b0_101001001010_000_0_101001001010;
      patterns[21073] = 29'b0_101001001010_001_0_001010101001;
      patterns[21074] = 29'b0_101001001010_010_1_010010010100;
      patterns[21075] = 29'b0_101001001010_011_0_100100101001;
      patterns[21076] = 29'b0_101001001010_100_0_010100100101;
      patterns[21077] = 29'b0_101001001010_101_1_001010010010;
      patterns[21078] = 29'b0_101001001010_110_0_101001001010;
      patterns[21079] = 29'b0_101001001010_111_0_101001001010;
      patterns[21080] = 29'b0_101001001011_000_0_101001001011;
      patterns[21081] = 29'b0_101001001011_001_0_001011101001;
      patterns[21082] = 29'b0_101001001011_010_1_010010010110;
      patterns[21083] = 29'b0_101001001011_011_0_100100101101;
      patterns[21084] = 29'b0_101001001011_100_1_010100100101;
      patterns[21085] = 29'b0_101001001011_101_1_101010010010;
      patterns[21086] = 29'b0_101001001011_110_0_101001001011;
      patterns[21087] = 29'b0_101001001011_111_0_101001001011;
      patterns[21088] = 29'b0_101001001100_000_0_101001001100;
      patterns[21089] = 29'b0_101001001100_001_0_001100101001;
      patterns[21090] = 29'b0_101001001100_010_1_010010011000;
      patterns[21091] = 29'b0_101001001100_011_0_100100110001;
      patterns[21092] = 29'b0_101001001100_100_0_010100100110;
      patterns[21093] = 29'b0_101001001100_101_0_001010010011;
      patterns[21094] = 29'b0_101001001100_110_0_101001001100;
      patterns[21095] = 29'b0_101001001100_111_0_101001001100;
      patterns[21096] = 29'b0_101001001101_000_0_101001001101;
      patterns[21097] = 29'b0_101001001101_001_0_001101101001;
      patterns[21098] = 29'b0_101001001101_010_1_010010011010;
      patterns[21099] = 29'b0_101001001101_011_0_100100110101;
      patterns[21100] = 29'b0_101001001101_100_1_010100100110;
      patterns[21101] = 29'b0_101001001101_101_0_101010010011;
      patterns[21102] = 29'b0_101001001101_110_0_101001001101;
      patterns[21103] = 29'b0_101001001101_111_0_101001001101;
      patterns[21104] = 29'b0_101001001110_000_0_101001001110;
      patterns[21105] = 29'b0_101001001110_001_0_001110101001;
      patterns[21106] = 29'b0_101001001110_010_1_010010011100;
      patterns[21107] = 29'b0_101001001110_011_0_100100111001;
      patterns[21108] = 29'b0_101001001110_100_0_010100100111;
      patterns[21109] = 29'b0_101001001110_101_1_001010010011;
      patterns[21110] = 29'b0_101001001110_110_0_101001001110;
      patterns[21111] = 29'b0_101001001110_111_0_101001001110;
      patterns[21112] = 29'b0_101001001111_000_0_101001001111;
      patterns[21113] = 29'b0_101001001111_001_0_001111101001;
      patterns[21114] = 29'b0_101001001111_010_1_010010011110;
      patterns[21115] = 29'b0_101001001111_011_0_100100111101;
      patterns[21116] = 29'b0_101001001111_100_1_010100100111;
      patterns[21117] = 29'b0_101001001111_101_1_101010010011;
      patterns[21118] = 29'b0_101001001111_110_0_101001001111;
      patterns[21119] = 29'b0_101001001111_111_0_101001001111;
      patterns[21120] = 29'b0_101001010000_000_0_101001010000;
      patterns[21121] = 29'b0_101001010000_001_0_010000101001;
      patterns[21122] = 29'b0_101001010000_010_1_010010100000;
      patterns[21123] = 29'b0_101001010000_011_0_100101000001;
      patterns[21124] = 29'b0_101001010000_100_0_010100101000;
      patterns[21125] = 29'b0_101001010000_101_0_001010010100;
      patterns[21126] = 29'b0_101001010000_110_0_101001010000;
      patterns[21127] = 29'b0_101001010000_111_0_101001010000;
      patterns[21128] = 29'b0_101001010001_000_0_101001010001;
      patterns[21129] = 29'b0_101001010001_001_0_010001101001;
      patterns[21130] = 29'b0_101001010001_010_1_010010100010;
      patterns[21131] = 29'b0_101001010001_011_0_100101000101;
      patterns[21132] = 29'b0_101001010001_100_1_010100101000;
      patterns[21133] = 29'b0_101001010001_101_0_101010010100;
      patterns[21134] = 29'b0_101001010001_110_0_101001010001;
      patterns[21135] = 29'b0_101001010001_111_0_101001010001;
      patterns[21136] = 29'b0_101001010010_000_0_101001010010;
      patterns[21137] = 29'b0_101001010010_001_0_010010101001;
      patterns[21138] = 29'b0_101001010010_010_1_010010100100;
      patterns[21139] = 29'b0_101001010010_011_0_100101001001;
      patterns[21140] = 29'b0_101001010010_100_0_010100101001;
      patterns[21141] = 29'b0_101001010010_101_1_001010010100;
      patterns[21142] = 29'b0_101001010010_110_0_101001010010;
      patterns[21143] = 29'b0_101001010010_111_0_101001010010;
      patterns[21144] = 29'b0_101001010011_000_0_101001010011;
      patterns[21145] = 29'b0_101001010011_001_0_010011101001;
      patterns[21146] = 29'b0_101001010011_010_1_010010100110;
      patterns[21147] = 29'b0_101001010011_011_0_100101001101;
      patterns[21148] = 29'b0_101001010011_100_1_010100101001;
      patterns[21149] = 29'b0_101001010011_101_1_101010010100;
      patterns[21150] = 29'b0_101001010011_110_0_101001010011;
      patterns[21151] = 29'b0_101001010011_111_0_101001010011;
      patterns[21152] = 29'b0_101001010100_000_0_101001010100;
      patterns[21153] = 29'b0_101001010100_001_0_010100101001;
      patterns[21154] = 29'b0_101001010100_010_1_010010101000;
      patterns[21155] = 29'b0_101001010100_011_0_100101010001;
      patterns[21156] = 29'b0_101001010100_100_0_010100101010;
      patterns[21157] = 29'b0_101001010100_101_0_001010010101;
      patterns[21158] = 29'b0_101001010100_110_0_101001010100;
      patterns[21159] = 29'b0_101001010100_111_0_101001010100;
      patterns[21160] = 29'b0_101001010101_000_0_101001010101;
      patterns[21161] = 29'b0_101001010101_001_0_010101101001;
      patterns[21162] = 29'b0_101001010101_010_1_010010101010;
      patterns[21163] = 29'b0_101001010101_011_0_100101010101;
      patterns[21164] = 29'b0_101001010101_100_1_010100101010;
      patterns[21165] = 29'b0_101001010101_101_0_101010010101;
      patterns[21166] = 29'b0_101001010101_110_0_101001010101;
      patterns[21167] = 29'b0_101001010101_111_0_101001010101;
      patterns[21168] = 29'b0_101001010110_000_0_101001010110;
      patterns[21169] = 29'b0_101001010110_001_0_010110101001;
      patterns[21170] = 29'b0_101001010110_010_1_010010101100;
      patterns[21171] = 29'b0_101001010110_011_0_100101011001;
      patterns[21172] = 29'b0_101001010110_100_0_010100101011;
      patterns[21173] = 29'b0_101001010110_101_1_001010010101;
      patterns[21174] = 29'b0_101001010110_110_0_101001010110;
      patterns[21175] = 29'b0_101001010110_111_0_101001010110;
      patterns[21176] = 29'b0_101001010111_000_0_101001010111;
      patterns[21177] = 29'b0_101001010111_001_0_010111101001;
      patterns[21178] = 29'b0_101001010111_010_1_010010101110;
      patterns[21179] = 29'b0_101001010111_011_0_100101011101;
      patterns[21180] = 29'b0_101001010111_100_1_010100101011;
      patterns[21181] = 29'b0_101001010111_101_1_101010010101;
      patterns[21182] = 29'b0_101001010111_110_0_101001010111;
      patterns[21183] = 29'b0_101001010111_111_0_101001010111;
      patterns[21184] = 29'b0_101001011000_000_0_101001011000;
      patterns[21185] = 29'b0_101001011000_001_0_011000101001;
      patterns[21186] = 29'b0_101001011000_010_1_010010110000;
      patterns[21187] = 29'b0_101001011000_011_0_100101100001;
      patterns[21188] = 29'b0_101001011000_100_0_010100101100;
      patterns[21189] = 29'b0_101001011000_101_0_001010010110;
      patterns[21190] = 29'b0_101001011000_110_0_101001011000;
      patterns[21191] = 29'b0_101001011000_111_0_101001011000;
      patterns[21192] = 29'b0_101001011001_000_0_101001011001;
      patterns[21193] = 29'b0_101001011001_001_0_011001101001;
      patterns[21194] = 29'b0_101001011001_010_1_010010110010;
      patterns[21195] = 29'b0_101001011001_011_0_100101100101;
      patterns[21196] = 29'b0_101001011001_100_1_010100101100;
      patterns[21197] = 29'b0_101001011001_101_0_101010010110;
      patterns[21198] = 29'b0_101001011001_110_0_101001011001;
      patterns[21199] = 29'b0_101001011001_111_0_101001011001;
      patterns[21200] = 29'b0_101001011010_000_0_101001011010;
      patterns[21201] = 29'b0_101001011010_001_0_011010101001;
      patterns[21202] = 29'b0_101001011010_010_1_010010110100;
      patterns[21203] = 29'b0_101001011010_011_0_100101101001;
      patterns[21204] = 29'b0_101001011010_100_0_010100101101;
      patterns[21205] = 29'b0_101001011010_101_1_001010010110;
      patterns[21206] = 29'b0_101001011010_110_0_101001011010;
      patterns[21207] = 29'b0_101001011010_111_0_101001011010;
      patterns[21208] = 29'b0_101001011011_000_0_101001011011;
      patterns[21209] = 29'b0_101001011011_001_0_011011101001;
      patterns[21210] = 29'b0_101001011011_010_1_010010110110;
      patterns[21211] = 29'b0_101001011011_011_0_100101101101;
      patterns[21212] = 29'b0_101001011011_100_1_010100101101;
      patterns[21213] = 29'b0_101001011011_101_1_101010010110;
      patterns[21214] = 29'b0_101001011011_110_0_101001011011;
      patterns[21215] = 29'b0_101001011011_111_0_101001011011;
      patterns[21216] = 29'b0_101001011100_000_0_101001011100;
      patterns[21217] = 29'b0_101001011100_001_0_011100101001;
      patterns[21218] = 29'b0_101001011100_010_1_010010111000;
      patterns[21219] = 29'b0_101001011100_011_0_100101110001;
      patterns[21220] = 29'b0_101001011100_100_0_010100101110;
      patterns[21221] = 29'b0_101001011100_101_0_001010010111;
      patterns[21222] = 29'b0_101001011100_110_0_101001011100;
      patterns[21223] = 29'b0_101001011100_111_0_101001011100;
      patterns[21224] = 29'b0_101001011101_000_0_101001011101;
      patterns[21225] = 29'b0_101001011101_001_0_011101101001;
      patterns[21226] = 29'b0_101001011101_010_1_010010111010;
      patterns[21227] = 29'b0_101001011101_011_0_100101110101;
      patterns[21228] = 29'b0_101001011101_100_1_010100101110;
      patterns[21229] = 29'b0_101001011101_101_0_101010010111;
      patterns[21230] = 29'b0_101001011101_110_0_101001011101;
      patterns[21231] = 29'b0_101001011101_111_0_101001011101;
      patterns[21232] = 29'b0_101001011110_000_0_101001011110;
      patterns[21233] = 29'b0_101001011110_001_0_011110101001;
      patterns[21234] = 29'b0_101001011110_010_1_010010111100;
      patterns[21235] = 29'b0_101001011110_011_0_100101111001;
      patterns[21236] = 29'b0_101001011110_100_0_010100101111;
      patterns[21237] = 29'b0_101001011110_101_1_001010010111;
      patterns[21238] = 29'b0_101001011110_110_0_101001011110;
      patterns[21239] = 29'b0_101001011110_111_0_101001011110;
      patterns[21240] = 29'b0_101001011111_000_0_101001011111;
      patterns[21241] = 29'b0_101001011111_001_0_011111101001;
      patterns[21242] = 29'b0_101001011111_010_1_010010111110;
      patterns[21243] = 29'b0_101001011111_011_0_100101111101;
      patterns[21244] = 29'b0_101001011111_100_1_010100101111;
      patterns[21245] = 29'b0_101001011111_101_1_101010010111;
      patterns[21246] = 29'b0_101001011111_110_0_101001011111;
      patterns[21247] = 29'b0_101001011111_111_0_101001011111;
      patterns[21248] = 29'b0_101001100000_000_0_101001100000;
      patterns[21249] = 29'b0_101001100000_001_0_100000101001;
      patterns[21250] = 29'b0_101001100000_010_1_010011000000;
      patterns[21251] = 29'b0_101001100000_011_0_100110000001;
      patterns[21252] = 29'b0_101001100000_100_0_010100110000;
      patterns[21253] = 29'b0_101001100000_101_0_001010011000;
      patterns[21254] = 29'b0_101001100000_110_0_101001100000;
      patterns[21255] = 29'b0_101001100000_111_0_101001100000;
      patterns[21256] = 29'b0_101001100001_000_0_101001100001;
      patterns[21257] = 29'b0_101001100001_001_0_100001101001;
      patterns[21258] = 29'b0_101001100001_010_1_010011000010;
      patterns[21259] = 29'b0_101001100001_011_0_100110000101;
      patterns[21260] = 29'b0_101001100001_100_1_010100110000;
      patterns[21261] = 29'b0_101001100001_101_0_101010011000;
      patterns[21262] = 29'b0_101001100001_110_0_101001100001;
      patterns[21263] = 29'b0_101001100001_111_0_101001100001;
      patterns[21264] = 29'b0_101001100010_000_0_101001100010;
      patterns[21265] = 29'b0_101001100010_001_0_100010101001;
      patterns[21266] = 29'b0_101001100010_010_1_010011000100;
      patterns[21267] = 29'b0_101001100010_011_0_100110001001;
      patterns[21268] = 29'b0_101001100010_100_0_010100110001;
      patterns[21269] = 29'b0_101001100010_101_1_001010011000;
      patterns[21270] = 29'b0_101001100010_110_0_101001100010;
      patterns[21271] = 29'b0_101001100010_111_0_101001100010;
      patterns[21272] = 29'b0_101001100011_000_0_101001100011;
      patterns[21273] = 29'b0_101001100011_001_0_100011101001;
      patterns[21274] = 29'b0_101001100011_010_1_010011000110;
      patterns[21275] = 29'b0_101001100011_011_0_100110001101;
      patterns[21276] = 29'b0_101001100011_100_1_010100110001;
      patterns[21277] = 29'b0_101001100011_101_1_101010011000;
      patterns[21278] = 29'b0_101001100011_110_0_101001100011;
      patterns[21279] = 29'b0_101001100011_111_0_101001100011;
      patterns[21280] = 29'b0_101001100100_000_0_101001100100;
      patterns[21281] = 29'b0_101001100100_001_0_100100101001;
      patterns[21282] = 29'b0_101001100100_010_1_010011001000;
      patterns[21283] = 29'b0_101001100100_011_0_100110010001;
      patterns[21284] = 29'b0_101001100100_100_0_010100110010;
      patterns[21285] = 29'b0_101001100100_101_0_001010011001;
      patterns[21286] = 29'b0_101001100100_110_0_101001100100;
      patterns[21287] = 29'b0_101001100100_111_0_101001100100;
      patterns[21288] = 29'b0_101001100101_000_0_101001100101;
      patterns[21289] = 29'b0_101001100101_001_0_100101101001;
      patterns[21290] = 29'b0_101001100101_010_1_010011001010;
      patterns[21291] = 29'b0_101001100101_011_0_100110010101;
      patterns[21292] = 29'b0_101001100101_100_1_010100110010;
      patterns[21293] = 29'b0_101001100101_101_0_101010011001;
      patterns[21294] = 29'b0_101001100101_110_0_101001100101;
      patterns[21295] = 29'b0_101001100101_111_0_101001100101;
      patterns[21296] = 29'b0_101001100110_000_0_101001100110;
      patterns[21297] = 29'b0_101001100110_001_0_100110101001;
      patterns[21298] = 29'b0_101001100110_010_1_010011001100;
      patterns[21299] = 29'b0_101001100110_011_0_100110011001;
      patterns[21300] = 29'b0_101001100110_100_0_010100110011;
      patterns[21301] = 29'b0_101001100110_101_1_001010011001;
      patterns[21302] = 29'b0_101001100110_110_0_101001100110;
      patterns[21303] = 29'b0_101001100110_111_0_101001100110;
      patterns[21304] = 29'b0_101001100111_000_0_101001100111;
      patterns[21305] = 29'b0_101001100111_001_0_100111101001;
      patterns[21306] = 29'b0_101001100111_010_1_010011001110;
      patterns[21307] = 29'b0_101001100111_011_0_100110011101;
      patterns[21308] = 29'b0_101001100111_100_1_010100110011;
      patterns[21309] = 29'b0_101001100111_101_1_101010011001;
      patterns[21310] = 29'b0_101001100111_110_0_101001100111;
      patterns[21311] = 29'b0_101001100111_111_0_101001100111;
      patterns[21312] = 29'b0_101001101000_000_0_101001101000;
      patterns[21313] = 29'b0_101001101000_001_0_101000101001;
      patterns[21314] = 29'b0_101001101000_010_1_010011010000;
      patterns[21315] = 29'b0_101001101000_011_0_100110100001;
      patterns[21316] = 29'b0_101001101000_100_0_010100110100;
      patterns[21317] = 29'b0_101001101000_101_0_001010011010;
      patterns[21318] = 29'b0_101001101000_110_0_101001101000;
      patterns[21319] = 29'b0_101001101000_111_0_101001101000;
      patterns[21320] = 29'b0_101001101001_000_0_101001101001;
      patterns[21321] = 29'b0_101001101001_001_0_101001101001;
      patterns[21322] = 29'b0_101001101001_010_1_010011010010;
      patterns[21323] = 29'b0_101001101001_011_0_100110100101;
      patterns[21324] = 29'b0_101001101001_100_1_010100110100;
      patterns[21325] = 29'b0_101001101001_101_0_101010011010;
      patterns[21326] = 29'b0_101001101001_110_0_101001101001;
      patterns[21327] = 29'b0_101001101001_111_0_101001101001;
      patterns[21328] = 29'b0_101001101010_000_0_101001101010;
      patterns[21329] = 29'b0_101001101010_001_0_101010101001;
      patterns[21330] = 29'b0_101001101010_010_1_010011010100;
      patterns[21331] = 29'b0_101001101010_011_0_100110101001;
      patterns[21332] = 29'b0_101001101010_100_0_010100110101;
      patterns[21333] = 29'b0_101001101010_101_1_001010011010;
      patterns[21334] = 29'b0_101001101010_110_0_101001101010;
      patterns[21335] = 29'b0_101001101010_111_0_101001101010;
      patterns[21336] = 29'b0_101001101011_000_0_101001101011;
      patterns[21337] = 29'b0_101001101011_001_0_101011101001;
      patterns[21338] = 29'b0_101001101011_010_1_010011010110;
      patterns[21339] = 29'b0_101001101011_011_0_100110101101;
      patterns[21340] = 29'b0_101001101011_100_1_010100110101;
      patterns[21341] = 29'b0_101001101011_101_1_101010011010;
      patterns[21342] = 29'b0_101001101011_110_0_101001101011;
      patterns[21343] = 29'b0_101001101011_111_0_101001101011;
      patterns[21344] = 29'b0_101001101100_000_0_101001101100;
      patterns[21345] = 29'b0_101001101100_001_0_101100101001;
      patterns[21346] = 29'b0_101001101100_010_1_010011011000;
      patterns[21347] = 29'b0_101001101100_011_0_100110110001;
      patterns[21348] = 29'b0_101001101100_100_0_010100110110;
      patterns[21349] = 29'b0_101001101100_101_0_001010011011;
      patterns[21350] = 29'b0_101001101100_110_0_101001101100;
      patterns[21351] = 29'b0_101001101100_111_0_101001101100;
      patterns[21352] = 29'b0_101001101101_000_0_101001101101;
      patterns[21353] = 29'b0_101001101101_001_0_101101101001;
      patterns[21354] = 29'b0_101001101101_010_1_010011011010;
      patterns[21355] = 29'b0_101001101101_011_0_100110110101;
      patterns[21356] = 29'b0_101001101101_100_1_010100110110;
      patterns[21357] = 29'b0_101001101101_101_0_101010011011;
      patterns[21358] = 29'b0_101001101101_110_0_101001101101;
      patterns[21359] = 29'b0_101001101101_111_0_101001101101;
      patterns[21360] = 29'b0_101001101110_000_0_101001101110;
      patterns[21361] = 29'b0_101001101110_001_0_101110101001;
      patterns[21362] = 29'b0_101001101110_010_1_010011011100;
      patterns[21363] = 29'b0_101001101110_011_0_100110111001;
      patterns[21364] = 29'b0_101001101110_100_0_010100110111;
      patterns[21365] = 29'b0_101001101110_101_1_001010011011;
      patterns[21366] = 29'b0_101001101110_110_0_101001101110;
      patterns[21367] = 29'b0_101001101110_111_0_101001101110;
      patterns[21368] = 29'b0_101001101111_000_0_101001101111;
      patterns[21369] = 29'b0_101001101111_001_0_101111101001;
      patterns[21370] = 29'b0_101001101111_010_1_010011011110;
      patterns[21371] = 29'b0_101001101111_011_0_100110111101;
      patterns[21372] = 29'b0_101001101111_100_1_010100110111;
      patterns[21373] = 29'b0_101001101111_101_1_101010011011;
      patterns[21374] = 29'b0_101001101111_110_0_101001101111;
      patterns[21375] = 29'b0_101001101111_111_0_101001101111;
      patterns[21376] = 29'b0_101001110000_000_0_101001110000;
      patterns[21377] = 29'b0_101001110000_001_0_110000101001;
      patterns[21378] = 29'b0_101001110000_010_1_010011100000;
      patterns[21379] = 29'b0_101001110000_011_0_100111000001;
      patterns[21380] = 29'b0_101001110000_100_0_010100111000;
      patterns[21381] = 29'b0_101001110000_101_0_001010011100;
      patterns[21382] = 29'b0_101001110000_110_0_101001110000;
      patterns[21383] = 29'b0_101001110000_111_0_101001110000;
      patterns[21384] = 29'b0_101001110001_000_0_101001110001;
      patterns[21385] = 29'b0_101001110001_001_0_110001101001;
      patterns[21386] = 29'b0_101001110001_010_1_010011100010;
      patterns[21387] = 29'b0_101001110001_011_0_100111000101;
      patterns[21388] = 29'b0_101001110001_100_1_010100111000;
      patterns[21389] = 29'b0_101001110001_101_0_101010011100;
      patterns[21390] = 29'b0_101001110001_110_0_101001110001;
      patterns[21391] = 29'b0_101001110001_111_0_101001110001;
      patterns[21392] = 29'b0_101001110010_000_0_101001110010;
      patterns[21393] = 29'b0_101001110010_001_0_110010101001;
      patterns[21394] = 29'b0_101001110010_010_1_010011100100;
      patterns[21395] = 29'b0_101001110010_011_0_100111001001;
      patterns[21396] = 29'b0_101001110010_100_0_010100111001;
      patterns[21397] = 29'b0_101001110010_101_1_001010011100;
      patterns[21398] = 29'b0_101001110010_110_0_101001110010;
      patterns[21399] = 29'b0_101001110010_111_0_101001110010;
      patterns[21400] = 29'b0_101001110011_000_0_101001110011;
      patterns[21401] = 29'b0_101001110011_001_0_110011101001;
      patterns[21402] = 29'b0_101001110011_010_1_010011100110;
      patterns[21403] = 29'b0_101001110011_011_0_100111001101;
      patterns[21404] = 29'b0_101001110011_100_1_010100111001;
      patterns[21405] = 29'b0_101001110011_101_1_101010011100;
      patterns[21406] = 29'b0_101001110011_110_0_101001110011;
      patterns[21407] = 29'b0_101001110011_111_0_101001110011;
      patterns[21408] = 29'b0_101001110100_000_0_101001110100;
      patterns[21409] = 29'b0_101001110100_001_0_110100101001;
      patterns[21410] = 29'b0_101001110100_010_1_010011101000;
      patterns[21411] = 29'b0_101001110100_011_0_100111010001;
      patterns[21412] = 29'b0_101001110100_100_0_010100111010;
      patterns[21413] = 29'b0_101001110100_101_0_001010011101;
      patterns[21414] = 29'b0_101001110100_110_0_101001110100;
      patterns[21415] = 29'b0_101001110100_111_0_101001110100;
      patterns[21416] = 29'b0_101001110101_000_0_101001110101;
      patterns[21417] = 29'b0_101001110101_001_0_110101101001;
      patterns[21418] = 29'b0_101001110101_010_1_010011101010;
      patterns[21419] = 29'b0_101001110101_011_0_100111010101;
      patterns[21420] = 29'b0_101001110101_100_1_010100111010;
      patterns[21421] = 29'b0_101001110101_101_0_101010011101;
      patterns[21422] = 29'b0_101001110101_110_0_101001110101;
      patterns[21423] = 29'b0_101001110101_111_0_101001110101;
      patterns[21424] = 29'b0_101001110110_000_0_101001110110;
      patterns[21425] = 29'b0_101001110110_001_0_110110101001;
      patterns[21426] = 29'b0_101001110110_010_1_010011101100;
      patterns[21427] = 29'b0_101001110110_011_0_100111011001;
      patterns[21428] = 29'b0_101001110110_100_0_010100111011;
      patterns[21429] = 29'b0_101001110110_101_1_001010011101;
      patterns[21430] = 29'b0_101001110110_110_0_101001110110;
      patterns[21431] = 29'b0_101001110110_111_0_101001110110;
      patterns[21432] = 29'b0_101001110111_000_0_101001110111;
      patterns[21433] = 29'b0_101001110111_001_0_110111101001;
      patterns[21434] = 29'b0_101001110111_010_1_010011101110;
      patterns[21435] = 29'b0_101001110111_011_0_100111011101;
      patterns[21436] = 29'b0_101001110111_100_1_010100111011;
      patterns[21437] = 29'b0_101001110111_101_1_101010011101;
      patterns[21438] = 29'b0_101001110111_110_0_101001110111;
      patterns[21439] = 29'b0_101001110111_111_0_101001110111;
      patterns[21440] = 29'b0_101001111000_000_0_101001111000;
      patterns[21441] = 29'b0_101001111000_001_0_111000101001;
      patterns[21442] = 29'b0_101001111000_010_1_010011110000;
      patterns[21443] = 29'b0_101001111000_011_0_100111100001;
      patterns[21444] = 29'b0_101001111000_100_0_010100111100;
      patterns[21445] = 29'b0_101001111000_101_0_001010011110;
      patterns[21446] = 29'b0_101001111000_110_0_101001111000;
      patterns[21447] = 29'b0_101001111000_111_0_101001111000;
      patterns[21448] = 29'b0_101001111001_000_0_101001111001;
      patterns[21449] = 29'b0_101001111001_001_0_111001101001;
      patterns[21450] = 29'b0_101001111001_010_1_010011110010;
      patterns[21451] = 29'b0_101001111001_011_0_100111100101;
      patterns[21452] = 29'b0_101001111001_100_1_010100111100;
      patterns[21453] = 29'b0_101001111001_101_0_101010011110;
      patterns[21454] = 29'b0_101001111001_110_0_101001111001;
      patterns[21455] = 29'b0_101001111001_111_0_101001111001;
      patterns[21456] = 29'b0_101001111010_000_0_101001111010;
      patterns[21457] = 29'b0_101001111010_001_0_111010101001;
      patterns[21458] = 29'b0_101001111010_010_1_010011110100;
      patterns[21459] = 29'b0_101001111010_011_0_100111101001;
      patterns[21460] = 29'b0_101001111010_100_0_010100111101;
      patterns[21461] = 29'b0_101001111010_101_1_001010011110;
      patterns[21462] = 29'b0_101001111010_110_0_101001111010;
      patterns[21463] = 29'b0_101001111010_111_0_101001111010;
      patterns[21464] = 29'b0_101001111011_000_0_101001111011;
      patterns[21465] = 29'b0_101001111011_001_0_111011101001;
      patterns[21466] = 29'b0_101001111011_010_1_010011110110;
      patterns[21467] = 29'b0_101001111011_011_0_100111101101;
      patterns[21468] = 29'b0_101001111011_100_1_010100111101;
      patterns[21469] = 29'b0_101001111011_101_1_101010011110;
      patterns[21470] = 29'b0_101001111011_110_0_101001111011;
      patterns[21471] = 29'b0_101001111011_111_0_101001111011;
      patterns[21472] = 29'b0_101001111100_000_0_101001111100;
      patterns[21473] = 29'b0_101001111100_001_0_111100101001;
      patterns[21474] = 29'b0_101001111100_010_1_010011111000;
      patterns[21475] = 29'b0_101001111100_011_0_100111110001;
      patterns[21476] = 29'b0_101001111100_100_0_010100111110;
      patterns[21477] = 29'b0_101001111100_101_0_001010011111;
      patterns[21478] = 29'b0_101001111100_110_0_101001111100;
      patterns[21479] = 29'b0_101001111100_111_0_101001111100;
      patterns[21480] = 29'b0_101001111101_000_0_101001111101;
      patterns[21481] = 29'b0_101001111101_001_0_111101101001;
      patterns[21482] = 29'b0_101001111101_010_1_010011111010;
      patterns[21483] = 29'b0_101001111101_011_0_100111110101;
      patterns[21484] = 29'b0_101001111101_100_1_010100111110;
      patterns[21485] = 29'b0_101001111101_101_0_101010011111;
      patterns[21486] = 29'b0_101001111101_110_0_101001111101;
      patterns[21487] = 29'b0_101001111101_111_0_101001111101;
      patterns[21488] = 29'b0_101001111110_000_0_101001111110;
      patterns[21489] = 29'b0_101001111110_001_0_111110101001;
      patterns[21490] = 29'b0_101001111110_010_1_010011111100;
      patterns[21491] = 29'b0_101001111110_011_0_100111111001;
      patterns[21492] = 29'b0_101001111110_100_0_010100111111;
      patterns[21493] = 29'b0_101001111110_101_1_001010011111;
      patterns[21494] = 29'b0_101001111110_110_0_101001111110;
      patterns[21495] = 29'b0_101001111110_111_0_101001111110;
      patterns[21496] = 29'b0_101001111111_000_0_101001111111;
      patterns[21497] = 29'b0_101001111111_001_0_111111101001;
      patterns[21498] = 29'b0_101001111111_010_1_010011111110;
      patterns[21499] = 29'b0_101001111111_011_0_100111111101;
      patterns[21500] = 29'b0_101001111111_100_1_010100111111;
      patterns[21501] = 29'b0_101001111111_101_1_101010011111;
      patterns[21502] = 29'b0_101001111111_110_0_101001111111;
      patterns[21503] = 29'b0_101001111111_111_0_101001111111;
      patterns[21504] = 29'b0_101010000000_000_0_101010000000;
      patterns[21505] = 29'b0_101010000000_001_0_000000101010;
      patterns[21506] = 29'b0_101010000000_010_1_010100000000;
      patterns[21507] = 29'b0_101010000000_011_0_101000000001;
      patterns[21508] = 29'b0_101010000000_100_0_010101000000;
      patterns[21509] = 29'b0_101010000000_101_0_001010100000;
      patterns[21510] = 29'b0_101010000000_110_0_101010000000;
      patterns[21511] = 29'b0_101010000000_111_0_101010000000;
      patterns[21512] = 29'b0_101010000001_000_0_101010000001;
      patterns[21513] = 29'b0_101010000001_001_0_000001101010;
      patterns[21514] = 29'b0_101010000001_010_1_010100000010;
      patterns[21515] = 29'b0_101010000001_011_0_101000000101;
      patterns[21516] = 29'b0_101010000001_100_1_010101000000;
      patterns[21517] = 29'b0_101010000001_101_0_101010100000;
      patterns[21518] = 29'b0_101010000001_110_0_101010000001;
      patterns[21519] = 29'b0_101010000001_111_0_101010000001;
      patterns[21520] = 29'b0_101010000010_000_0_101010000010;
      patterns[21521] = 29'b0_101010000010_001_0_000010101010;
      patterns[21522] = 29'b0_101010000010_010_1_010100000100;
      patterns[21523] = 29'b0_101010000010_011_0_101000001001;
      patterns[21524] = 29'b0_101010000010_100_0_010101000001;
      patterns[21525] = 29'b0_101010000010_101_1_001010100000;
      patterns[21526] = 29'b0_101010000010_110_0_101010000010;
      patterns[21527] = 29'b0_101010000010_111_0_101010000010;
      patterns[21528] = 29'b0_101010000011_000_0_101010000011;
      patterns[21529] = 29'b0_101010000011_001_0_000011101010;
      patterns[21530] = 29'b0_101010000011_010_1_010100000110;
      patterns[21531] = 29'b0_101010000011_011_0_101000001101;
      patterns[21532] = 29'b0_101010000011_100_1_010101000001;
      patterns[21533] = 29'b0_101010000011_101_1_101010100000;
      patterns[21534] = 29'b0_101010000011_110_0_101010000011;
      patterns[21535] = 29'b0_101010000011_111_0_101010000011;
      patterns[21536] = 29'b0_101010000100_000_0_101010000100;
      patterns[21537] = 29'b0_101010000100_001_0_000100101010;
      patterns[21538] = 29'b0_101010000100_010_1_010100001000;
      patterns[21539] = 29'b0_101010000100_011_0_101000010001;
      patterns[21540] = 29'b0_101010000100_100_0_010101000010;
      patterns[21541] = 29'b0_101010000100_101_0_001010100001;
      patterns[21542] = 29'b0_101010000100_110_0_101010000100;
      patterns[21543] = 29'b0_101010000100_111_0_101010000100;
      patterns[21544] = 29'b0_101010000101_000_0_101010000101;
      patterns[21545] = 29'b0_101010000101_001_0_000101101010;
      patterns[21546] = 29'b0_101010000101_010_1_010100001010;
      patterns[21547] = 29'b0_101010000101_011_0_101000010101;
      patterns[21548] = 29'b0_101010000101_100_1_010101000010;
      patterns[21549] = 29'b0_101010000101_101_0_101010100001;
      patterns[21550] = 29'b0_101010000101_110_0_101010000101;
      patterns[21551] = 29'b0_101010000101_111_0_101010000101;
      patterns[21552] = 29'b0_101010000110_000_0_101010000110;
      patterns[21553] = 29'b0_101010000110_001_0_000110101010;
      patterns[21554] = 29'b0_101010000110_010_1_010100001100;
      patterns[21555] = 29'b0_101010000110_011_0_101000011001;
      patterns[21556] = 29'b0_101010000110_100_0_010101000011;
      patterns[21557] = 29'b0_101010000110_101_1_001010100001;
      patterns[21558] = 29'b0_101010000110_110_0_101010000110;
      patterns[21559] = 29'b0_101010000110_111_0_101010000110;
      patterns[21560] = 29'b0_101010000111_000_0_101010000111;
      patterns[21561] = 29'b0_101010000111_001_0_000111101010;
      patterns[21562] = 29'b0_101010000111_010_1_010100001110;
      patterns[21563] = 29'b0_101010000111_011_0_101000011101;
      patterns[21564] = 29'b0_101010000111_100_1_010101000011;
      patterns[21565] = 29'b0_101010000111_101_1_101010100001;
      patterns[21566] = 29'b0_101010000111_110_0_101010000111;
      patterns[21567] = 29'b0_101010000111_111_0_101010000111;
      patterns[21568] = 29'b0_101010001000_000_0_101010001000;
      patterns[21569] = 29'b0_101010001000_001_0_001000101010;
      patterns[21570] = 29'b0_101010001000_010_1_010100010000;
      patterns[21571] = 29'b0_101010001000_011_0_101000100001;
      patterns[21572] = 29'b0_101010001000_100_0_010101000100;
      patterns[21573] = 29'b0_101010001000_101_0_001010100010;
      patterns[21574] = 29'b0_101010001000_110_0_101010001000;
      patterns[21575] = 29'b0_101010001000_111_0_101010001000;
      patterns[21576] = 29'b0_101010001001_000_0_101010001001;
      patterns[21577] = 29'b0_101010001001_001_0_001001101010;
      patterns[21578] = 29'b0_101010001001_010_1_010100010010;
      patterns[21579] = 29'b0_101010001001_011_0_101000100101;
      patterns[21580] = 29'b0_101010001001_100_1_010101000100;
      patterns[21581] = 29'b0_101010001001_101_0_101010100010;
      patterns[21582] = 29'b0_101010001001_110_0_101010001001;
      patterns[21583] = 29'b0_101010001001_111_0_101010001001;
      patterns[21584] = 29'b0_101010001010_000_0_101010001010;
      patterns[21585] = 29'b0_101010001010_001_0_001010101010;
      patterns[21586] = 29'b0_101010001010_010_1_010100010100;
      patterns[21587] = 29'b0_101010001010_011_0_101000101001;
      patterns[21588] = 29'b0_101010001010_100_0_010101000101;
      patterns[21589] = 29'b0_101010001010_101_1_001010100010;
      patterns[21590] = 29'b0_101010001010_110_0_101010001010;
      patterns[21591] = 29'b0_101010001010_111_0_101010001010;
      patterns[21592] = 29'b0_101010001011_000_0_101010001011;
      patterns[21593] = 29'b0_101010001011_001_0_001011101010;
      patterns[21594] = 29'b0_101010001011_010_1_010100010110;
      patterns[21595] = 29'b0_101010001011_011_0_101000101101;
      patterns[21596] = 29'b0_101010001011_100_1_010101000101;
      patterns[21597] = 29'b0_101010001011_101_1_101010100010;
      patterns[21598] = 29'b0_101010001011_110_0_101010001011;
      patterns[21599] = 29'b0_101010001011_111_0_101010001011;
      patterns[21600] = 29'b0_101010001100_000_0_101010001100;
      patterns[21601] = 29'b0_101010001100_001_0_001100101010;
      patterns[21602] = 29'b0_101010001100_010_1_010100011000;
      patterns[21603] = 29'b0_101010001100_011_0_101000110001;
      patterns[21604] = 29'b0_101010001100_100_0_010101000110;
      patterns[21605] = 29'b0_101010001100_101_0_001010100011;
      patterns[21606] = 29'b0_101010001100_110_0_101010001100;
      patterns[21607] = 29'b0_101010001100_111_0_101010001100;
      patterns[21608] = 29'b0_101010001101_000_0_101010001101;
      patterns[21609] = 29'b0_101010001101_001_0_001101101010;
      patterns[21610] = 29'b0_101010001101_010_1_010100011010;
      patterns[21611] = 29'b0_101010001101_011_0_101000110101;
      patterns[21612] = 29'b0_101010001101_100_1_010101000110;
      patterns[21613] = 29'b0_101010001101_101_0_101010100011;
      patterns[21614] = 29'b0_101010001101_110_0_101010001101;
      patterns[21615] = 29'b0_101010001101_111_0_101010001101;
      patterns[21616] = 29'b0_101010001110_000_0_101010001110;
      patterns[21617] = 29'b0_101010001110_001_0_001110101010;
      patterns[21618] = 29'b0_101010001110_010_1_010100011100;
      patterns[21619] = 29'b0_101010001110_011_0_101000111001;
      patterns[21620] = 29'b0_101010001110_100_0_010101000111;
      patterns[21621] = 29'b0_101010001110_101_1_001010100011;
      patterns[21622] = 29'b0_101010001110_110_0_101010001110;
      patterns[21623] = 29'b0_101010001110_111_0_101010001110;
      patterns[21624] = 29'b0_101010001111_000_0_101010001111;
      patterns[21625] = 29'b0_101010001111_001_0_001111101010;
      patterns[21626] = 29'b0_101010001111_010_1_010100011110;
      patterns[21627] = 29'b0_101010001111_011_0_101000111101;
      patterns[21628] = 29'b0_101010001111_100_1_010101000111;
      patterns[21629] = 29'b0_101010001111_101_1_101010100011;
      patterns[21630] = 29'b0_101010001111_110_0_101010001111;
      patterns[21631] = 29'b0_101010001111_111_0_101010001111;
      patterns[21632] = 29'b0_101010010000_000_0_101010010000;
      patterns[21633] = 29'b0_101010010000_001_0_010000101010;
      patterns[21634] = 29'b0_101010010000_010_1_010100100000;
      patterns[21635] = 29'b0_101010010000_011_0_101001000001;
      patterns[21636] = 29'b0_101010010000_100_0_010101001000;
      patterns[21637] = 29'b0_101010010000_101_0_001010100100;
      patterns[21638] = 29'b0_101010010000_110_0_101010010000;
      patterns[21639] = 29'b0_101010010000_111_0_101010010000;
      patterns[21640] = 29'b0_101010010001_000_0_101010010001;
      patterns[21641] = 29'b0_101010010001_001_0_010001101010;
      patterns[21642] = 29'b0_101010010001_010_1_010100100010;
      patterns[21643] = 29'b0_101010010001_011_0_101001000101;
      patterns[21644] = 29'b0_101010010001_100_1_010101001000;
      patterns[21645] = 29'b0_101010010001_101_0_101010100100;
      patterns[21646] = 29'b0_101010010001_110_0_101010010001;
      patterns[21647] = 29'b0_101010010001_111_0_101010010001;
      patterns[21648] = 29'b0_101010010010_000_0_101010010010;
      patterns[21649] = 29'b0_101010010010_001_0_010010101010;
      patterns[21650] = 29'b0_101010010010_010_1_010100100100;
      patterns[21651] = 29'b0_101010010010_011_0_101001001001;
      patterns[21652] = 29'b0_101010010010_100_0_010101001001;
      patterns[21653] = 29'b0_101010010010_101_1_001010100100;
      patterns[21654] = 29'b0_101010010010_110_0_101010010010;
      patterns[21655] = 29'b0_101010010010_111_0_101010010010;
      patterns[21656] = 29'b0_101010010011_000_0_101010010011;
      patterns[21657] = 29'b0_101010010011_001_0_010011101010;
      patterns[21658] = 29'b0_101010010011_010_1_010100100110;
      patterns[21659] = 29'b0_101010010011_011_0_101001001101;
      patterns[21660] = 29'b0_101010010011_100_1_010101001001;
      patterns[21661] = 29'b0_101010010011_101_1_101010100100;
      patterns[21662] = 29'b0_101010010011_110_0_101010010011;
      patterns[21663] = 29'b0_101010010011_111_0_101010010011;
      patterns[21664] = 29'b0_101010010100_000_0_101010010100;
      patterns[21665] = 29'b0_101010010100_001_0_010100101010;
      patterns[21666] = 29'b0_101010010100_010_1_010100101000;
      patterns[21667] = 29'b0_101010010100_011_0_101001010001;
      patterns[21668] = 29'b0_101010010100_100_0_010101001010;
      patterns[21669] = 29'b0_101010010100_101_0_001010100101;
      patterns[21670] = 29'b0_101010010100_110_0_101010010100;
      patterns[21671] = 29'b0_101010010100_111_0_101010010100;
      patterns[21672] = 29'b0_101010010101_000_0_101010010101;
      patterns[21673] = 29'b0_101010010101_001_0_010101101010;
      patterns[21674] = 29'b0_101010010101_010_1_010100101010;
      patterns[21675] = 29'b0_101010010101_011_0_101001010101;
      patterns[21676] = 29'b0_101010010101_100_1_010101001010;
      patterns[21677] = 29'b0_101010010101_101_0_101010100101;
      patterns[21678] = 29'b0_101010010101_110_0_101010010101;
      patterns[21679] = 29'b0_101010010101_111_0_101010010101;
      patterns[21680] = 29'b0_101010010110_000_0_101010010110;
      patterns[21681] = 29'b0_101010010110_001_0_010110101010;
      patterns[21682] = 29'b0_101010010110_010_1_010100101100;
      patterns[21683] = 29'b0_101010010110_011_0_101001011001;
      patterns[21684] = 29'b0_101010010110_100_0_010101001011;
      patterns[21685] = 29'b0_101010010110_101_1_001010100101;
      patterns[21686] = 29'b0_101010010110_110_0_101010010110;
      patterns[21687] = 29'b0_101010010110_111_0_101010010110;
      patterns[21688] = 29'b0_101010010111_000_0_101010010111;
      patterns[21689] = 29'b0_101010010111_001_0_010111101010;
      patterns[21690] = 29'b0_101010010111_010_1_010100101110;
      patterns[21691] = 29'b0_101010010111_011_0_101001011101;
      patterns[21692] = 29'b0_101010010111_100_1_010101001011;
      patterns[21693] = 29'b0_101010010111_101_1_101010100101;
      patterns[21694] = 29'b0_101010010111_110_0_101010010111;
      patterns[21695] = 29'b0_101010010111_111_0_101010010111;
      patterns[21696] = 29'b0_101010011000_000_0_101010011000;
      patterns[21697] = 29'b0_101010011000_001_0_011000101010;
      patterns[21698] = 29'b0_101010011000_010_1_010100110000;
      patterns[21699] = 29'b0_101010011000_011_0_101001100001;
      patterns[21700] = 29'b0_101010011000_100_0_010101001100;
      patterns[21701] = 29'b0_101010011000_101_0_001010100110;
      patterns[21702] = 29'b0_101010011000_110_0_101010011000;
      patterns[21703] = 29'b0_101010011000_111_0_101010011000;
      patterns[21704] = 29'b0_101010011001_000_0_101010011001;
      patterns[21705] = 29'b0_101010011001_001_0_011001101010;
      patterns[21706] = 29'b0_101010011001_010_1_010100110010;
      patterns[21707] = 29'b0_101010011001_011_0_101001100101;
      patterns[21708] = 29'b0_101010011001_100_1_010101001100;
      patterns[21709] = 29'b0_101010011001_101_0_101010100110;
      patterns[21710] = 29'b0_101010011001_110_0_101010011001;
      patterns[21711] = 29'b0_101010011001_111_0_101010011001;
      patterns[21712] = 29'b0_101010011010_000_0_101010011010;
      patterns[21713] = 29'b0_101010011010_001_0_011010101010;
      patterns[21714] = 29'b0_101010011010_010_1_010100110100;
      patterns[21715] = 29'b0_101010011010_011_0_101001101001;
      patterns[21716] = 29'b0_101010011010_100_0_010101001101;
      patterns[21717] = 29'b0_101010011010_101_1_001010100110;
      patterns[21718] = 29'b0_101010011010_110_0_101010011010;
      patterns[21719] = 29'b0_101010011010_111_0_101010011010;
      patterns[21720] = 29'b0_101010011011_000_0_101010011011;
      patterns[21721] = 29'b0_101010011011_001_0_011011101010;
      patterns[21722] = 29'b0_101010011011_010_1_010100110110;
      patterns[21723] = 29'b0_101010011011_011_0_101001101101;
      patterns[21724] = 29'b0_101010011011_100_1_010101001101;
      patterns[21725] = 29'b0_101010011011_101_1_101010100110;
      patterns[21726] = 29'b0_101010011011_110_0_101010011011;
      patterns[21727] = 29'b0_101010011011_111_0_101010011011;
      patterns[21728] = 29'b0_101010011100_000_0_101010011100;
      patterns[21729] = 29'b0_101010011100_001_0_011100101010;
      patterns[21730] = 29'b0_101010011100_010_1_010100111000;
      patterns[21731] = 29'b0_101010011100_011_0_101001110001;
      patterns[21732] = 29'b0_101010011100_100_0_010101001110;
      patterns[21733] = 29'b0_101010011100_101_0_001010100111;
      patterns[21734] = 29'b0_101010011100_110_0_101010011100;
      patterns[21735] = 29'b0_101010011100_111_0_101010011100;
      patterns[21736] = 29'b0_101010011101_000_0_101010011101;
      patterns[21737] = 29'b0_101010011101_001_0_011101101010;
      patterns[21738] = 29'b0_101010011101_010_1_010100111010;
      patterns[21739] = 29'b0_101010011101_011_0_101001110101;
      patterns[21740] = 29'b0_101010011101_100_1_010101001110;
      patterns[21741] = 29'b0_101010011101_101_0_101010100111;
      patterns[21742] = 29'b0_101010011101_110_0_101010011101;
      patterns[21743] = 29'b0_101010011101_111_0_101010011101;
      patterns[21744] = 29'b0_101010011110_000_0_101010011110;
      patterns[21745] = 29'b0_101010011110_001_0_011110101010;
      patterns[21746] = 29'b0_101010011110_010_1_010100111100;
      patterns[21747] = 29'b0_101010011110_011_0_101001111001;
      patterns[21748] = 29'b0_101010011110_100_0_010101001111;
      patterns[21749] = 29'b0_101010011110_101_1_001010100111;
      patterns[21750] = 29'b0_101010011110_110_0_101010011110;
      patterns[21751] = 29'b0_101010011110_111_0_101010011110;
      patterns[21752] = 29'b0_101010011111_000_0_101010011111;
      patterns[21753] = 29'b0_101010011111_001_0_011111101010;
      patterns[21754] = 29'b0_101010011111_010_1_010100111110;
      patterns[21755] = 29'b0_101010011111_011_0_101001111101;
      patterns[21756] = 29'b0_101010011111_100_1_010101001111;
      patterns[21757] = 29'b0_101010011111_101_1_101010100111;
      patterns[21758] = 29'b0_101010011111_110_0_101010011111;
      patterns[21759] = 29'b0_101010011111_111_0_101010011111;
      patterns[21760] = 29'b0_101010100000_000_0_101010100000;
      patterns[21761] = 29'b0_101010100000_001_0_100000101010;
      patterns[21762] = 29'b0_101010100000_010_1_010101000000;
      patterns[21763] = 29'b0_101010100000_011_0_101010000001;
      patterns[21764] = 29'b0_101010100000_100_0_010101010000;
      patterns[21765] = 29'b0_101010100000_101_0_001010101000;
      patterns[21766] = 29'b0_101010100000_110_0_101010100000;
      patterns[21767] = 29'b0_101010100000_111_0_101010100000;
      patterns[21768] = 29'b0_101010100001_000_0_101010100001;
      patterns[21769] = 29'b0_101010100001_001_0_100001101010;
      patterns[21770] = 29'b0_101010100001_010_1_010101000010;
      patterns[21771] = 29'b0_101010100001_011_0_101010000101;
      patterns[21772] = 29'b0_101010100001_100_1_010101010000;
      patterns[21773] = 29'b0_101010100001_101_0_101010101000;
      patterns[21774] = 29'b0_101010100001_110_0_101010100001;
      patterns[21775] = 29'b0_101010100001_111_0_101010100001;
      patterns[21776] = 29'b0_101010100010_000_0_101010100010;
      patterns[21777] = 29'b0_101010100010_001_0_100010101010;
      patterns[21778] = 29'b0_101010100010_010_1_010101000100;
      patterns[21779] = 29'b0_101010100010_011_0_101010001001;
      patterns[21780] = 29'b0_101010100010_100_0_010101010001;
      patterns[21781] = 29'b0_101010100010_101_1_001010101000;
      patterns[21782] = 29'b0_101010100010_110_0_101010100010;
      patterns[21783] = 29'b0_101010100010_111_0_101010100010;
      patterns[21784] = 29'b0_101010100011_000_0_101010100011;
      patterns[21785] = 29'b0_101010100011_001_0_100011101010;
      patterns[21786] = 29'b0_101010100011_010_1_010101000110;
      patterns[21787] = 29'b0_101010100011_011_0_101010001101;
      patterns[21788] = 29'b0_101010100011_100_1_010101010001;
      patterns[21789] = 29'b0_101010100011_101_1_101010101000;
      patterns[21790] = 29'b0_101010100011_110_0_101010100011;
      patterns[21791] = 29'b0_101010100011_111_0_101010100011;
      patterns[21792] = 29'b0_101010100100_000_0_101010100100;
      patterns[21793] = 29'b0_101010100100_001_0_100100101010;
      patterns[21794] = 29'b0_101010100100_010_1_010101001000;
      patterns[21795] = 29'b0_101010100100_011_0_101010010001;
      patterns[21796] = 29'b0_101010100100_100_0_010101010010;
      patterns[21797] = 29'b0_101010100100_101_0_001010101001;
      patterns[21798] = 29'b0_101010100100_110_0_101010100100;
      patterns[21799] = 29'b0_101010100100_111_0_101010100100;
      patterns[21800] = 29'b0_101010100101_000_0_101010100101;
      patterns[21801] = 29'b0_101010100101_001_0_100101101010;
      patterns[21802] = 29'b0_101010100101_010_1_010101001010;
      patterns[21803] = 29'b0_101010100101_011_0_101010010101;
      patterns[21804] = 29'b0_101010100101_100_1_010101010010;
      patterns[21805] = 29'b0_101010100101_101_0_101010101001;
      patterns[21806] = 29'b0_101010100101_110_0_101010100101;
      patterns[21807] = 29'b0_101010100101_111_0_101010100101;
      patterns[21808] = 29'b0_101010100110_000_0_101010100110;
      patterns[21809] = 29'b0_101010100110_001_0_100110101010;
      patterns[21810] = 29'b0_101010100110_010_1_010101001100;
      patterns[21811] = 29'b0_101010100110_011_0_101010011001;
      patterns[21812] = 29'b0_101010100110_100_0_010101010011;
      patterns[21813] = 29'b0_101010100110_101_1_001010101001;
      patterns[21814] = 29'b0_101010100110_110_0_101010100110;
      patterns[21815] = 29'b0_101010100110_111_0_101010100110;
      patterns[21816] = 29'b0_101010100111_000_0_101010100111;
      patterns[21817] = 29'b0_101010100111_001_0_100111101010;
      patterns[21818] = 29'b0_101010100111_010_1_010101001110;
      patterns[21819] = 29'b0_101010100111_011_0_101010011101;
      patterns[21820] = 29'b0_101010100111_100_1_010101010011;
      patterns[21821] = 29'b0_101010100111_101_1_101010101001;
      patterns[21822] = 29'b0_101010100111_110_0_101010100111;
      patterns[21823] = 29'b0_101010100111_111_0_101010100111;
      patterns[21824] = 29'b0_101010101000_000_0_101010101000;
      patterns[21825] = 29'b0_101010101000_001_0_101000101010;
      patterns[21826] = 29'b0_101010101000_010_1_010101010000;
      patterns[21827] = 29'b0_101010101000_011_0_101010100001;
      patterns[21828] = 29'b0_101010101000_100_0_010101010100;
      patterns[21829] = 29'b0_101010101000_101_0_001010101010;
      patterns[21830] = 29'b0_101010101000_110_0_101010101000;
      patterns[21831] = 29'b0_101010101000_111_0_101010101000;
      patterns[21832] = 29'b0_101010101001_000_0_101010101001;
      patterns[21833] = 29'b0_101010101001_001_0_101001101010;
      patterns[21834] = 29'b0_101010101001_010_1_010101010010;
      patterns[21835] = 29'b0_101010101001_011_0_101010100101;
      patterns[21836] = 29'b0_101010101001_100_1_010101010100;
      patterns[21837] = 29'b0_101010101001_101_0_101010101010;
      patterns[21838] = 29'b0_101010101001_110_0_101010101001;
      patterns[21839] = 29'b0_101010101001_111_0_101010101001;
      patterns[21840] = 29'b0_101010101010_000_0_101010101010;
      patterns[21841] = 29'b0_101010101010_001_0_101010101010;
      patterns[21842] = 29'b0_101010101010_010_1_010101010100;
      patterns[21843] = 29'b0_101010101010_011_0_101010101001;
      patterns[21844] = 29'b0_101010101010_100_0_010101010101;
      patterns[21845] = 29'b0_101010101010_101_1_001010101010;
      patterns[21846] = 29'b0_101010101010_110_0_101010101010;
      patterns[21847] = 29'b0_101010101010_111_0_101010101010;
      patterns[21848] = 29'b0_101010101011_000_0_101010101011;
      patterns[21849] = 29'b0_101010101011_001_0_101011101010;
      patterns[21850] = 29'b0_101010101011_010_1_010101010110;
      patterns[21851] = 29'b0_101010101011_011_0_101010101101;
      patterns[21852] = 29'b0_101010101011_100_1_010101010101;
      patterns[21853] = 29'b0_101010101011_101_1_101010101010;
      patterns[21854] = 29'b0_101010101011_110_0_101010101011;
      patterns[21855] = 29'b0_101010101011_111_0_101010101011;
      patterns[21856] = 29'b0_101010101100_000_0_101010101100;
      patterns[21857] = 29'b0_101010101100_001_0_101100101010;
      patterns[21858] = 29'b0_101010101100_010_1_010101011000;
      patterns[21859] = 29'b0_101010101100_011_0_101010110001;
      patterns[21860] = 29'b0_101010101100_100_0_010101010110;
      patterns[21861] = 29'b0_101010101100_101_0_001010101011;
      patterns[21862] = 29'b0_101010101100_110_0_101010101100;
      patterns[21863] = 29'b0_101010101100_111_0_101010101100;
      patterns[21864] = 29'b0_101010101101_000_0_101010101101;
      patterns[21865] = 29'b0_101010101101_001_0_101101101010;
      patterns[21866] = 29'b0_101010101101_010_1_010101011010;
      patterns[21867] = 29'b0_101010101101_011_0_101010110101;
      patterns[21868] = 29'b0_101010101101_100_1_010101010110;
      patterns[21869] = 29'b0_101010101101_101_0_101010101011;
      patterns[21870] = 29'b0_101010101101_110_0_101010101101;
      patterns[21871] = 29'b0_101010101101_111_0_101010101101;
      patterns[21872] = 29'b0_101010101110_000_0_101010101110;
      patterns[21873] = 29'b0_101010101110_001_0_101110101010;
      patterns[21874] = 29'b0_101010101110_010_1_010101011100;
      patterns[21875] = 29'b0_101010101110_011_0_101010111001;
      patterns[21876] = 29'b0_101010101110_100_0_010101010111;
      patterns[21877] = 29'b0_101010101110_101_1_001010101011;
      patterns[21878] = 29'b0_101010101110_110_0_101010101110;
      patterns[21879] = 29'b0_101010101110_111_0_101010101110;
      patterns[21880] = 29'b0_101010101111_000_0_101010101111;
      patterns[21881] = 29'b0_101010101111_001_0_101111101010;
      patterns[21882] = 29'b0_101010101111_010_1_010101011110;
      patterns[21883] = 29'b0_101010101111_011_0_101010111101;
      patterns[21884] = 29'b0_101010101111_100_1_010101010111;
      patterns[21885] = 29'b0_101010101111_101_1_101010101011;
      patterns[21886] = 29'b0_101010101111_110_0_101010101111;
      patterns[21887] = 29'b0_101010101111_111_0_101010101111;
      patterns[21888] = 29'b0_101010110000_000_0_101010110000;
      patterns[21889] = 29'b0_101010110000_001_0_110000101010;
      patterns[21890] = 29'b0_101010110000_010_1_010101100000;
      patterns[21891] = 29'b0_101010110000_011_0_101011000001;
      patterns[21892] = 29'b0_101010110000_100_0_010101011000;
      patterns[21893] = 29'b0_101010110000_101_0_001010101100;
      patterns[21894] = 29'b0_101010110000_110_0_101010110000;
      patterns[21895] = 29'b0_101010110000_111_0_101010110000;
      patterns[21896] = 29'b0_101010110001_000_0_101010110001;
      patterns[21897] = 29'b0_101010110001_001_0_110001101010;
      patterns[21898] = 29'b0_101010110001_010_1_010101100010;
      patterns[21899] = 29'b0_101010110001_011_0_101011000101;
      patterns[21900] = 29'b0_101010110001_100_1_010101011000;
      patterns[21901] = 29'b0_101010110001_101_0_101010101100;
      patterns[21902] = 29'b0_101010110001_110_0_101010110001;
      patterns[21903] = 29'b0_101010110001_111_0_101010110001;
      patterns[21904] = 29'b0_101010110010_000_0_101010110010;
      patterns[21905] = 29'b0_101010110010_001_0_110010101010;
      patterns[21906] = 29'b0_101010110010_010_1_010101100100;
      patterns[21907] = 29'b0_101010110010_011_0_101011001001;
      patterns[21908] = 29'b0_101010110010_100_0_010101011001;
      patterns[21909] = 29'b0_101010110010_101_1_001010101100;
      patterns[21910] = 29'b0_101010110010_110_0_101010110010;
      patterns[21911] = 29'b0_101010110010_111_0_101010110010;
      patterns[21912] = 29'b0_101010110011_000_0_101010110011;
      patterns[21913] = 29'b0_101010110011_001_0_110011101010;
      patterns[21914] = 29'b0_101010110011_010_1_010101100110;
      patterns[21915] = 29'b0_101010110011_011_0_101011001101;
      patterns[21916] = 29'b0_101010110011_100_1_010101011001;
      patterns[21917] = 29'b0_101010110011_101_1_101010101100;
      patterns[21918] = 29'b0_101010110011_110_0_101010110011;
      patterns[21919] = 29'b0_101010110011_111_0_101010110011;
      patterns[21920] = 29'b0_101010110100_000_0_101010110100;
      patterns[21921] = 29'b0_101010110100_001_0_110100101010;
      patterns[21922] = 29'b0_101010110100_010_1_010101101000;
      patterns[21923] = 29'b0_101010110100_011_0_101011010001;
      patterns[21924] = 29'b0_101010110100_100_0_010101011010;
      patterns[21925] = 29'b0_101010110100_101_0_001010101101;
      patterns[21926] = 29'b0_101010110100_110_0_101010110100;
      patterns[21927] = 29'b0_101010110100_111_0_101010110100;
      patterns[21928] = 29'b0_101010110101_000_0_101010110101;
      patterns[21929] = 29'b0_101010110101_001_0_110101101010;
      patterns[21930] = 29'b0_101010110101_010_1_010101101010;
      patterns[21931] = 29'b0_101010110101_011_0_101011010101;
      patterns[21932] = 29'b0_101010110101_100_1_010101011010;
      patterns[21933] = 29'b0_101010110101_101_0_101010101101;
      patterns[21934] = 29'b0_101010110101_110_0_101010110101;
      patterns[21935] = 29'b0_101010110101_111_0_101010110101;
      patterns[21936] = 29'b0_101010110110_000_0_101010110110;
      patterns[21937] = 29'b0_101010110110_001_0_110110101010;
      patterns[21938] = 29'b0_101010110110_010_1_010101101100;
      patterns[21939] = 29'b0_101010110110_011_0_101011011001;
      patterns[21940] = 29'b0_101010110110_100_0_010101011011;
      patterns[21941] = 29'b0_101010110110_101_1_001010101101;
      patterns[21942] = 29'b0_101010110110_110_0_101010110110;
      patterns[21943] = 29'b0_101010110110_111_0_101010110110;
      patterns[21944] = 29'b0_101010110111_000_0_101010110111;
      patterns[21945] = 29'b0_101010110111_001_0_110111101010;
      patterns[21946] = 29'b0_101010110111_010_1_010101101110;
      patterns[21947] = 29'b0_101010110111_011_0_101011011101;
      patterns[21948] = 29'b0_101010110111_100_1_010101011011;
      patterns[21949] = 29'b0_101010110111_101_1_101010101101;
      patterns[21950] = 29'b0_101010110111_110_0_101010110111;
      patterns[21951] = 29'b0_101010110111_111_0_101010110111;
      patterns[21952] = 29'b0_101010111000_000_0_101010111000;
      patterns[21953] = 29'b0_101010111000_001_0_111000101010;
      patterns[21954] = 29'b0_101010111000_010_1_010101110000;
      patterns[21955] = 29'b0_101010111000_011_0_101011100001;
      patterns[21956] = 29'b0_101010111000_100_0_010101011100;
      patterns[21957] = 29'b0_101010111000_101_0_001010101110;
      patterns[21958] = 29'b0_101010111000_110_0_101010111000;
      patterns[21959] = 29'b0_101010111000_111_0_101010111000;
      patterns[21960] = 29'b0_101010111001_000_0_101010111001;
      patterns[21961] = 29'b0_101010111001_001_0_111001101010;
      patterns[21962] = 29'b0_101010111001_010_1_010101110010;
      patterns[21963] = 29'b0_101010111001_011_0_101011100101;
      patterns[21964] = 29'b0_101010111001_100_1_010101011100;
      patterns[21965] = 29'b0_101010111001_101_0_101010101110;
      patterns[21966] = 29'b0_101010111001_110_0_101010111001;
      patterns[21967] = 29'b0_101010111001_111_0_101010111001;
      patterns[21968] = 29'b0_101010111010_000_0_101010111010;
      patterns[21969] = 29'b0_101010111010_001_0_111010101010;
      patterns[21970] = 29'b0_101010111010_010_1_010101110100;
      patterns[21971] = 29'b0_101010111010_011_0_101011101001;
      patterns[21972] = 29'b0_101010111010_100_0_010101011101;
      patterns[21973] = 29'b0_101010111010_101_1_001010101110;
      patterns[21974] = 29'b0_101010111010_110_0_101010111010;
      patterns[21975] = 29'b0_101010111010_111_0_101010111010;
      patterns[21976] = 29'b0_101010111011_000_0_101010111011;
      patterns[21977] = 29'b0_101010111011_001_0_111011101010;
      patterns[21978] = 29'b0_101010111011_010_1_010101110110;
      patterns[21979] = 29'b0_101010111011_011_0_101011101101;
      patterns[21980] = 29'b0_101010111011_100_1_010101011101;
      patterns[21981] = 29'b0_101010111011_101_1_101010101110;
      patterns[21982] = 29'b0_101010111011_110_0_101010111011;
      patterns[21983] = 29'b0_101010111011_111_0_101010111011;
      patterns[21984] = 29'b0_101010111100_000_0_101010111100;
      patterns[21985] = 29'b0_101010111100_001_0_111100101010;
      patterns[21986] = 29'b0_101010111100_010_1_010101111000;
      patterns[21987] = 29'b0_101010111100_011_0_101011110001;
      patterns[21988] = 29'b0_101010111100_100_0_010101011110;
      patterns[21989] = 29'b0_101010111100_101_0_001010101111;
      patterns[21990] = 29'b0_101010111100_110_0_101010111100;
      patterns[21991] = 29'b0_101010111100_111_0_101010111100;
      patterns[21992] = 29'b0_101010111101_000_0_101010111101;
      patterns[21993] = 29'b0_101010111101_001_0_111101101010;
      patterns[21994] = 29'b0_101010111101_010_1_010101111010;
      patterns[21995] = 29'b0_101010111101_011_0_101011110101;
      patterns[21996] = 29'b0_101010111101_100_1_010101011110;
      patterns[21997] = 29'b0_101010111101_101_0_101010101111;
      patterns[21998] = 29'b0_101010111101_110_0_101010111101;
      patterns[21999] = 29'b0_101010111101_111_0_101010111101;
      patterns[22000] = 29'b0_101010111110_000_0_101010111110;
      patterns[22001] = 29'b0_101010111110_001_0_111110101010;
      patterns[22002] = 29'b0_101010111110_010_1_010101111100;
      patterns[22003] = 29'b0_101010111110_011_0_101011111001;
      patterns[22004] = 29'b0_101010111110_100_0_010101011111;
      patterns[22005] = 29'b0_101010111110_101_1_001010101111;
      patterns[22006] = 29'b0_101010111110_110_0_101010111110;
      patterns[22007] = 29'b0_101010111110_111_0_101010111110;
      patterns[22008] = 29'b0_101010111111_000_0_101010111111;
      patterns[22009] = 29'b0_101010111111_001_0_111111101010;
      patterns[22010] = 29'b0_101010111111_010_1_010101111110;
      patterns[22011] = 29'b0_101010111111_011_0_101011111101;
      patterns[22012] = 29'b0_101010111111_100_1_010101011111;
      patterns[22013] = 29'b0_101010111111_101_1_101010101111;
      patterns[22014] = 29'b0_101010111111_110_0_101010111111;
      patterns[22015] = 29'b0_101010111111_111_0_101010111111;
      patterns[22016] = 29'b0_101011000000_000_0_101011000000;
      patterns[22017] = 29'b0_101011000000_001_0_000000101011;
      patterns[22018] = 29'b0_101011000000_010_1_010110000000;
      patterns[22019] = 29'b0_101011000000_011_0_101100000001;
      patterns[22020] = 29'b0_101011000000_100_0_010101100000;
      patterns[22021] = 29'b0_101011000000_101_0_001010110000;
      patterns[22022] = 29'b0_101011000000_110_0_101011000000;
      patterns[22023] = 29'b0_101011000000_111_0_101011000000;
      patterns[22024] = 29'b0_101011000001_000_0_101011000001;
      patterns[22025] = 29'b0_101011000001_001_0_000001101011;
      patterns[22026] = 29'b0_101011000001_010_1_010110000010;
      patterns[22027] = 29'b0_101011000001_011_0_101100000101;
      patterns[22028] = 29'b0_101011000001_100_1_010101100000;
      patterns[22029] = 29'b0_101011000001_101_0_101010110000;
      patterns[22030] = 29'b0_101011000001_110_0_101011000001;
      patterns[22031] = 29'b0_101011000001_111_0_101011000001;
      patterns[22032] = 29'b0_101011000010_000_0_101011000010;
      patterns[22033] = 29'b0_101011000010_001_0_000010101011;
      patterns[22034] = 29'b0_101011000010_010_1_010110000100;
      patterns[22035] = 29'b0_101011000010_011_0_101100001001;
      patterns[22036] = 29'b0_101011000010_100_0_010101100001;
      patterns[22037] = 29'b0_101011000010_101_1_001010110000;
      patterns[22038] = 29'b0_101011000010_110_0_101011000010;
      patterns[22039] = 29'b0_101011000010_111_0_101011000010;
      patterns[22040] = 29'b0_101011000011_000_0_101011000011;
      patterns[22041] = 29'b0_101011000011_001_0_000011101011;
      patterns[22042] = 29'b0_101011000011_010_1_010110000110;
      patterns[22043] = 29'b0_101011000011_011_0_101100001101;
      patterns[22044] = 29'b0_101011000011_100_1_010101100001;
      patterns[22045] = 29'b0_101011000011_101_1_101010110000;
      patterns[22046] = 29'b0_101011000011_110_0_101011000011;
      patterns[22047] = 29'b0_101011000011_111_0_101011000011;
      patterns[22048] = 29'b0_101011000100_000_0_101011000100;
      patterns[22049] = 29'b0_101011000100_001_0_000100101011;
      patterns[22050] = 29'b0_101011000100_010_1_010110001000;
      patterns[22051] = 29'b0_101011000100_011_0_101100010001;
      patterns[22052] = 29'b0_101011000100_100_0_010101100010;
      patterns[22053] = 29'b0_101011000100_101_0_001010110001;
      patterns[22054] = 29'b0_101011000100_110_0_101011000100;
      patterns[22055] = 29'b0_101011000100_111_0_101011000100;
      patterns[22056] = 29'b0_101011000101_000_0_101011000101;
      patterns[22057] = 29'b0_101011000101_001_0_000101101011;
      patterns[22058] = 29'b0_101011000101_010_1_010110001010;
      patterns[22059] = 29'b0_101011000101_011_0_101100010101;
      patterns[22060] = 29'b0_101011000101_100_1_010101100010;
      patterns[22061] = 29'b0_101011000101_101_0_101010110001;
      patterns[22062] = 29'b0_101011000101_110_0_101011000101;
      patterns[22063] = 29'b0_101011000101_111_0_101011000101;
      patterns[22064] = 29'b0_101011000110_000_0_101011000110;
      patterns[22065] = 29'b0_101011000110_001_0_000110101011;
      patterns[22066] = 29'b0_101011000110_010_1_010110001100;
      patterns[22067] = 29'b0_101011000110_011_0_101100011001;
      patterns[22068] = 29'b0_101011000110_100_0_010101100011;
      patterns[22069] = 29'b0_101011000110_101_1_001010110001;
      patterns[22070] = 29'b0_101011000110_110_0_101011000110;
      patterns[22071] = 29'b0_101011000110_111_0_101011000110;
      patterns[22072] = 29'b0_101011000111_000_0_101011000111;
      patterns[22073] = 29'b0_101011000111_001_0_000111101011;
      patterns[22074] = 29'b0_101011000111_010_1_010110001110;
      patterns[22075] = 29'b0_101011000111_011_0_101100011101;
      patterns[22076] = 29'b0_101011000111_100_1_010101100011;
      patterns[22077] = 29'b0_101011000111_101_1_101010110001;
      patterns[22078] = 29'b0_101011000111_110_0_101011000111;
      patterns[22079] = 29'b0_101011000111_111_0_101011000111;
      patterns[22080] = 29'b0_101011001000_000_0_101011001000;
      patterns[22081] = 29'b0_101011001000_001_0_001000101011;
      patterns[22082] = 29'b0_101011001000_010_1_010110010000;
      patterns[22083] = 29'b0_101011001000_011_0_101100100001;
      patterns[22084] = 29'b0_101011001000_100_0_010101100100;
      patterns[22085] = 29'b0_101011001000_101_0_001010110010;
      patterns[22086] = 29'b0_101011001000_110_0_101011001000;
      patterns[22087] = 29'b0_101011001000_111_0_101011001000;
      patterns[22088] = 29'b0_101011001001_000_0_101011001001;
      patterns[22089] = 29'b0_101011001001_001_0_001001101011;
      patterns[22090] = 29'b0_101011001001_010_1_010110010010;
      patterns[22091] = 29'b0_101011001001_011_0_101100100101;
      patterns[22092] = 29'b0_101011001001_100_1_010101100100;
      patterns[22093] = 29'b0_101011001001_101_0_101010110010;
      patterns[22094] = 29'b0_101011001001_110_0_101011001001;
      patterns[22095] = 29'b0_101011001001_111_0_101011001001;
      patterns[22096] = 29'b0_101011001010_000_0_101011001010;
      patterns[22097] = 29'b0_101011001010_001_0_001010101011;
      patterns[22098] = 29'b0_101011001010_010_1_010110010100;
      patterns[22099] = 29'b0_101011001010_011_0_101100101001;
      patterns[22100] = 29'b0_101011001010_100_0_010101100101;
      patterns[22101] = 29'b0_101011001010_101_1_001010110010;
      patterns[22102] = 29'b0_101011001010_110_0_101011001010;
      patterns[22103] = 29'b0_101011001010_111_0_101011001010;
      patterns[22104] = 29'b0_101011001011_000_0_101011001011;
      patterns[22105] = 29'b0_101011001011_001_0_001011101011;
      patterns[22106] = 29'b0_101011001011_010_1_010110010110;
      patterns[22107] = 29'b0_101011001011_011_0_101100101101;
      patterns[22108] = 29'b0_101011001011_100_1_010101100101;
      patterns[22109] = 29'b0_101011001011_101_1_101010110010;
      patterns[22110] = 29'b0_101011001011_110_0_101011001011;
      patterns[22111] = 29'b0_101011001011_111_0_101011001011;
      patterns[22112] = 29'b0_101011001100_000_0_101011001100;
      patterns[22113] = 29'b0_101011001100_001_0_001100101011;
      patterns[22114] = 29'b0_101011001100_010_1_010110011000;
      patterns[22115] = 29'b0_101011001100_011_0_101100110001;
      patterns[22116] = 29'b0_101011001100_100_0_010101100110;
      patterns[22117] = 29'b0_101011001100_101_0_001010110011;
      patterns[22118] = 29'b0_101011001100_110_0_101011001100;
      patterns[22119] = 29'b0_101011001100_111_0_101011001100;
      patterns[22120] = 29'b0_101011001101_000_0_101011001101;
      patterns[22121] = 29'b0_101011001101_001_0_001101101011;
      patterns[22122] = 29'b0_101011001101_010_1_010110011010;
      patterns[22123] = 29'b0_101011001101_011_0_101100110101;
      patterns[22124] = 29'b0_101011001101_100_1_010101100110;
      patterns[22125] = 29'b0_101011001101_101_0_101010110011;
      patterns[22126] = 29'b0_101011001101_110_0_101011001101;
      patterns[22127] = 29'b0_101011001101_111_0_101011001101;
      patterns[22128] = 29'b0_101011001110_000_0_101011001110;
      patterns[22129] = 29'b0_101011001110_001_0_001110101011;
      patterns[22130] = 29'b0_101011001110_010_1_010110011100;
      patterns[22131] = 29'b0_101011001110_011_0_101100111001;
      patterns[22132] = 29'b0_101011001110_100_0_010101100111;
      patterns[22133] = 29'b0_101011001110_101_1_001010110011;
      patterns[22134] = 29'b0_101011001110_110_0_101011001110;
      patterns[22135] = 29'b0_101011001110_111_0_101011001110;
      patterns[22136] = 29'b0_101011001111_000_0_101011001111;
      patterns[22137] = 29'b0_101011001111_001_0_001111101011;
      patterns[22138] = 29'b0_101011001111_010_1_010110011110;
      patterns[22139] = 29'b0_101011001111_011_0_101100111101;
      patterns[22140] = 29'b0_101011001111_100_1_010101100111;
      patterns[22141] = 29'b0_101011001111_101_1_101010110011;
      patterns[22142] = 29'b0_101011001111_110_0_101011001111;
      patterns[22143] = 29'b0_101011001111_111_0_101011001111;
      patterns[22144] = 29'b0_101011010000_000_0_101011010000;
      patterns[22145] = 29'b0_101011010000_001_0_010000101011;
      patterns[22146] = 29'b0_101011010000_010_1_010110100000;
      patterns[22147] = 29'b0_101011010000_011_0_101101000001;
      patterns[22148] = 29'b0_101011010000_100_0_010101101000;
      patterns[22149] = 29'b0_101011010000_101_0_001010110100;
      patterns[22150] = 29'b0_101011010000_110_0_101011010000;
      patterns[22151] = 29'b0_101011010000_111_0_101011010000;
      patterns[22152] = 29'b0_101011010001_000_0_101011010001;
      patterns[22153] = 29'b0_101011010001_001_0_010001101011;
      patterns[22154] = 29'b0_101011010001_010_1_010110100010;
      patterns[22155] = 29'b0_101011010001_011_0_101101000101;
      patterns[22156] = 29'b0_101011010001_100_1_010101101000;
      patterns[22157] = 29'b0_101011010001_101_0_101010110100;
      patterns[22158] = 29'b0_101011010001_110_0_101011010001;
      patterns[22159] = 29'b0_101011010001_111_0_101011010001;
      patterns[22160] = 29'b0_101011010010_000_0_101011010010;
      patterns[22161] = 29'b0_101011010010_001_0_010010101011;
      patterns[22162] = 29'b0_101011010010_010_1_010110100100;
      patterns[22163] = 29'b0_101011010010_011_0_101101001001;
      patterns[22164] = 29'b0_101011010010_100_0_010101101001;
      patterns[22165] = 29'b0_101011010010_101_1_001010110100;
      patterns[22166] = 29'b0_101011010010_110_0_101011010010;
      patterns[22167] = 29'b0_101011010010_111_0_101011010010;
      patterns[22168] = 29'b0_101011010011_000_0_101011010011;
      patterns[22169] = 29'b0_101011010011_001_0_010011101011;
      patterns[22170] = 29'b0_101011010011_010_1_010110100110;
      patterns[22171] = 29'b0_101011010011_011_0_101101001101;
      patterns[22172] = 29'b0_101011010011_100_1_010101101001;
      patterns[22173] = 29'b0_101011010011_101_1_101010110100;
      patterns[22174] = 29'b0_101011010011_110_0_101011010011;
      patterns[22175] = 29'b0_101011010011_111_0_101011010011;
      patterns[22176] = 29'b0_101011010100_000_0_101011010100;
      patterns[22177] = 29'b0_101011010100_001_0_010100101011;
      patterns[22178] = 29'b0_101011010100_010_1_010110101000;
      patterns[22179] = 29'b0_101011010100_011_0_101101010001;
      patterns[22180] = 29'b0_101011010100_100_0_010101101010;
      patterns[22181] = 29'b0_101011010100_101_0_001010110101;
      patterns[22182] = 29'b0_101011010100_110_0_101011010100;
      patterns[22183] = 29'b0_101011010100_111_0_101011010100;
      patterns[22184] = 29'b0_101011010101_000_0_101011010101;
      patterns[22185] = 29'b0_101011010101_001_0_010101101011;
      patterns[22186] = 29'b0_101011010101_010_1_010110101010;
      patterns[22187] = 29'b0_101011010101_011_0_101101010101;
      patterns[22188] = 29'b0_101011010101_100_1_010101101010;
      patterns[22189] = 29'b0_101011010101_101_0_101010110101;
      patterns[22190] = 29'b0_101011010101_110_0_101011010101;
      patterns[22191] = 29'b0_101011010101_111_0_101011010101;
      patterns[22192] = 29'b0_101011010110_000_0_101011010110;
      patterns[22193] = 29'b0_101011010110_001_0_010110101011;
      patterns[22194] = 29'b0_101011010110_010_1_010110101100;
      patterns[22195] = 29'b0_101011010110_011_0_101101011001;
      patterns[22196] = 29'b0_101011010110_100_0_010101101011;
      patterns[22197] = 29'b0_101011010110_101_1_001010110101;
      patterns[22198] = 29'b0_101011010110_110_0_101011010110;
      patterns[22199] = 29'b0_101011010110_111_0_101011010110;
      patterns[22200] = 29'b0_101011010111_000_0_101011010111;
      patterns[22201] = 29'b0_101011010111_001_0_010111101011;
      patterns[22202] = 29'b0_101011010111_010_1_010110101110;
      patterns[22203] = 29'b0_101011010111_011_0_101101011101;
      patterns[22204] = 29'b0_101011010111_100_1_010101101011;
      patterns[22205] = 29'b0_101011010111_101_1_101010110101;
      patterns[22206] = 29'b0_101011010111_110_0_101011010111;
      patterns[22207] = 29'b0_101011010111_111_0_101011010111;
      patterns[22208] = 29'b0_101011011000_000_0_101011011000;
      patterns[22209] = 29'b0_101011011000_001_0_011000101011;
      patterns[22210] = 29'b0_101011011000_010_1_010110110000;
      patterns[22211] = 29'b0_101011011000_011_0_101101100001;
      patterns[22212] = 29'b0_101011011000_100_0_010101101100;
      patterns[22213] = 29'b0_101011011000_101_0_001010110110;
      patterns[22214] = 29'b0_101011011000_110_0_101011011000;
      patterns[22215] = 29'b0_101011011000_111_0_101011011000;
      patterns[22216] = 29'b0_101011011001_000_0_101011011001;
      patterns[22217] = 29'b0_101011011001_001_0_011001101011;
      patterns[22218] = 29'b0_101011011001_010_1_010110110010;
      patterns[22219] = 29'b0_101011011001_011_0_101101100101;
      patterns[22220] = 29'b0_101011011001_100_1_010101101100;
      patterns[22221] = 29'b0_101011011001_101_0_101010110110;
      patterns[22222] = 29'b0_101011011001_110_0_101011011001;
      patterns[22223] = 29'b0_101011011001_111_0_101011011001;
      patterns[22224] = 29'b0_101011011010_000_0_101011011010;
      patterns[22225] = 29'b0_101011011010_001_0_011010101011;
      patterns[22226] = 29'b0_101011011010_010_1_010110110100;
      patterns[22227] = 29'b0_101011011010_011_0_101101101001;
      patterns[22228] = 29'b0_101011011010_100_0_010101101101;
      patterns[22229] = 29'b0_101011011010_101_1_001010110110;
      patterns[22230] = 29'b0_101011011010_110_0_101011011010;
      patterns[22231] = 29'b0_101011011010_111_0_101011011010;
      patterns[22232] = 29'b0_101011011011_000_0_101011011011;
      patterns[22233] = 29'b0_101011011011_001_0_011011101011;
      patterns[22234] = 29'b0_101011011011_010_1_010110110110;
      patterns[22235] = 29'b0_101011011011_011_0_101101101101;
      patterns[22236] = 29'b0_101011011011_100_1_010101101101;
      patterns[22237] = 29'b0_101011011011_101_1_101010110110;
      patterns[22238] = 29'b0_101011011011_110_0_101011011011;
      patterns[22239] = 29'b0_101011011011_111_0_101011011011;
      patterns[22240] = 29'b0_101011011100_000_0_101011011100;
      patterns[22241] = 29'b0_101011011100_001_0_011100101011;
      patterns[22242] = 29'b0_101011011100_010_1_010110111000;
      patterns[22243] = 29'b0_101011011100_011_0_101101110001;
      patterns[22244] = 29'b0_101011011100_100_0_010101101110;
      patterns[22245] = 29'b0_101011011100_101_0_001010110111;
      patterns[22246] = 29'b0_101011011100_110_0_101011011100;
      patterns[22247] = 29'b0_101011011100_111_0_101011011100;
      patterns[22248] = 29'b0_101011011101_000_0_101011011101;
      patterns[22249] = 29'b0_101011011101_001_0_011101101011;
      patterns[22250] = 29'b0_101011011101_010_1_010110111010;
      patterns[22251] = 29'b0_101011011101_011_0_101101110101;
      patterns[22252] = 29'b0_101011011101_100_1_010101101110;
      patterns[22253] = 29'b0_101011011101_101_0_101010110111;
      patterns[22254] = 29'b0_101011011101_110_0_101011011101;
      patterns[22255] = 29'b0_101011011101_111_0_101011011101;
      patterns[22256] = 29'b0_101011011110_000_0_101011011110;
      patterns[22257] = 29'b0_101011011110_001_0_011110101011;
      patterns[22258] = 29'b0_101011011110_010_1_010110111100;
      patterns[22259] = 29'b0_101011011110_011_0_101101111001;
      patterns[22260] = 29'b0_101011011110_100_0_010101101111;
      patterns[22261] = 29'b0_101011011110_101_1_001010110111;
      patterns[22262] = 29'b0_101011011110_110_0_101011011110;
      patterns[22263] = 29'b0_101011011110_111_0_101011011110;
      patterns[22264] = 29'b0_101011011111_000_0_101011011111;
      patterns[22265] = 29'b0_101011011111_001_0_011111101011;
      patterns[22266] = 29'b0_101011011111_010_1_010110111110;
      patterns[22267] = 29'b0_101011011111_011_0_101101111101;
      patterns[22268] = 29'b0_101011011111_100_1_010101101111;
      patterns[22269] = 29'b0_101011011111_101_1_101010110111;
      patterns[22270] = 29'b0_101011011111_110_0_101011011111;
      patterns[22271] = 29'b0_101011011111_111_0_101011011111;
      patterns[22272] = 29'b0_101011100000_000_0_101011100000;
      patterns[22273] = 29'b0_101011100000_001_0_100000101011;
      patterns[22274] = 29'b0_101011100000_010_1_010111000000;
      patterns[22275] = 29'b0_101011100000_011_0_101110000001;
      patterns[22276] = 29'b0_101011100000_100_0_010101110000;
      patterns[22277] = 29'b0_101011100000_101_0_001010111000;
      patterns[22278] = 29'b0_101011100000_110_0_101011100000;
      patterns[22279] = 29'b0_101011100000_111_0_101011100000;
      patterns[22280] = 29'b0_101011100001_000_0_101011100001;
      patterns[22281] = 29'b0_101011100001_001_0_100001101011;
      patterns[22282] = 29'b0_101011100001_010_1_010111000010;
      patterns[22283] = 29'b0_101011100001_011_0_101110000101;
      patterns[22284] = 29'b0_101011100001_100_1_010101110000;
      patterns[22285] = 29'b0_101011100001_101_0_101010111000;
      patterns[22286] = 29'b0_101011100001_110_0_101011100001;
      patterns[22287] = 29'b0_101011100001_111_0_101011100001;
      patterns[22288] = 29'b0_101011100010_000_0_101011100010;
      patterns[22289] = 29'b0_101011100010_001_0_100010101011;
      patterns[22290] = 29'b0_101011100010_010_1_010111000100;
      patterns[22291] = 29'b0_101011100010_011_0_101110001001;
      patterns[22292] = 29'b0_101011100010_100_0_010101110001;
      patterns[22293] = 29'b0_101011100010_101_1_001010111000;
      patterns[22294] = 29'b0_101011100010_110_0_101011100010;
      patterns[22295] = 29'b0_101011100010_111_0_101011100010;
      patterns[22296] = 29'b0_101011100011_000_0_101011100011;
      patterns[22297] = 29'b0_101011100011_001_0_100011101011;
      patterns[22298] = 29'b0_101011100011_010_1_010111000110;
      patterns[22299] = 29'b0_101011100011_011_0_101110001101;
      patterns[22300] = 29'b0_101011100011_100_1_010101110001;
      patterns[22301] = 29'b0_101011100011_101_1_101010111000;
      patterns[22302] = 29'b0_101011100011_110_0_101011100011;
      patterns[22303] = 29'b0_101011100011_111_0_101011100011;
      patterns[22304] = 29'b0_101011100100_000_0_101011100100;
      patterns[22305] = 29'b0_101011100100_001_0_100100101011;
      patterns[22306] = 29'b0_101011100100_010_1_010111001000;
      patterns[22307] = 29'b0_101011100100_011_0_101110010001;
      patterns[22308] = 29'b0_101011100100_100_0_010101110010;
      patterns[22309] = 29'b0_101011100100_101_0_001010111001;
      patterns[22310] = 29'b0_101011100100_110_0_101011100100;
      patterns[22311] = 29'b0_101011100100_111_0_101011100100;
      patterns[22312] = 29'b0_101011100101_000_0_101011100101;
      patterns[22313] = 29'b0_101011100101_001_0_100101101011;
      patterns[22314] = 29'b0_101011100101_010_1_010111001010;
      patterns[22315] = 29'b0_101011100101_011_0_101110010101;
      patterns[22316] = 29'b0_101011100101_100_1_010101110010;
      patterns[22317] = 29'b0_101011100101_101_0_101010111001;
      patterns[22318] = 29'b0_101011100101_110_0_101011100101;
      patterns[22319] = 29'b0_101011100101_111_0_101011100101;
      patterns[22320] = 29'b0_101011100110_000_0_101011100110;
      patterns[22321] = 29'b0_101011100110_001_0_100110101011;
      patterns[22322] = 29'b0_101011100110_010_1_010111001100;
      patterns[22323] = 29'b0_101011100110_011_0_101110011001;
      patterns[22324] = 29'b0_101011100110_100_0_010101110011;
      patterns[22325] = 29'b0_101011100110_101_1_001010111001;
      patterns[22326] = 29'b0_101011100110_110_0_101011100110;
      patterns[22327] = 29'b0_101011100110_111_0_101011100110;
      patterns[22328] = 29'b0_101011100111_000_0_101011100111;
      patterns[22329] = 29'b0_101011100111_001_0_100111101011;
      patterns[22330] = 29'b0_101011100111_010_1_010111001110;
      patterns[22331] = 29'b0_101011100111_011_0_101110011101;
      patterns[22332] = 29'b0_101011100111_100_1_010101110011;
      patterns[22333] = 29'b0_101011100111_101_1_101010111001;
      patterns[22334] = 29'b0_101011100111_110_0_101011100111;
      patterns[22335] = 29'b0_101011100111_111_0_101011100111;
      patterns[22336] = 29'b0_101011101000_000_0_101011101000;
      patterns[22337] = 29'b0_101011101000_001_0_101000101011;
      patterns[22338] = 29'b0_101011101000_010_1_010111010000;
      patterns[22339] = 29'b0_101011101000_011_0_101110100001;
      patterns[22340] = 29'b0_101011101000_100_0_010101110100;
      patterns[22341] = 29'b0_101011101000_101_0_001010111010;
      patterns[22342] = 29'b0_101011101000_110_0_101011101000;
      patterns[22343] = 29'b0_101011101000_111_0_101011101000;
      patterns[22344] = 29'b0_101011101001_000_0_101011101001;
      patterns[22345] = 29'b0_101011101001_001_0_101001101011;
      patterns[22346] = 29'b0_101011101001_010_1_010111010010;
      patterns[22347] = 29'b0_101011101001_011_0_101110100101;
      patterns[22348] = 29'b0_101011101001_100_1_010101110100;
      patterns[22349] = 29'b0_101011101001_101_0_101010111010;
      patterns[22350] = 29'b0_101011101001_110_0_101011101001;
      patterns[22351] = 29'b0_101011101001_111_0_101011101001;
      patterns[22352] = 29'b0_101011101010_000_0_101011101010;
      patterns[22353] = 29'b0_101011101010_001_0_101010101011;
      patterns[22354] = 29'b0_101011101010_010_1_010111010100;
      patterns[22355] = 29'b0_101011101010_011_0_101110101001;
      patterns[22356] = 29'b0_101011101010_100_0_010101110101;
      patterns[22357] = 29'b0_101011101010_101_1_001010111010;
      patterns[22358] = 29'b0_101011101010_110_0_101011101010;
      patterns[22359] = 29'b0_101011101010_111_0_101011101010;
      patterns[22360] = 29'b0_101011101011_000_0_101011101011;
      patterns[22361] = 29'b0_101011101011_001_0_101011101011;
      patterns[22362] = 29'b0_101011101011_010_1_010111010110;
      patterns[22363] = 29'b0_101011101011_011_0_101110101101;
      patterns[22364] = 29'b0_101011101011_100_1_010101110101;
      patterns[22365] = 29'b0_101011101011_101_1_101010111010;
      patterns[22366] = 29'b0_101011101011_110_0_101011101011;
      patterns[22367] = 29'b0_101011101011_111_0_101011101011;
      patterns[22368] = 29'b0_101011101100_000_0_101011101100;
      patterns[22369] = 29'b0_101011101100_001_0_101100101011;
      patterns[22370] = 29'b0_101011101100_010_1_010111011000;
      patterns[22371] = 29'b0_101011101100_011_0_101110110001;
      patterns[22372] = 29'b0_101011101100_100_0_010101110110;
      patterns[22373] = 29'b0_101011101100_101_0_001010111011;
      patterns[22374] = 29'b0_101011101100_110_0_101011101100;
      patterns[22375] = 29'b0_101011101100_111_0_101011101100;
      patterns[22376] = 29'b0_101011101101_000_0_101011101101;
      patterns[22377] = 29'b0_101011101101_001_0_101101101011;
      patterns[22378] = 29'b0_101011101101_010_1_010111011010;
      patterns[22379] = 29'b0_101011101101_011_0_101110110101;
      patterns[22380] = 29'b0_101011101101_100_1_010101110110;
      patterns[22381] = 29'b0_101011101101_101_0_101010111011;
      patterns[22382] = 29'b0_101011101101_110_0_101011101101;
      patterns[22383] = 29'b0_101011101101_111_0_101011101101;
      patterns[22384] = 29'b0_101011101110_000_0_101011101110;
      patterns[22385] = 29'b0_101011101110_001_0_101110101011;
      patterns[22386] = 29'b0_101011101110_010_1_010111011100;
      patterns[22387] = 29'b0_101011101110_011_0_101110111001;
      patterns[22388] = 29'b0_101011101110_100_0_010101110111;
      patterns[22389] = 29'b0_101011101110_101_1_001010111011;
      patterns[22390] = 29'b0_101011101110_110_0_101011101110;
      patterns[22391] = 29'b0_101011101110_111_0_101011101110;
      patterns[22392] = 29'b0_101011101111_000_0_101011101111;
      patterns[22393] = 29'b0_101011101111_001_0_101111101011;
      patterns[22394] = 29'b0_101011101111_010_1_010111011110;
      patterns[22395] = 29'b0_101011101111_011_0_101110111101;
      patterns[22396] = 29'b0_101011101111_100_1_010101110111;
      patterns[22397] = 29'b0_101011101111_101_1_101010111011;
      patterns[22398] = 29'b0_101011101111_110_0_101011101111;
      patterns[22399] = 29'b0_101011101111_111_0_101011101111;
      patterns[22400] = 29'b0_101011110000_000_0_101011110000;
      patterns[22401] = 29'b0_101011110000_001_0_110000101011;
      patterns[22402] = 29'b0_101011110000_010_1_010111100000;
      patterns[22403] = 29'b0_101011110000_011_0_101111000001;
      patterns[22404] = 29'b0_101011110000_100_0_010101111000;
      patterns[22405] = 29'b0_101011110000_101_0_001010111100;
      patterns[22406] = 29'b0_101011110000_110_0_101011110000;
      patterns[22407] = 29'b0_101011110000_111_0_101011110000;
      patterns[22408] = 29'b0_101011110001_000_0_101011110001;
      patterns[22409] = 29'b0_101011110001_001_0_110001101011;
      patterns[22410] = 29'b0_101011110001_010_1_010111100010;
      patterns[22411] = 29'b0_101011110001_011_0_101111000101;
      patterns[22412] = 29'b0_101011110001_100_1_010101111000;
      patterns[22413] = 29'b0_101011110001_101_0_101010111100;
      patterns[22414] = 29'b0_101011110001_110_0_101011110001;
      patterns[22415] = 29'b0_101011110001_111_0_101011110001;
      patterns[22416] = 29'b0_101011110010_000_0_101011110010;
      patterns[22417] = 29'b0_101011110010_001_0_110010101011;
      patterns[22418] = 29'b0_101011110010_010_1_010111100100;
      patterns[22419] = 29'b0_101011110010_011_0_101111001001;
      patterns[22420] = 29'b0_101011110010_100_0_010101111001;
      patterns[22421] = 29'b0_101011110010_101_1_001010111100;
      patterns[22422] = 29'b0_101011110010_110_0_101011110010;
      patterns[22423] = 29'b0_101011110010_111_0_101011110010;
      patterns[22424] = 29'b0_101011110011_000_0_101011110011;
      patterns[22425] = 29'b0_101011110011_001_0_110011101011;
      patterns[22426] = 29'b0_101011110011_010_1_010111100110;
      patterns[22427] = 29'b0_101011110011_011_0_101111001101;
      patterns[22428] = 29'b0_101011110011_100_1_010101111001;
      patterns[22429] = 29'b0_101011110011_101_1_101010111100;
      patterns[22430] = 29'b0_101011110011_110_0_101011110011;
      patterns[22431] = 29'b0_101011110011_111_0_101011110011;
      patterns[22432] = 29'b0_101011110100_000_0_101011110100;
      patterns[22433] = 29'b0_101011110100_001_0_110100101011;
      patterns[22434] = 29'b0_101011110100_010_1_010111101000;
      patterns[22435] = 29'b0_101011110100_011_0_101111010001;
      patterns[22436] = 29'b0_101011110100_100_0_010101111010;
      patterns[22437] = 29'b0_101011110100_101_0_001010111101;
      patterns[22438] = 29'b0_101011110100_110_0_101011110100;
      patterns[22439] = 29'b0_101011110100_111_0_101011110100;
      patterns[22440] = 29'b0_101011110101_000_0_101011110101;
      patterns[22441] = 29'b0_101011110101_001_0_110101101011;
      patterns[22442] = 29'b0_101011110101_010_1_010111101010;
      patterns[22443] = 29'b0_101011110101_011_0_101111010101;
      patterns[22444] = 29'b0_101011110101_100_1_010101111010;
      patterns[22445] = 29'b0_101011110101_101_0_101010111101;
      patterns[22446] = 29'b0_101011110101_110_0_101011110101;
      patterns[22447] = 29'b0_101011110101_111_0_101011110101;
      patterns[22448] = 29'b0_101011110110_000_0_101011110110;
      patterns[22449] = 29'b0_101011110110_001_0_110110101011;
      patterns[22450] = 29'b0_101011110110_010_1_010111101100;
      patterns[22451] = 29'b0_101011110110_011_0_101111011001;
      patterns[22452] = 29'b0_101011110110_100_0_010101111011;
      patterns[22453] = 29'b0_101011110110_101_1_001010111101;
      patterns[22454] = 29'b0_101011110110_110_0_101011110110;
      patterns[22455] = 29'b0_101011110110_111_0_101011110110;
      patterns[22456] = 29'b0_101011110111_000_0_101011110111;
      patterns[22457] = 29'b0_101011110111_001_0_110111101011;
      patterns[22458] = 29'b0_101011110111_010_1_010111101110;
      patterns[22459] = 29'b0_101011110111_011_0_101111011101;
      patterns[22460] = 29'b0_101011110111_100_1_010101111011;
      patterns[22461] = 29'b0_101011110111_101_1_101010111101;
      patterns[22462] = 29'b0_101011110111_110_0_101011110111;
      patterns[22463] = 29'b0_101011110111_111_0_101011110111;
      patterns[22464] = 29'b0_101011111000_000_0_101011111000;
      patterns[22465] = 29'b0_101011111000_001_0_111000101011;
      patterns[22466] = 29'b0_101011111000_010_1_010111110000;
      patterns[22467] = 29'b0_101011111000_011_0_101111100001;
      patterns[22468] = 29'b0_101011111000_100_0_010101111100;
      patterns[22469] = 29'b0_101011111000_101_0_001010111110;
      patterns[22470] = 29'b0_101011111000_110_0_101011111000;
      patterns[22471] = 29'b0_101011111000_111_0_101011111000;
      patterns[22472] = 29'b0_101011111001_000_0_101011111001;
      patterns[22473] = 29'b0_101011111001_001_0_111001101011;
      patterns[22474] = 29'b0_101011111001_010_1_010111110010;
      patterns[22475] = 29'b0_101011111001_011_0_101111100101;
      patterns[22476] = 29'b0_101011111001_100_1_010101111100;
      patterns[22477] = 29'b0_101011111001_101_0_101010111110;
      patterns[22478] = 29'b0_101011111001_110_0_101011111001;
      patterns[22479] = 29'b0_101011111001_111_0_101011111001;
      patterns[22480] = 29'b0_101011111010_000_0_101011111010;
      patterns[22481] = 29'b0_101011111010_001_0_111010101011;
      patterns[22482] = 29'b0_101011111010_010_1_010111110100;
      patterns[22483] = 29'b0_101011111010_011_0_101111101001;
      patterns[22484] = 29'b0_101011111010_100_0_010101111101;
      patterns[22485] = 29'b0_101011111010_101_1_001010111110;
      patterns[22486] = 29'b0_101011111010_110_0_101011111010;
      patterns[22487] = 29'b0_101011111010_111_0_101011111010;
      patterns[22488] = 29'b0_101011111011_000_0_101011111011;
      patterns[22489] = 29'b0_101011111011_001_0_111011101011;
      patterns[22490] = 29'b0_101011111011_010_1_010111110110;
      patterns[22491] = 29'b0_101011111011_011_0_101111101101;
      patterns[22492] = 29'b0_101011111011_100_1_010101111101;
      patterns[22493] = 29'b0_101011111011_101_1_101010111110;
      patterns[22494] = 29'b0_101011111011_110_0_101011111011;
      patterns[22495] = 29'b0_101011111011_111_0_101011111011;
      patterns[22496] = 29'b0_101011111100_000_0_101011111100;
      patterns[22497] = 29'b0_101011111100_001_0_111100101011;
      patterns[22498] = 29'b0_101011111100_010_1_010111111000;
      patterns[22499] = 29'b0_101011111100_011_0_101111110001;
      patterns[22500] = 29'b0_101011111100_100_0_010101111110;
      patterns[22501] = 29'b0_101011111100_101_0_001010111111;
      patterns[22502] = 29'b0_101011111100_110_0_101011111100;
      patterns[22503] = 29'b0_101011111100_111_0_101011111100;
      patterns[22504] = 29'b0_101011111101_000_0_101011111101;
      patterns[22505] = 29'b0_101011111101_001_0_111101101011;
      patterns[22506] = 29'b0_101011111101_010_1_010111111010;
      patterns[22507] = 29'b0_101011111101_011_0_101111110101;
      patterns[22508] = 29'b0_101011111101_100_1_010101111110;
      patterns[22509] = 29'b0_101011111101_101_0_101010111111;
      patterns[22510] = 29'b0_101011111101_110_0_101011111101;
      patterns[22511] = 29'b0_101011111101_111_0_101011111101;
      patterns[22512] = 29'b0_101011111110_000_0_101011111110;
      patterns[22513] = 29'b0_101011111110_001_0_111110101011;
      patterns[22514] = 29'b0_101011111110_010_1_010111111100;
      patterns[22515] = 29'b0_101011111110_011_0_101111111001;
      patterns[22516] = 29'b0_101011111110_100_0_010101111111;
      patterns[22517] = 29'b0_101011111110_101_1_001010111111;
      patterns[22518] = 29'b0_101011111110_110_0_101011111110;
      patterns[22519] = 29'b0_101011111110_111_0_101011111110;
      patterns[22520] = 29'b0_101011111111_000_0_101011111111;
      patterns[22521] = 29'b0_101011111111_001_0_111111101011;
      patterns[22522] = 29'b0_101011111111_010_1_010111111110;
      patterns[22523] = 29'b0_101011111111_011_0_101111111101;
      patterns[22524] = 29'b0_101011111111_100_1_010101111111;
      patterns[22525] = 29'b0_101011111111_101_1_101010111111;
      patterns[22526] = 29'b0_101011111111_110_0_101011111111;
      patterns[22527] = 29'b0_101011111111_111_0_101011111111;
      patterns[22528] = 29'b0_101100000000_000_0_101100000000;
      patterns[22529] = 29'b0_101100000000_001_0_000000101100;
      patterns[22530] = 29'b0_101100000000_010_1_011000000000;
      patterns[22531] = 29'b0_101100000000_011_0_110000000001;
      patterns[22532] = 29'b0_101100000000_100_0_010110000000;
      patterns[22533] = 29'b0_101100000000_101_0_001011000000;
      patterns[22534] = 29'b0_101100000000_110_0_101100000000;
      patterns[22535] = 29'b0_101100000000_111_0_101100000000;
      patterns[22536] = 29'b0_101100000001_000_0_101100000001;
      patterns[22537] = 29'b0_101100000001_001_0_000001101100;
      patterns[22538] = 29'b0_101100000001_010_1_011000000010;
      patterns[22539] = 29'b0_101100000001_011_0_110000000101;
      patterns[22540] = 29'b0_101100000001_100_1_010110000000;
      patterns[22541] = 29'b0_101100000001_101_0_101011000000;
      patterns[22542] = 29'b0_101100000001_110_0_101100000001;
      patterns[22543] = 29'b0_101100000001_111_0_101100000001;
      patterns[22544] = 29'b0_101100000010_000_0_101100000010;
      patterns[22545] = 29'b0_101100000010_001_0_000010101100;
      patterns[22546] = 29'b0_101100000010_010_1_011000000100;
      patterns[22547] = 29'b0_101100000010_011_0_110000001001;
      patterns[22548] = 29'b0_101100000010_100_0_010110000001;
      patterns[22549] = 29'b0_101100000010_101_1_001011000000;
      patterns[22550] = 29'b0_101100000010_110_0_101100000010;
      patterns[22551] = 29'b0_101100000010_111_0_101100000010;
      patterns[22552] = 29'b0_101100000011_000_0_101100000011;
      patterns[22553] = 29'b0_101100000011_001_0_000011101100;
      patterns[22554] = 29'b0_101100000011_010_1_011000000110;
      patterns[22555] = 29'b0_101100000011_011_0_110000001101;
      patterns[22556] = 29'b0_101100000011_100_1_010110000001;
      patterns[22557] = 29'b0_101100000011_101_1_101011000000;
      patterns[22558] = 29'b0_101100000011_110_0_101100000011;
      patterns[22559] = 29'b0_101100000011_111_0_101100000011;
      patterns[22560] = 29'b0_101100000100_000_0_101100000100;
      patterns[22561] = 29'b0_101100000100_001_0_000100101100;
      patterns[22562] = 29'b0_101100000100_010_1_011000001000;
      patterns[22563] = 29'b0_101100000100_011_0_110000010001;
      patterns[22564] = 29'b0_101100000100_100_0_010110000010;
      patterns[22565] = 29'b0_101100000100_101_0_001011000001;
      patterns[22566] = 29'b0_101100000100_110_0_101100000100;
      patterns[22567] = 29'b0_101100000100_111_0_101100000100;
      patterns[22568] = 29'b0_101100000101_000_0_101100000101;
      patterns[22569] = 29'b0_101100000101_001_0_000101101100;
      patterns[22570] = 29'b0_101100000101_010_1_011000001010;
      patterns[22571] = 29'b0_101100000101_011_0_110000010101;
      patterns[22572] = 29'b0_101100000101_100_1_010110000010;
      patterns[22573] = 29'b0_101100000101_101_0_101011000001;
      patterns[22574] = 29'b0_101100000101_110_0_101100000101;
      patterns[22575] = 29'b0_101100000101_111_0_101100000101;
      patterns[22576] = 29'b0_101100000110_000_0_101100000110;
      patterns[22577] = 29'b0_101100000110_001_0_000110101100;
      patterns[22578] = 29'b0_101100000110_010_1_011000001100;
      patterns[22579] = 29'b0_101100000110_011_0_110000011001;
      patterns[22580] = 29'b0_101100000110_100_0_010110000011;
      patterns[22581] = 29'b0_101100000110_101_1_001011000001;
      patterns[22582] = 29'b0_101100000110_110_0_101100000110;
      patterns[22583] = 29'b0_101100000110_111_0_101100000110;
      patterns[22584] = 29'b0_101100000111_000_0_101100000111;
      patterns[22585] = 29'b0_101100000111_001_0_000111101100;
      patterns[22586] = 29'b0_101100000111_010_1_011000001110;
      patterns[22587] = 29'b0_101100000111_011_0_110000011101;
      patterns[22588] = 29'b0_101100000111_100_1_010110000011;
      patterns[22589] = 29'b0_101100000111_101_1_101011000001;
      patterns[22590] = 29'b0_101100000111_110_0_101100000111;
      patterns[22591] = 29'b0_101100000111_111_0_101100000111;
      patterns[22592] = 29'b0_101100001000_000_0_101100001000;
      patterns[22593] = 29'b0_101100001000_001_0_001000101100;
      patterns[22594] = 29'b0_101100001000_010_1_011000010000;
      patterns[22595] = 29'b0_101100001000_011_0_110000100001;
      patterns[22596] = 29'b0_101100001000_100_0_010110000100;
      patterns[22597] = 29'b0_101100001000_101_0_001011000010;
      patterns[22598] = 29'b0_101100001000_110_0_101100001000;
      patterns[22599] = 29'b0_101100001000_111_0_101100001000;
      patterns[22600] = 29'b0_101100001001_000_0_101100001001;
      patterns[22601] = 29'b0_101100001001_001_0_001001101100;
      patterns[22602] = 29'b0_101100001001_010_1_011000010010;
      patterns[22603] = 29'b0_101100001001_011_0_110000100101;
      patterns[22604] = 29'b0_101100001001_100_1_010110000100;
      patterns[22605] = 29'b0_101100001001_101_0_101011000010;
      patterns[22606] = 29'b0_101100001001_110_0_101100001001;
      patterns[22607] = 29'b0_101100001001_111_0_101100001001;
      patterns[22608] = 29'b0_101100001010_000_0_101100001010;
      patterns[22609] = 29'b0_101100001010_001_0_001010101100;
      patterns[22610] = 29'b0_101100001010_010_1_011000010100;
      patterns[22611] = 29'b0_101100001010_011_0_110000101001;
      patterns[22612] = 29'b0_101100001010_100_0_010110000101;
      patterns[22613] = 29'b0_101100001010_101_1_001011000010;
      patterns[22614] = 29'b0_101100001010_110_0_101100001010;
      patterns[22615] = 29'b0_101100001010_111_0_101100001010;
      patterns[22616] = 29'b0_101100001011_000_0_101100001011;
      patterns[22617] = 29'b0_101100001011_001_0_001011101100;
      patterns[22618] = 29'b0_101100001011_010_1_011000010110;
      patterns[22619] = 29'b0_101100001011_011_0_110000101101;
      patterns[22620] = 29'b0_101100001011_100_1_010110000101;
      patterns[22621] = 29'b0_101100001011_101_1_101011000010;
      patterns[22622] = 29'b0_101100001011_110_0_101100001011;
      patterns[22623] = 29'b0_101100001011_111_0_101100001011;
      patterns[22624] = 29'b0_101100001100_000_0_101100001100;
      patterns[22625] = 29'b0_101100001100_001_0_001100101100;
      patterns[22626] = 29'b0_101100001100_010_1_011000011000;
      patterns[22627] = 29'b0_101100001100_011_0_110000110001;
      patterns[22628] = 29'b0_101100001100_100_0_010110000110;
      patterns[22629] = 29'b0_101100001100_101_0_001011000011;
      patterns[22630] = 29'b0_101100001100_110_0_101100001100;
      patterns[22631] = 29'b0_101100001100_111_0_101100001100;
      patterns[22632] = 29'b0_101100001101_000_0_101100001101;
      patterns[22633] = 29'b0_101100001101_001_0_001101101100;
      patterns[22634] = 29'b0_101100001101_010_1_011000011010;
      patterns[22635] = 29'b0_101100001101_011_0_110000110101;
      patterns[22636] = 29'b0_101100001101_100_1_010110000110;
      patterns[22637] = 29'b0_101100001101_101_0_101011000011;
      patterns[22638] = 29'b0_101100001101_110_0_101100001101;
      patterns[22639] = 29'b0_101100001101_111_0_101100001101;
      patterns[22640] = 29'b0_101100001110_000_0_101100001110;
      patterns[22641] = 29'b0_101100001110_001_0_001110101100;
      patterns[22642] = 29'b0_101100001110_010_1_011000011100;
      patterns[22643] = 29'b0_101100001110_011_0_110000111001;
      patterns[22644] = 29'b0_101100001110_100_0_010110000111;
      patterns[22645] = 29'b0_101100001110_101_1_001011000011;
      patterns[22646] = 29'b0_101100001110_110_0_101100001110;
      patterns[22647] = 29'b0_101100001110_111_0_101100001110;
      patterns[22648] = 29'b0_101100001111_000_0_101100001111;
      patterns[22649] = 29'b0_101100001111_001_0_001111101100;
      patterns[22650] = 29'b0_101100001111_010_1_011000011110;
      patterns[22651] = 29'b0_101100001111_011_0_110000111101;
      patterns[22652] = 29'b0_101100001111_100_1_010110000111;
      patterns[22653] = 29'b0_101100001111_101_1_101011000011;
      patterns[22654] = 29'b0_101100001111_110_0_101100001111;
      patterns[22655] = 29'b0_101100001111_111_0_101100001111;
      patterns[22656] = 29'b0_101100010000_000_0_101100010000;
      patterns[22657] = 29'b0_101100010000_001_0_010000101100;
      patterns[22658] = 29'b0_101100010000_010_1_011000100000;
      patterns[22659] = 29'b0_101100010000_011_0_110001000001;
      patterns[22660] = 29'b0_101100010000_100_0_010110001000;
      patterns[22661] = 29'b0_101100010000_101_0_001011000100;
      patterns[22662] = 29'b0_101100010000_110_0_101100010000;
      patterns[22663] = 29'b0_101100010000_111_0_101100010000;
      patterns[22664] = 29'b0_101100010001_000_0_101100010001;
      patterns[22665] = 29'b0_101100010001_001_0_010001101100;
      patterns[22666] = 29'b0_101100010001_010_1_011000100010;
      patterns[22667] = 29'b0_101100010001_011_0_110001000101;
      patterns[22668] = 29'b0_101100010001_100_1_010110001000;
      patterns[22669] = 29'b0_101100010001_101_0_101011000100;
      patterns[22670] = 29'b0_101100010001_110_0_101100010001;
      patterns[22671] = 29'b0_101100010001_111_0_101100010001;
      patterns[22672] = 29'b0_101100010010_000_0_101100010010;
      patterns[22673] = 29'b0_101100010010_001_0_010010101100;
      patterns[22674] = 29'b0_101100010010_010_1_011000100100;
      patterns[22675] = 29'b0_101100010010_011_0_110001001001;
      patterns[22676] = 29'b0_101100010010_100_0_010110001001;
      patterns[22677] = 29'b0_101100010010_101_1_001011000100;
      patterns[22678] = 29'b0_101100010010_110_0_101100010010;
      patterns[22679] = 29'b0_101100010010_111_0_101100010010;
      patterns[22680] = 29'b0_101100010011_000_0_101100010011;
      patterns[22681] = 29'b0_101100010011_001_0_010011101100;
      patterns[22682] = 29'b0_101100010011_010_1_011000100110;
      patterns[22683] = 29'b0_101100010011_011_0_110001001101;
      patterns[22684] = 29'b0_101100010011_100_1_010110001001;
      patterns[22685] = 29'b0_101100010011_101_1_101011000100;
      patterns[22686] = 29'b0_101100010011_110_0_101100010011;
      patterns[22687] = 29'b0_101100010011_111_0_101100010011;
      patterns[22688] = 29'b0_101100010100_000_0_101100010100;
      patterns[22689] = 29'b0_101100010100_001_0_010100101100;
      patterns[22690] = 29'b0_101100010100_010_1_011000101000;
      patterns[22691] = 29'b0_101100010100_011_0_110001010001;
      patterns[22692] = 29'b0_101100010100_100_0_010110001010;
      patterns[22693] = 29'b0_101100010100_101_0_001011000101;
      patterns[22694] = 29'b0_101100010100_110_0_101100010100;
      patterns[22695] = 29'b0_101100010100_111_0_101100010100;
      patterns[22696] = 29'b0_101100010101_000_0_101100010101;
      patterns[22697] = 29'b0_101100010101_001_0_010101101100;
      patterns[22698] = 29'b0_101100010101_010_1_011000101010;
      patterns[22699] = 29'b0_101100010101_011_0_110001010101;
      patterns[22700] = 29'b0_101100010101_100_1_010110001010;
      patterns[22701] = 29'b0_101100010101_101_0_101011000101;
      patterns[22702] = 29'b0_101100010101_110_0_101100010101;
      patterns[22703] = 29'b0_101100010101_111_0_101100010101;
      patterns[22704] = 29'b0_101100010110_000_0_101100010110;
      patterns[22705] = 29'b0_101100010110_001_0_010110101100;
      patterns[22706] = 29'b0_101100010110_010_1_011000101100;
      patterns[22707] = 29'b0_101100010110_011_0_110001011001;
      patterns[22708] = 29'b0_101100010110_100_0_010110001011;
      patterns[22709] = 29'b0_101100010110_101_1_001011000101;
      patterns[22710] = 29'b0_101100010110_110_0_101100010110;
      patterns[22711] = 29'b0_101100010110_111_0_101100010110;
      patterns[22712] = 29'b0_101100010111_000_0_101100010111;
      patterns[22713] = 29'b0_101100010111_001_0_010111101100;
      patterns[22714] = 29'b0_101100010111_010_1_011000101110;
      patterns[22715] = 29'b0_101100010111_011_0_110001011101;
      patterns[22716] = 29'b0_101100010111_100_1_010110001011;
      patterns[22717] = 29'b0_101100010111_101_1_101011000101;
      patterns[22718] = 29'b0_101100010111_110_0_101100010111;
      patterns[22719] = 29'b0_101100010111_111_0_101100010111;
      patterns[22720] = 29'b0_101100011000_000_0_101100011000;
      patterns[22721] = 29'b0_101100011000_001_0_011000101100;
      patterns[22722] = 29'b0_101100011000_010_1_011000110000;
      patterns[22723] = 29'b0_101100011000_011_0_110001100001;
      patterns[22724] = 29'b0_101100011000_100_0_010110001100;
      patterns[22725] = 29'b0_101100011000_101_0_001011000110;
      patterns[22726] = 29'b0_101100011000_110_0_101100011000;
      patterns[22727] = 29'b0_101100011000_111_0_101100011000;
      patterns[22728] = 29'b0_101100011001_000_0_101100011001;
      patterns[22729] = 29'b0_101100011001_001_0_011001101100;
      patterns[22730] = 29'b0_101100011001_010_1_011000110010;
      patterns[22731] = 29'b0_101100011001_011_0_110001100101;
      patterns[22732] = 29'b0_101100011001_100_1_010110001100;
      patterns[22733] = 29'b0_101100011001_101_0_101011000110;
      patterns[22734] = 29'b0_101100011001_110_0_101100011001;
      patterns[22735] = 29'b0_101100011001_111_0_101100011001;
      patterns[22736] = 29'b0_101100011010_000_0_101100011010;
      patterns[22737] = 29'b0_101100011010_001_0_011010101100;
      patterns[22738] = 29'b0_101100011010_010_1_011000110100;
      patterns[22739] = 29'b0_101100011010_011_0_110001101001;
      patterns[22740] = 29'b0_101100011010_100_0_010110001101;
      patterns[22741] = 29'b0_101100011010_101_1_001011000110;
      patterns[22742] = 29'b0_101100011010_110_0_101100011010;
      patterns[22743] = 29'b0_101100011010_111_0_101100011010;
      patterns[22744] = 29'b0_101100011011_000_0_101100011011;
      patterns[22745] = 29'b0_101100011011_001_0_011011101100;
      patterns[22746] = 29'b0_101100011011_010_1_011000110110;
      patterns[22747] = 29'b0_101100011011_011_0_110001101101;
      patterns[22748] = 29'b0_101100011011_100_1_010110001101;
      patterns[22749] = 29'b0_101100011011_101_1_101011000110;
      patterns[22750] = 29'b0_101100011011_110_0_101100011011;
      patterns[22751] = 29'b0_101100011011_111_0_101100011011;
      patterns[22752] = 29'b0_101100011100_000_0_101100011100;
      patterns[22753] = 29'b0_101100011100_001_0_011100101100;
      patterns[22754] = 29'b0_101100011100_010_1_011000111000;
      patterns[22755] = 29'b0_101100011100_011_0_110001110001;
      patterns[22756] = 29'b0_101100011100_100_0_010110001110;
      patterns[22757] = 29'b0_101100011100_101_0_001011000111;
      patterns[22758] = 29'b0_101100011100_110_0_101100011100;
      patterns[22759] = 29'b0_101100011100_111_0_101100011100;
      patterns[22760] = 29'b0_101100011101_000_0_101100011101;
      patterns[22761] = 29'b0_101100011101_001_0_011101101100;
      patterns[22762] = 29'b0_101100011101_010_1_011000111010;
      patterns[22763] = 29'b0_101100011101_011_0_110001110101;
      patterns[22764] = 29'b0_101100011101_100_1_010110001110;
      patterns[22765] = 29'b0_101100011101_101_0_101011000111;
      patterns[22766] = 29'b0_101100011101_110_0_101100011101;
      patterns[22767] = 29'b0_101100011101_111_0_101100011101;
      patterns[22768] = 29'b0_101100011110_000_0_101100011110;
      patterns[22769] = 29'b0_101100011110_001_0_011110101100;
      patterns[22770] = 29'b0_101100011110_010_1_011000111100;
      patterns[22771] = 29'b0_101100011110_011_0_110001111001;
      patterns[22772] = 29'b0_101100011110_100_0_010110001111;
      patterns[22773] = 29'b0_101100011110_101_1_001011000111;
      patterns[22774] = 29'b0_101100011110_110_0_101100011110;
      patterns[22775] = 29'b0_101100011110_111_0_101100011110;
      patterns[22776] = 29'b0_101100011111_000_0_101100011111;
      patterns[22777] = 29'b0_101100011111_001_0_011111101100;
      patterns[22778] = 29'b0_101100011111_010_1_011000111110;
      patterns[22779] = 29'b0_101100011111_011_0_110001111101;
      patterns[22780] = 29'b0_101100011111_100_1_010110001111;
      patterns[22781] = 29'b0_101100011111_101_1_101011000111;
      patterns[22782] = 29'b0_101100011111_110_0_101100011111;
      patterns[22783] = 29'b0_101100011111_111_0_101100011111;
      patterns[22784] = 29'b0_101100100000_000_0_101100100000;
      patterns[22785] = 29'b0_101100100000_001_0_100000101100;
      patterns[22786] = 29'b0_101100100000_010_1_011001000000;
      patterns[22787] = 29'b0_101100100000_011_0_110010000001;
      patterns[22788] = 29'b0_101100100000_100_0_010110010000;
      patterns[22789] = 29'b0_101100100000_101_0_001011001000;
      patterns[22790] = 29'b0_101100100000_110_0_101100100000;
      patterns[22791] = 29'b0_101100100000_111_0_101100100000;
      patterns[22792] = 29'b0_101100100001_000_0_101100100001;
      patterns[22793] = 29'b0_101100100001_001_0_100001101100;
      patterns[22794] = 29'b0_101100100001_010_1_011001000010;
      patterns[22795] = 29'b0_101100100001_011_0_110010000101;
      patterns[22796] = 29'b0_101100100001_100_1_010110010000;
      patterns[22797] = 29'b0_101100100001_101_0_101011001000;
      patterns[22798] = 29'b0_101100100001_110_0_101100100001;
      patterns[22799] = 29'b0_101100100001_111_0_101100100001;
      patterns[22800] = 29'b0_101100100010_000_0_101100100010;
      patterns[22801] = 29'b0_101100100010_001_0_100010101100;
      patterns[22802] = 29'b0_101100100010_010_1_011001000100;
      patterns[22803] = 29'b0_101100100010_011_0_110010001001;
      patterns[22804] = 29'b0_101100100010_100_0_010110010001;
      patterns[22805] = 29'b0_101100100010_101_1_001011001000;
      patterns[22806] = 29'b0_101100100010_110_0_101100100010;
      patterns[22807] = 29'b0_101100100010_111_0_101100100010;
      patterns[22808] = 29'b0_101100100011_000_0_101100100011;
      patterns[22809] = 29'b0_101100100011_001_0_100011101100;
      patterns[22810] = 29'b0_101100100011_010_1_011001000110;
      patterns[22811] = 29'b0_101100100011_011_0_110010001101;
      patterns[22812] = 29'b0_101100100011_100_1_010110010001;
      patterns[22813] = 29'b0_101100100011_101_1_101011001000;
      patterns[22814] = 29'b0_101100100011_110_0_101100100011;
      patterns[22815] = 29'b0_101100100011_111_0_101100100011;
      patterns[22816] = 29'b0_101100100100_000_0_101100100100;
      patterns[22817] = 29'b0_101100100100_001_0_100100101100;
      patterns[22818] = 29'b0_101100100100_010_1_011001001000;
      patterns[22819] = 29'b0_101100100100_011_0_110010010001;
      patterns[22820] = 29'b0_101100100100_100_0_010110010010;
      patterns[22821] = 29'b0_101100100100_101_0_001011001001;
      patterns[22822] = 29'b0_101100100100_110_0_101100100100;
      patterns[22823] = 29'b0_101100100100_111_0_101100100100;
      patterns[22824] = 29'b0_101100100101_000_0_101100100101;
      patterns[22825] = 29'b0_101100100101_001_0_100101101100;
      patterns[22826] = 29'b0_101100100101_010_1_011001001010;
      patterns[22827] = 29'b0_101100100101_011_0_110010010101;
      patterns[22828] = 29'b0_101100100101_100_1_010110010010;
      patterns[22829] = 29'b0_101100100101_101_0_101011001001;
      patterns[22830] = 29'b0_101100100101_110_0_101100100101;
      patterns[22831] = 29'b0_101100100101_111_0_101100100101;
      patterns[22832] = 29'b0_101100100110_000_0_101100100110;
      patterns[22833] = 29'b0_101100100110_001_0_100110101100;
      patterns[22834] = 29'b0_101100100110_010_1_011001001100;
      patterns[22835] = 29'b0_101100100110_011_0_110010011001;
      patterns[22836] = 29'b0_101100100110_100_0_010110010011;
      patterns[22837] = 29'b0_101100100110_101_1_001011001001;
      patterns[22838] = 29'b0_101100100110_110_0_101100100110;
      patterns[22839] = 29'b0_101100100110_111_0_101100100110;
      patterns[22840] = 29'b0_101100100111_000_0_101100100111;
      patterns[22841] = 29'b0_101100100111_001_0_100111101100;
      patterns[22842] = 29'b0_101100100111_010_1_011001001110;
      patterns[22843] = 29'b0_101100100111_011_0_110010011101;
      patterns[22844] = 29'b0_101100100111_100_1_010110010011;
      patterns[22845] = 29'b0_101100100111_101_1_101011001001;
      patterns[22846] = 29'b0_101100100111_110_0_101100100111;
      patterns[22847] = 29'b0_101100100111_111_0_101100100111;
      patterns[22848] = 29'b0_101100101000_000_0_101100101000;
      patterns[22849] = 29'b0_101100101000_001_0_101000101100;
      patterns[22850] = 29'b0_101100101000_010_1_011001010000;
      patterns[22851] = 29'b0_101100101000_011_0_110010100001;
      patterns[22852] = 29'b0_101100101000_100_0_010110010100;
      patterns[22853] = 29'b0_101100101000_101_0_001011001010;
      patterns[22854] = 29'b0_101100101000_110_0_101100101000;
      patterns[22855] = 29'b0_101100101000_111_0_101100101000;
      patterns[22856] = 29'b0_101100101001_000_0_101100101001;
      patterns[22857] = 29'b0_101100101001_001_0_101001101100;
      patterns[22858] = 29'b0_101100101001_010_1_011001010010;
      patterns[22859] = 29'b0_101100101001_011_0_110010100101;
      patterns[22860] = 29'b0_101100101001_100_1_010110010100;
      patterns[22861] = 29'b0_101100101001_101_0_101011001010;
      patterns[22862] = 29'b0_101100101001_110_0_101100101001;
      patterns[22863] = 29'b0_101100101001_111_0_101100101001;
      patterns[22864] = 29'b0_101100101010_000_0_101100101010;
      patterns[22865] = 29'b0_101100101010_001_0_101010101100;
      patterns[22866] = 29'b0_101100101010_010_1_011001010100;
      patterns[22867] = 29'b0_101100101010_011_0_110010101001;
      patterns[22868] = 29'b0_101100101010_100_0_010110010101;
      patterns[22869] = 29'b0_101100101010_101_1_001011001010;
      patterns[22870] = 29'b0_101100101010_110_0_101100101010;
      patterns[22871] = 29'b0_101100101010_111_0_101100101010;
      patterns[22872] = 29'b0_101100101011_000_0_101100101011;
      patterns[22873] = 29'b0_101100101011_001_0_101011101100;
      patterns[22874] = 29'b0_101100101011_010_1_011001010110;
      patterns[22875] = 29'b0_101100101011_011_0_110010101101;
      patterns[22876] = 29'b0_101100101011_100_1_010110010101;
      patterns[22877] = 29'b0_101100101011_101_1_101011001010;
      patterns[22878] = 29'b0_101100101011_110_0_101100101011;
      patterns[22879] = 29'b0_101100101011_111_0_101100101011;
      patterns[22880] = 29'b0_101100101100_000_0_101100101100;
      patterns[22881] = 29'b0_101100101100_001_0_101100101100;
      patterns[22882] = 29'b0_101100101100_010_1_011001011000;
      patterns[22883] = 29'b0_101100101100_011_0_110010110001;
      patterns[22884] = 29'b0_101100101100_100_0_010110010110;
      patterns[22885] = 29'b0_101100101100_101_0_001011001011;
      patterns[22886] = 29'b0_101100101100_110_0_101100101100;
      patterns[22887] = 29'b0_101100101100_111_0_101100101100;
      patterns[22888] = 29'b0_101100101101_000_0_101100101101;
      patterns[22889] = 29'b0_101100101101_001_0_101101101100;
      patterns[22890] = 29'b0_101100101101_010_1_011001011010;
      patterns[22891] = 29'b0_101100101101_011_0_110010110101;
      patterns[22892] = 29'b0_101100101101_100_1_010110010110;
      patterns[22893] = 29'b0_101100101101_101_0_101011001011;
      patterns[22894] = 29'b0_101100101101_110_0_101100101101;
      patterns[22895] = 29'b0_101100101101_111_0_101100101101;
      patterns[22896] = 29'b0_101100101110_000_0_101100101110;
      patterns[22897] = 29'b0_101100101110_001_0_101110101100;
      patterns[22898] = 29'b0_101100101110_010_1_011001011100;
      patterns[22899] = 29'b0_101100101110_011_0_110010111001;
      patterns[22900] = 29'b0_101100101110_100_0_010110010111;
      patterns[22901] = 29'b0_101100101110_101_1_001011001011;
      patterns[22902] = 29'b0_101100101110_110_0_101100101110;
      patterns[22903] = 29'b0_101100101110_111_0_101100101110;
      patterns[22904] = 29'b0_101100101111_000_0_101100101111;
      patterns[22905] = 29'b0_101100101111_001_0_101111101100;
      patterns[22906] = 29'b0_101100101111_010_1_011001011110;
      patterns[22907] = 29'b0_101100101111_011_0_110010111101;
      patterns[22908] = 29'b0_101100101111_100_1_010110010111;
      patterns[22909] = 29'b0_101100101111_101_1_101011001011;
      patterns[22910] = 29'b0_101100101111_110_0_101100101111;
      patterns[22911] = 29'b0_101100101111_111_0_101100101111;
      patterns[22912] = 29'b0_101100110000_000_0_101100110000;
      patterns[22913] = 29'b0_101100110000_001_0_110000101100;
      patterns[22914] = 29'b0_101100110000_010_1_011001100000;
      patterns[22915] = 29'b0_101100110000_011_0_110011000001;
      patterns[22916] = 29'b0_101100110000_100_0_010110011000;
      patterns[22917] = 29'b0_101100110000_101_0_001011001100;
      patterns[22918] = 29'b0_101100110000_110_0_101100110000;
      patterns[22919] = 29'b0_101100110000_111_0_101100110000;
      patterns[22920] = 29'b0_101100110001_000_0_101100110001;
      patterns[22921] = 29'b0_101100110001_001_0_110001101100;
      patterns[22922] = 29'b0_101100110001_010_1_011001100010;
      patterns[22923] = 29'b0_101100110001_011_0_110011000101;
      patterns[22924] = 29'b0_101100110001_100_1_010110011000;
      patterns[22925] = 29'b0_101100110001_101_0_101011001100;
      patterns[22926] = 29'b0_101100110001_110_0_101100110001;
      patterns[22927] = 29'b0_101100110001_111_0_101100110001;
      patterns[22928] = 29'b0_101100110010_000_0_101100110010;
      patterns[22929] = 29'b0_101100110010_001_0_110010101100;
      patterns[22930] = 29'b0_101100110010_010_1_011001100100;
      patterns[22931] = 29'b0_101100110010_011_0_110011001001;
      patterns[22932] = 29'b0_101100110010_100_0_010110011001;
      patterns[22933] = 29'b0_101100110010_101_1_001011001100;
      patterns[22934] = 29'b0_101100110010_110_0_101100110010;
      patterns[22935] = 29'b0_101100110010_111_0_101100110010;
      patterns[22936] = 29'b0_101100110011_000_0_101100110011;
      patterns[22937] = 29'b0_101100110011_001_0_110011101100;
      patterns[22938] = 29'b0_101100110011_010_1_011001100110;
      patterns[22939] = 29'b0_101100110011_011_0_110011001101;
      patterns[22940] = 29'b0_101100110011_100_1_010110011001;
      patterns[22941] = 29'b0_101100110011_101_1_101011001100;
      patterns[22942] = 29'b0_101100110011_110_0_101100110011;
      patterns[22943] = 29'b0_101100110011_111_0_101100110011;
      patterns[22944] = 29'b0_101100110100_000_0_101100110100;
      patterns[22945] = 29'b0_101100110100_001_0_110100101100;
      patterns[22946] = 29'b0_101100110100_010_1_011001101000;
      patterns[22947] = 29'b0_101100110100_011_0_110011010001;
      patterns[22948] = 29'b0_101100110100_100_0_010110011010;
      patterns[22949] = 29'b0_101100110100_101_0_001011001101;
      patterns[22950] = 29'b0_101100110100_110_0_101100110100;
      patterns[22951] = 29'b0_101100110100_111_0_101100110100;
      patterns[22952] = 29'b0_101100110101_000_0_101100110101;
      patterns[22953] = 29'b0_101100110101_001_0_110101101100;
      patterns[22954] = 29'b0_101100110101_010_1_011001101010;
      patterns[22955] = 29'b0_101100110101_011_0_110011010101;
      patterns[22956] = 29'b0_101100110101_100_1_010110011010;
      patterns[22957] = 29'b0_101100110101_101_0_101011001101;
      patterns[22958] = 29'b0_101100110101_110_0_101100110101;
      patterns[22959] = 29'b0_101100110101_111_0_101100110101;
      patterns[22960] = 29'b0_101100110110_000_0_101100110110;
      patterns[22961] = 29'b0_101100110110_001_0_110110101100;
      patterns[22962] = 29'b0_101100110110_010_1_011001101100;
      patterns[22963] = 29'b0_101100110110_011_0_110011011001;
      patterns[22964] = 29'b0_101100110110_100_0_010110011011;
      patterns[22965] = 29'b0_101100110110_101_1_001011001101;
      patterns[22966] = 29'b0_101100110110_110_0_101100110110;
      patterns[22967] = 29'b0_101100110110_111_0_101100110110;
      patterns[22968] = 29'b0_101100110111_000_0_101100110111;
      patterns[22969] = 29'b0_101100110111_001_0_110111101100;
      patterns[22970] = 29'b0_101100110111_010_1_011001101110;
      patterns[22971] = 29'b0_101100110111_011_0_110011011101;
      patterns[22972] = 29'b0_101100110111_100_1_010110011011;
      patterns[22973] = 29'b0_101100110111_101_1_101011001101;
      patterns[22974] = 29'b0_101100110111_110_0_101100110111;
      patterns[22975] = 29'b0_101100110111_111_0_101100110111;
      patterns[22976] = 29'b0_101100111000_000_0_101100111000;
      patterns[22977] = 29'b0_101100111000_001_0_111000101100;
      patterns[22978] = 29'b0_101100111000_010_1_011001110000;
      patterns[22979] = 29'b0_101100111000_011_0_110011100001;
      patterns[22980] = 29'b0_101100111000_100_0_010110011100;
      patterns[22981] = 29'b0_101100111000_101_0_001011001110;
      patterns[22982] = 29'b0_101100111000_110_0_101100111000;
      patterns[22983] = 29'b0_101100111000_111_0_101100111000;
      patterns[22984] = 29'b0_101100111001_000_0_101100111001;
      patterns[22985] = 29'b0_101100111001_001_0_111001101100;
      patterns[22986] = 29'b0_101100111001_010_1_011001110010;
      patterns[22987] = 29'b0_101100111001_011_0_110011100101;
      patterns[22988] = 29'b0_101100111001_100_1_010110011100;
      patterns[22989] = 29'b0_101100111001_101_0_101011001110;
      patterns[22990] = 29'b0_101100111001_110_0_101100111001;
      patterns[22991] = 29'b0_101100111001_111_0_101100111001;
      patterns[22992] = 29'b0_101100111010_000_0_101100111010;
      patterns[22993] = 29'b0_101100111010_001_0_111010101100;
      patterns[22994] = 29'b0_101100111010_010_1_011001110100;
      patterns[22995] = 29'b0_101100111010_011_0_110011101001;
      patterns[22996] = 29'b0_101100111010_100_0_010110011101;
      patterns[22997] = 29'b0_101100111010_101_1_001011001110;
      patterns[22998] = 29'b0_101100111010_110_0_101100111010;
      patterns[22999] = 29'b0_101100111010_111_0_101100111010;
      patterns[23000] = 29'b0_101100111011_000_0_101100111011;
      patterns[23001] = 29'b0_101100111011_001_0_111011101100;
      patterns[23002] = 29'b0_101100111011_010_1_011001110110;
      patterns[23003] = 29'b0_101100111011_011_0_110011101101;
      patterns[23004] = 29'b0_101100111011_100_1_010110011101;
      patterns[23005] = 29'b0_101100111011_101_1_101011001110;
      patterns[23006] = 29'b0_101100111011_110_0_101100111011;
      patterns[23007] = 29'b0_101100111011_111_0_101100111011;
      patterns[23008] = 29'b0_101100111100_000_0_101100111100;
      patterns[23009] = 29'b0_101100111100_001_0_111100101100;
      patterns[23010] = 29'b0_101100111100_010_1_011001111000;
      patterns[23011] = 29'b0_101100111100_011_0_110011110001;
      patterns[23012] = 29'b0_101100111100_100_0_010110011110;
      patterns[23013] = 29'b0_101100111100_101_0_001011001111;
      patterns[23014] = 29'b0_101100111100_110_0_101100111100;
      patterns[23015] = 29'b0_101100111100_111_0_101100111100;
      patterns[23016] = 29'b0_101100111101_000_0_101100111101;
      patterns[23017] = 29'b0_101100111101_001_0_111101101100;
      patterns[23018] = 29'b0_101100111101_010_1_011001111010;
      patterns[23019] = 29'b0_101100111101_011_0_110011110101;
      patterns[23020] = 29'b0_101100111101_100_1_010110011110;
      patterns[23021] = 29'b0_101100111101_101_0_101011001111;
      patterns[23022] = 29'b0_101100111101_110_0_101100111101;
      patterns[23023] = 29'b0_101100111101_111_0_101100111101;
      patterns[23024] = 29'b0_101100111110_000_0_101100111110;
      patterns[23025] = 29'b0_101100111110_001_0_111110101100;
      patterns[23026] = 29'b0_101100111110_010_1_011001111100;
      patterns[23027] = 29'b0_101100111110_011_0_110011111001;
      patterns[23028] = 29'b0_101100111110_100_0_010110011111;
      patterns[23029] = 29'b0_101100111110_101_1_001011001111;
      patterns[23030] = 29'b0_101100111110_110_0_101100111110;
      patterns[23031] = 29'b0_101100111110_111_0_101100111110;
      patterns[23032] = 29'b0_101100111111_000_0_101100111111;
      patterns[23033] = 29'b0_101100111111_001_0_111111101100;
      patterns[23034] = 29'b0_101100111111_010_1_011001111110;
      patterns[23035] = 29'b0_101100111111_011_0_110011111101;
      patterns[23036] = 29'b0_101100111111_100_1_010110011111;
      patterns[23037] = 29'b0_101100111111_101_1_101011001111;
      patterns[23038] = 29'b0_101100111111_110_0_101100111111;
      patterns[23039] = 29'b0_101100111111_111_0_101100111111;
      patterns[23040] = 29'b0_101101000000_000_0_101101000000;
      patterns[23041] = 29'b0_101101000000_001_0_000000101101;
      patterns[23042] = 29'b0_101101000000_010_1_011010000000;
      patterns[23043] = 29'b0_101101000000_011_0_110100000001;
      patterns[23044] = 29'b0_101101000000_100_0_010110100000;
      patterns[23045] = 29'b0_101101000000_101_0_001011010000;
      patterns[23046] = 29'b0_101101000000_110_0_101101000000;
      patterns[23047] = 29'b0_101101000000_111_0_101101000000;
      patterns[23048] = 29'b0_101101000001_000_0_101101000001;
      patterns[23049] = 29'b0_101101000001_001_0_000001101101;
      patterns[23050] = 29'b0_101101000001_010_1_011010000010;
      patterns[23051] = 29'b0_101101000001_011_0_110100000101;
      patterns[23052] = 29'b0_101101000001_100_1_010110100000;
      patterns[23053] = 29'b0_101101000001_101_0_101011010000;
      patterns[23054] = 29'b0_101101000001_110_0_101101000001;
      patterns[23055] = 29'b0_101101000001_111_0_101101000001;
      patterns[23056] = 29'b0_101101000010_000_0_101101000010;
      patterns[23057] = 29'b0_101101000010_001_0_000010101101;
      patterns[23058] = 29'b0_101101000010_010_1_011010000100;
      patterns[23059] = 29'b0_101101000010_011_0_110100001001;
      patterns[23060] = 29'b0_101101000010_100_0_010110100001;
      patterns[23061] = 29'b0_101101000010_101_1_001011010000;
      patterns[23062] = 29'b0_101101000010_110_0_101101000010;
      patterns[23063] = 29'b0_101101000010_111_0_101101000010;
      patterns[23064] = 29'b0_101101000011_000_0_101101000011;
      patterns[23065] = 29'b0_101101000011_001_0_000011101101;
      patterns[23066] = 29'b0_101101000011_010_1_011010000110;
      patterns[23067] = 29'b0_101101000011_011_0_110100001101;
      patterns[23068] = 29'b0_101101000011_100_1_010110100001;
      patterns[23069] = 29'b0_101101000011_101_1_101011010000;
      patterns[23070] = 29'b0_101101000011_110_0_101101000011;
      patterns[23071] = 29'b0_101101000011_111_0_101101000011;
      patterns[23072] = 29'b0_101101000100_000_0_101101000100;
      patterns[23073] = 29'b0_101101000100_001_0_000100101101;
      patterns[23074] = 29'b0_101101000100_010_1_011010001000;
      patterns[23075] = 29'b0_101101000100_011_0_110100010001;
      patterns[23076] = 29'b0_101101000100_100_0_010110100010;
      patterns[23077] = 29'b0_101101000100_101_0_001011010001;
      patterns[23078] = 29'b0_101101000100_110_0_101101000100;
      patterns[23079] = 29'b0_101101000100_111_0_101101000100;
      patterns[23080] = 29'b0_101101000101_000_0_101101000101;
      patterns[23081] = 29'b0_101101000101_001_0_000101101101;
      patterns[23082] = 29'b0_101101000101_010_1_011010001010;
      patterns[23083] = 29'b0_101101000101_011_0_110100010101;
      patterns[23084] = 29'b0_101101000101_100_1_010110100010;
      patterns[23085] = 29'b0_101101000101_101_0_101011010001;
      patterns[23086] = 29'b0_101101000101_110_0_101101000101;
      patterns[23087] = 29'b0_101101000101_111_0_101101000101;
      patterns[23088] = 29'b0_101101000110_000_0_101101000110;
      patterns[23089] = 29'b0_101101000110_001_0_000110101101;
      patterns[23090] = 29'b0_101101000110_010_1_011010001100;
      patterns[23091] = 29'b0_101101000110_011_0_110100011001;
      patterns[23092] = 29'b0_101101000110_100_0_010110100011;
      patterns[23093] = 29'b0_101101000110_101_1_001011010001;
      patterns[23094] = 29'b0_101101000110_110_0_101101000110;
      patterns[23095] = 29'b0_101101000110_111_0_101101000110;
      patterns[23096] = 29'b0_101101000111_000_0_101101000111;
      patterns[23097] = 29'b0_101101000111_001_0_000111101101;
      patterns[23098] = 29'b0_101101000111_010_1_011010001110;
      patterns[23099] = 29'b0_101101000111_011_0_110100011101;
      patterns[23100] = 29'b0_101101000111_100_1_010110100011;
      patterns[23101] = 29'b0_101101000111_101_1_101011010001;
      patterns[23102] = 29'b0_101101000111_110_0_101101000111;
      patterns[23103] = 29'b0_101101000111_111_0_101101000111;
      patterns[23104] = 29'b0_101101001000_000_0_101101001000;
      patterns[23105] = 29'b0_101101001000_001_0_001000101101;
      patterns[23106] = 29'b0_101101001000_010_1_011010010000;
      patterns[23107] = 29'b0_101101001000_011_0_110100100001;
      patterns[23108] = 29'b0_101101001000_100_0_010110100100;
      patterns[23109] = 29'b0_101101001000_101_0_001011010010;
      patterns[23110] = 29'b0_101101001000_110_0_101101001000;
      patterns[23111] = 29'b0_101101001000_111_0_101101001000;
      patterns[23112] = 29'b0_101101001001_000_0_101101001001;
      patterns[23113] = 29'b0_101101001001_001_0_001001101101;
      patterns[23114] = 29'b0_101101001001_010_1_011010010010;
      patterns[23115] = 29'b0_101101001001_011_0_110100100101;
      patterns[23116] = 29'b0_101101001001_100_1_010110100100;
      patterns[23117] = 29'b0_101101001001_101_0_101011010010;
      patterns[23118] = 29'b0_101101001001_110_0_101101001001;
      patterns[23119] = 29'b0_101101001001_111_0_101101001001;
      patterns[23120] = 29'b0_101101001010_000_0_101101001010;
      patterns[23121] = 29'b0_101101001010_001_0_001010101101;
      patterns[23122] = 29'b0_101101001010_010_1_011010010100;
      patterns[23123] = 29'b0_101101001010_011_0_110100101001;
      patterns[23124] = 29'b0_101101001010_100_0_010110100101;
      patterns[23125] = 29'b0_101101001010_101_1_001011010010;
      patterns[23126] = 29'b0_101101001010_110_0_101101001010;
      patterns[23127] = 29'b0_101101001010_111_0_101101001010;
      patterns[23128] = 29'b0_101101001011_000_0_101101001011;
      patterns[23129] = 29'b0_101101001011_001_0_001011101101;
      patterns[23130] = 29'b0_101101001011_010_1_011010010110;
      patterns[23131] = 29'b0_101101001011_011_0_110100101101;
      patterns[23132] = 29'b0_101101001011_100_1_010110100101;
      patterns[23133] = 29'b0_101101001011_101_1_101011010010;
      patterns[23134] = 29'b0_101101001011_110_0_101101001011;
      patterns[23135] = 29'b0_101101001011_111_0_101101001011;
      patterns[23136] = 29'b0_101101001100_000_0_101101001100;
      patterns[23137] = 29'b0_101101001100_001_0_001100101101;
      patterns[23138] = 29'b0_101101001100_010_1_011010011000;
      patterns[23139] = 29'b0_101101001100_011_0_110100110001;
      patterns[23140] = 29'b0_101101001100_100_0_010110100110;
      patterns[23141] = 29'b0_101101001100_101_0_001011010011;
      patterns[23142] = 29'b0_101101001100_110_0_101101001100;
      patterns[23143] = 29'b0_101101001100_111_0_101101001100;
      patterns[23144] = 29'b0_101101001101_000_0_101101001101;
      patterns[23145] = 29'b0_101101001101_001_0_001101101101;
      patterns[23146] = 29'b0_101101001101_010_1_011010011010;
      patterns[23147] = 29'b0_101101001101_011_0_110100110101;
      patterns[23148] = 29'b0_101101001101_100_1_010110100110;
      patterns[23149] = 29'b0_101101001101_101_0_101011010011;
      patterns[23150] = 29'b0_101101001101_110_0_101101001101;
      patterns[23151] = 29'b0_101101001101_111_0_101101001101;
      patterns[23152] = 29'b0_101101001110_000_0_101101001110;
      patterns[23153] = 29'b0_101101001110_001_0_001110101101;
      patterns[23154] = 29'b0_101101001110_010_1_011010011100;
      patterns[23155] = 29'b0_101101001110_011_0_110100111001;
      patterns[23156] = 29'b0_101101001110_100_0_010110100111;
      patterns[23157] = 29'b0_101101001110_101_1_001011010011;
      patterns[23158] = 29'b0_101101001110_110_0_101101001110;
      patterns[23159] = 29'b0_101101001110_111_0_101101001110;
      patterns[23160] = 29'b0_101101001111_000_0_101101001111;
      patterns[23161] = 29'b0_101101001111_001_0_001111101101;
      patterns[23162] = 29'b0_101101001111_010_1_011010011110;
      patterns[23163] = 29'b0_101101001111_011_0_110100111101;
      patterns[23164] = 29'b0_101101001111_100_1_010110100111;
      patterns[23165] = 29'b0_101101001111_101_1_101011010011;
      patterns[23166] = 29'b0_101101001111_110_0_101101001111;
      patterns[23167] = 29'b0_101101001111_111_0_101101001111;
      patterns[23168] = 29'b0_101101010000_000_0_101101010000;
      patterns[23169] = 29'b0_101101010000_001_0_010000101101;
      patterns[23170] = 29'b0_101101010000_010_1_011010100000;
      patterns[23171] = 29'b0_101101010000_011_0_110101000001;
      patterns[23172] = 29'b0_101101010000_100_0_010110101000;
      patterns[23173] = 29'b0_101101010000_101_0_001011010100;
      patterns[23174] = 29'b0_101101010000_110_0_101101010000;
      patterns[23175] = 29'b0_101101010000_111_0_101101010000;
      patterns[23176] = 29'b0_101101010001_000_0_101101010001;
      patterns[23177] = 29'b0_101101010001_001_0_010001101101;
      patterns[23178] = 29'b0_101101010001_010_1_011010100010;
      patterns[23179] = 29'b0_101101010001_011_0_110101000101;
      patterns[23180] = 29'b0_101101010001_100_1_010110101000;
      patterns[23181] = 29'b0_101101010001_101_0_101011010100;
      patterns[23182] = 29'b0_101101010001_110_0_101101010001;
      patterns[23183] = 29'b0_101101010001_111_0_101101010001;
      patterns[23184] = 29'b0_101101010010_000_0_101101010010;
      patterns[23185] = 29'b0_101101010010_001_0_010010101101;
      patterns[23186] = 29'b0_101101010010_010_1_011010100100;
      patterns[23187] = 29'b0_101101010010_011_0_110101001001;
      patterns[23188] = 29'b0_101101010010_100_0_010110101001;
      patterns[23189] = 29'b0_101101010010_101_1_001011010100;
      patterns[23190] = 29'b0_101101010010_110_0_101101010010;
      patterns[23191] = 29'b0_101101010010_111_0_101101010010;
      patterns[23192] = 29'b0_101101010011_000_0_101101010011;
      patterns[23193] = 29'b0_101101010011_001_0_010011101101;
      patterns[23194] = 29'b0_101101010011_010_1_011010100110;
      patterns[23195] = 29'b0_101101010011_011_0_110101001101;
      patterns[23196] = 29'b0_101101010011_100_1_010110101001;
      patterns[23197] = 29'b0_101101010011_101_1_101011010100;
      patterns[23198] = 29'b0_101101010011_110_0_101101010011;
      patterns[23199] = 29'b0_101101010011_111_0_101101010011;
      patterns[23200] = 29'b0_101101010100_000_0_101101010100;
      patterns[23201] = 29'b0_101101010100_001_0_010100101101;
      patterns[23202] = 29'b0_101101010100_010_1_011010101000;
      patterns[23203] = 29'b0_101101010100_011_0_110101010001;
      patterns[23204] = 29'b0_101101010100_100_0_010110101010;
      patterns[23205] = 29'b0_101101010100_101_0_001011010101;
      patterns[23206] = 29'b0_101101010100_110_0_101101010100;
      patterns[23207] = 29'b0_101101010100_111_0_101101010100;
      patterns[23208] = 29'b0_101101010101_000_0_101101010101;
      patterns[23209] = 29'b0_101101010101_001_0_010101101101;
      patterns[23210] = 29'b0_101101010101_010_1_011010101010;
      patterns[23211] = 29'b0_101101010101_011_0_110101010101;
      patterns[23212] = 29'b0_101101010101_100_1_010110101010;
      patterns[23213] = 29'b0_101101010101_101_0_101011010101;
      patterns[23214] = 29'b0_101101010101_110_0_101101010101;
      patterns[23215] = 29'b0_101101010101_111_0_101101010101;
      patterns[23216] = 29'b0_101101010110_000_0_101101010110;
      patterns[23217] = 29'b0_101101010110_001_0_010110101101;
      patterns[23218] = 29'b0_101101010110_010_1_011010101100;
      patterns[23219] = 29'b0_101101010110_011_0_110101011001;
      patterns[23220] = 29'b0_101101010110_100_0_010110101011;
      patterns[23221] = 29'b0_101101010110_101_1_001011010101;
      patterns[23222] = 29'b0_101101010110_110_0_101101010110;
      patterns[23223] = 29'b0_101101010110_111_0_101101010110;
      patterns[23224] = 29'b0_101101010111_000_0_101101010111;
      patterns[23225] = 29'b0_101101010111_001_0_010111101101;
      patterns[23226] = 29'b0_101101010111_010_1_011010101110;
      patterns[23227] = 29'b0_101101010111_011_0_110101011101;
      patterns[23228] = 29'b0_101101010111_100_1_010110101011;
      patterns[23229] = 29'b0_101101010111_101_1_101011010101;
      patterns[23230] = 29'b0_101101010111_110_0_101101010111;
      patterns[23231] = 29'b0_101101010111_111_0_101101010111;
      patterns[23232] = 29'b0_101101011000_000_0_101101011000;
      patterns[23233] = 29'b0_101101011000_001_0_011000101101;
      patterns[23234] = 29'b0_101101011000_010_1_011010110000;
      patterns[23235] = 29'b0_101101011000_011_0_110101100001;
      patterns[23236] = 29'b0_101101011000_100_0_010110101100;
      patterns[23237] = 29'b0_101101011000_101_0_001011010110;
      patterns[23238] = 29'b0_101101011000_110_0_101101011000;
      patterns[23239] = 29'b0_101101011000_111_0_101101011000;
      patterns[23240] = 29'b0_101101011001_000_0_101101011001;
      patterns[23241] = 29'b0_101101011001_001_0_011001101101;
      patterns[23242] = 29'b0_101101011001_010_1_011010110010;
      patterns[23243] = 29'b0_101101011001_011_0_110101100101;
      patterns[23244] = 29'b0_101101011001_100_1_010110101100;
      patterns[23245] = 29'b0_101101011001_101_0_101011010110;
      patterns[23246] = 29'b0_101101011001_110_0_101101011001;
      patterns[23247] = 29'b0_101101011001_111_0_101101011001;
      patterns[23248] = 29'b0_101101011010_000_0_101101011010;
      patterns[23249] = 29'b0_101101011010_001_0_011010101101;
      patterns[23250] = 29'b0_101101011010_010_1_011010110100;
      patterns[23251] = 29'b0_101101011010_011_0_110101101001;
      patterns[23252] = 29'b0_101101011010_100_0_010110101101;
      patterns[23253] = 29'b0_101101011010_101_1_001011010110;
      patterns[23254] = 29'b0_101101011010_110_0_101101011010;
      patterns[23255] = 29'b0_101101011010_111_0_101101011010;
      patterns[23256] = 29'b0_101101011011_000_0_101101011011;
      patterns[23257] = 29'b0_101101011011_001_0_011011101101;
      patterns[23258] = 29'b0_101101011011_010_1_011010110110;
      patterns[23259] = 29'b0_101101011011_011_0_110101101101;
      patterns[23260] = 29'b0_101101011011_100_1_010110101101;
      patterns[23261] = 29'b0_101101011011_101_1_101011010110;
      patterns[23262] = 29'b0_101101011011_110_0_101101011011;
      patterns[23263] = 29'b0_101101011011_111_0_101101011011;
      patterns[23264] = 29'b0_101101011100_000_0_101101011100;
      patterns[23265] = 29'b0_101101011100_001_0_011100101101;
      patterns[23266] = 29'b0_101101011100_010_1_011010111000;
      patterns[23267] = 29'b0_101101011100_011_0_110101110001;
      patterns[23268] = 29'b0_101101011100_100_0_010110101110;
      patterns[23269] = 29'b0_101101011100_101_0_001011010111;
      patterns[23270] = 29'b0_101101011100_110_0_101101011100;
      patterns[23271] = 29'b0_101101011100_111_0_101101011100;
      patterns[23272] = 29'b0_101101011101_000_0_101101011101;
      patterns[23273] = 29'b0_101101011101_001_0_011101101101;
      patterns[23274] = 29'b0_101101011101_010_1_011010111010;
      patterns[23275] = 29'b0_101101011101_011_0_110101110101;
      patterns[23276] = 29'b0_101101011101_100_1_010110101110;
      patterns[23277] = 29'b0_101101011101_101_0_101011010111;
      patterns[23278] = 29'b0_101101011101_110_0_101101011101;
      patterns[23279] = 29'b0_101101011101_111_0_101101011101;
      patterns[23280] = 29'b0_101101011110_000_0_101101011110;
      patterns[23281] = 29'b0_101101011110_001_0_011110101101;
      patterns[23282] = 29'b0_101101011110_010_1_011010111100;
      patterns[23283] = 29'b0_101101011110_011_0_110101111001;
      patterns[23284] = 29'b0_101101011110_100_0_010110101111;
      patterns[23285] = 29'b0_101101011110_101_1_001011010111;
      patterns[23286] = 29'b0_101101011110_110_0_101101011110;
      patterns[23287] = 29'b0_101101011110_111_0_101101011110;
      patterns[23288] = 29'b0_101101011111_000_0_101101011111;
      patterns[23289] = 29'b0_101101011111_001_0_011111101101;
      patterns[23290] = 29'b0_101101011111_010_1_011010111110;
      patterns[23291] = 29'b0_101101011111_011_0_110101111101;
      patterns[23292] = 29'b0_101101011111_100_1_010110101111;
      patterns[23293] = 29'b0_101101011111_101_1_101011010111;
      patterns[23294] = 29'b0_101101011111_110_0_101101011111;
      patterns[23295] = 29'b0_101101011111_111_0_101101011111;
      patterns[23296] = 29'b0_101101100000_000_0_101101100000;
      patterns[23297] = 29'b0_101101100000_001_0_100000101101;
      patterns[23298] = 29'b0_101101100000_010_1_011011000000;
      patterns[23299] = 29'b0_101101100000_011_0_110110000001;
      patterns[23300] = 29'b0_101101100000_100_0_010110110000;
      patterns[23301] = 29'b0_101101100000_101_0_001011011000;
      patterns[23302] = 29'b0_101101100000_110_0_101101100000;
      patterns[23303] = 29'b0_101101100000_111_0_101101100000;
      patterns[23304] = 29'b0_101101100001_000_0_101101100001;
      patterns[23305] = 29'b0_101101100001_001_0_100001101101;
      patterns[23306] = 29'b0_101101100001_010_1_011011000010;
      patterns[23307] = 29'b0_101101100001_011_0_110110000101;
      patterns[23308] = 29'b0_101101100001_100_1_010110110000;
      patterns[23309] = 29'b0_101101100001_101_0_101011011000;
      patterns[23310] = 29'b0_101101100001_110_0_101101100001;
      patterns[23311] = 29'b0_101101100001_111_0_101101100001;
      patterns[23312] = 29'b0_101101100010_000_0_101101100010;
      patterns[23313] = 29'b0_101101100010_001_0_100010101101;
      patterns[23314] = 29'b0_101101100010_010_1_011011000100;
      patterns[23315] = 29'b0_101101100010_011_0_110110001001;
      patterns[23316] = 29'b0_101101100010_100_0_010110110001;
      patterns[23317] = 29'b0_101101100010_101_1_001011011000;
      patterns[23318] = 29'b0_101101100010_110_0_101101100010;
      patterns[23319] = 29'b0_101101100010_111_0_101101100010;
      patterns[23320] = 29'b0_101101100011_000_0_101101100011;
      patterns[23321] = 29'b0_101101100011_001_0_100011101101;
      patterns[23322] = 29'b0_101101100011_010_1_011011000110;
      patterns[23323] = 29'b0_101101100011_011_0_110110001101;
      patterns[23324] = 29'b0_101101100011_100_1_010110110001;
      patterns[23325] = 29'b0_101101100011_101_1_101011011000;
      patterns[23326] = 29'b0_101101100011_110_0_101101100011;
      patterns[23327] = 29'b0_101101100011_111_0_101101100011;
      patterns[23328] = 29'b0_101101100100_000_0_101101100100;
      patterns[23329] = 29'b0_101101100100_001_0_100100101101;
      patterns[23330] = 29'b0_101101100100_010_1_011011001000;
      patterns[23331] = 29'b0_101101100100_011_0_110110010001;
      patterns[23332] = 29'b0_101101100100_100_0_010110110010;
      patterns[23333] = 29'b0_101101100100_101_0_001011011001;
      patterns[23334] = 29'b0_101101100100_110_0_101101100100;
      patterns[23335] = 29'b0_101101100100_111_0_101101100100;
      patterns[23336] = 29'b0_101101100101_000_0_101101100101;
      patterns[23337] = 29'b0_101101100101_001_0_100101101101;
      patterns[23338] = 29'b0_101101100101_010_1_011011001010;
      patterns[23339] = 29'b0_101101100101_011_0_110110010101;
      patterns[23340] = 29'b0_101101100101_100_1_010110110010;
      patterns[23341] = 29'b0_101101100101_101_0_101011011001;
      patterns[23342] = 29'b0_101101100101_110_0_101101100101;
      patterns[23343] = 29'b0_101101100101_111_0_101101100101;
      patterns[23344] = 29'b0_101101100110_000_0_101101100110;
      patterns[23345] = 29'b0_101101100110_001_0_100110101101;
      patterns[23346] = 29'b0_101101100110_010_1_011011001100;
      patterns[23347] = 29'b0_101101100110_011_0_110110011001;
      patterns[23348] = 29'b0_101101100110_100_0_010110110011;
      patterns[23349] = 29'b0_101101100110_101_1_001011011001;
      patterns[23350] = 29'b0_101101100110_110_0_101101100110;
      patterns[23351] = 29'b0_101101100110_111_0_101101100110;
      patterns[23352] = 29'b0_101101100111_000_0_101101100111;
      patterns[23353] = 29'b0_101101100111_001_0_100111101101;
      patterns[23354] = 29'b0_101101100111_010_1_011011001110;
      patterns[23355] = 29'b0_101101100111_011_0_110110011101;
      patterns[23356] = 29'b0_101101100111_100_1_010110110011;
      patterns[23357] = 29'b0_101101100111_101_1_101011011001;
      patterns[23358] = 29'b0_101101100111_110_0_101101100111;
      patterns[23359] = 29'b0_101101100111_111_0_101101100111;
      patterns[23360] = 29'b0_101101101000_000_0_101101101000;
      patterns[23361] = 29'b0_101101101000_001_0_101000101101;
      patterns[23362] = 29'b0_101101101000_010_1_011011010000;
      patterns[23363] = 29'b0_101101101000_011_0_110110100001;
      patterns[23364] = 29'b0_101101101000_100_0_010110110100;
      patterns[23365] = 29'b0_101101101000_101_0_001011011010;
      patterns[23366] = 29'b0_101101101000_110_0_101101101000;
      patterns[23367] = 29'b0_101101101000_111_0_101101101000;
      patterns[23368] = 29'b0_101101101001_000_0_101101101001;
      patterns[23369] = 29'b0_101101101001_001_0_101001101101;
      patterns[23370] = 29'b0_101101101001_010_1_011011010010;
      patterns[23371] = 29'b0_101101101001_011_0_110110100101;
      patterns[23372] = 29'b0_101101101001_100_1_010110110100;
      patterns[23373] = 29'b0_101101101001_101_0_101011011010;
      patterns[23374] = 29'b0_101101101001_110_0_101101101001;
      patterns[23375] = 29'b0_101101101001_111_0_101101101001;
      patterns[23376] = 29'b0_101101101010_000_0_101101101010;
      patterns[23377] = 29'b0_101101101010_001_0_101010101101;
      patterns[23378] = 29'b0_101101101010_010_1_011011010100;
      patterns[23379] = 29'b0_101101101010_011_0_110110101001;
      patterns[23380] = 29'b0_101101101010_100_0_010110110101;
      patterns[23381] = 29'b0_101101101010_101_1_001011011010;
      patterns[23382] = 29'b0_101101101010_110_0_101101101010;
      patterns[23383] = 29'b0_101101101010_111_0_101101101010;
      patterns[23384] = 29'b0_101101101011_000_0_101101101011;
      patterns[23385] = 29'b0_101101101011_001_0_101011101101;
      patterns[23386] = 29'b0_101101101011_010_1_011011010110;
      patterns[23387] = 29'b0_101101101011_011_0_110110101101;
      patterns[23388] = 29'b0_101101101011_100_1_010110110101;
      patterns[23389] = 29'b0_101101101011_101_1_101011011010;
      patterns[23390] = 29'b0_101101101011_110_0_101101101011;
      patterns[23391] = 29'b0_101101101011_111_0_101101101011;
      patterns[23392] = 29'b0_101101101100_000_0_101101101100;
      patterns[23393] = 29'b0_101101101100_001_0_101100101101;
      patterns[23394] = 29'b0_101101101100_010_1_011011011000;
      patterns[23395] = 29'b0_101101101100_011_0_110110110001;
      patterns[23396] = 29'b0_101101101100_100_0_010110110110;
      patterns[23397] = 29'b0_101101101100_101_0_001011011011;
      patterns[23398] = 29'b0_101101101100_110_0_101101101100;
      patterns[23399] = 29'b0_101101101100_111_0_101101101100;
      patterns[23400] = 29'b0_101101101101_000_0_101101101101;
      patterns[23401] = 29'b0_101101101101_001_0_101101101101;
      patterns[23402] = 29'b0_101101101101_010_1_011011011010;
      patterns[23403] = 29'b0_101101101101_011_0_110110110101;
      patterns[23404] = 29'b0_101101101101_100_1_010110110110;
      patterns[23405] = 29'b0_101101101101_101_0_101011011011;
      patterns[23406] = 29'b0_101101101101_110_0_101101101101;
      patterns[23407] = 29'b0_101101101101_111_0_101101101101;
      patterns[23408] = 29'b0_101101101110_000_0_101101101110;
      patterns[23409] = 29'b0_101101101110_001_0_101110101101;
      patterns[23410] = 29'b0_101101101110_010_1_011011011100;
      patterns[23411] = 29'b0_101101101110_011_0_110110111001;
      patterns[23412] = 29'b0_101101101110_100_0_010110110111;
      patterns[23413] = 29'b0_101101101110_101_1_001011011011;
      patterns[23414] = 29'b0_101101101110_110_0_101101101110;
      patterns[23415] = 29'b0_101101101110_111_0_101101101110;
      patterns[23416] = 29'b0_101101101111_000_0_101101101111;
      patterns[23417] = 29'b0_101101101111_001_0_101111101101;
      patterns[23418] = 29'b0_101101101111_010_1_011011011110;
      patterns[23419] = 29'b0_101101101111_011_0_110110111101;
      patterns[23420] = 29'b0_101101101111_100_1_010110110111;
      patterns[23421] = 29'b0_101101101111_101_1_101011011011;
      patterns[23422] = 29'b0_101101101111_110_0_101101101111;
      patterns[23423] = 29'b0_101101101111_111_0_101101101111;
      patterns[23424] = 29'b0_101101110000_000_0_101101110000;
      patterns[23425] = 29'b0_101101110000_001_0_110000101101;
      patterns[23426] = 29'b0_101101110000_010_1_011011100000;
      patterns[23427] = 29'b0_101101110000_011_0_110111000001;
      patterns[23428] = 29'b0_101101110000_100_0_010110111000;
      patterns[23429] = 29'b0_101101110000_101_0_001011011100;
      patterns[23430] = 29'b0_101101110000_110_0_101101110000;
      patterns[23431] = 29'b0_101101110000_111_0_101101110000;
      patterns[23432] = 29'b0_101101110001_000_0_101101110001;
      patterns[23433] = 29'b0_101101110001_001_0_110001101101;
      patterns[23434] = 29'b0_101101110001_010_1_011011100010;
      patterns[23435] = 29'b0_101101110001_011_0_110111000101;
      patterns[23436] = 29'b0_101101110001_100_1_010110111000;
      patterns[23437] = 29'b0_101101110001_101_0_101011011100;
      patterns[23438] = 29'b0_101101110001_110_0_101101110001;
      patterns[23439] = 29'b0_101101110001_111_0_101101110001;
      patterns[23440] = 29'b0_101101110010_000_0_101101110010;
      patterns[23441] = 29'b0_101101110010_001_0_110010101101;
      patterns[23442] = 29'b0_101101110010_010_1_011011100100;
      patterns[23443] = 29'b0_101101110010_011_0_110111001001;
      patterns[23444] = 29'b0_101101110010_100_0_010110111001;
      patterns[23445] = 29'b0_101101110010_101_1_001011011100;
      patterns[23446] = 29'b0_101101110010_110_0_101101110010;
      patterns[23447] = 29'b0_101101110010_111_0_101101110010;
      patterns[23448] = 29'b0_101101110011_000_0_101101110011;
      patterns[23449] = 29'b0_101101110011_001_0_110011101101;
      patterns[23450] = 29'b0_101101110011_010_1_011011100110;
      patterns[23451] = 29'b0_101101110011_011_0_110111001101;
      patterns[23452] = 29'b0_101101110011_100_1_010110111001;
      patterns[23453] = 29'b0_101101110011_101_1_101011011100;
      patterns[23454] = 29'b0_101101110011_110_0_101101110011;
      patterns[23455] = 29'b0_101101110011_111_0_101101110011;
      patterns[23456] = 29'b0_101101110100_000_0_101101110100;
      patterns[23457] = 29'b0_101101110100_001_0_110100101101;
      patterns[23458] = 29'b0_101101110100_010_1_011011101000;
      patterns[23459] = 29'b0_101101110100_011_0_110111010001;
      patterns[23460] = 29'b0_101101110100_100_0_010110111010;
      patterns[23461] = 29'b0_101101110100_101_0_001011011101;
      patterns[23462] = 29'b0_101101110100_110_0_101101110100;
      patterns[23463] = 29'b0_101101110100_111_0_101101110100;
      patterns[23464] = 29'b0_101101110101_000_0_101101110101;
      patterns[23465] = 29'b0_101101110101_001_0_110101101101;
      patterns[23466] = 29'b0_101101110101_010_1_011011101010;
      patterns[23467] = 29'b0_101101110101_011_0_110111010101;
      patterns[23468] = 29'b0_101101110101_100_1_010110111010;
      patterns[23469] = 29'b0_101101110101_101_0_101011011101;
      patterns[23470] = 29'b0_101101110101_110_0_101101110101;
      patterns[23471] = 29'b0_101101110101_111_0_101101110101;
      patterns[23472] = 29'b0_101101110110_000_0_101101110110;
      patterns[23473] = 29'b0_101101110110_001_0_110110101101;
      patterns[23474] = 29'b0_101101110110_010_1_011011101100;
      patterns[23475] = 29'b0_101101110110_011_0_110111011001;
      patterns[23476] = 29'b0_101101110110_100_0_010110111011;
      patterns[23477] = 29'b0_101101110110_101_1_001011011101;
      patterns[23478] = 29'b0_101101110110_110_0_101101110110;
      patterns[23479] = 29'b0_101101110110_111_0_101101110110;
      patterns[23480] = 29'b0_101101110111_000_0_101101110111;
      patterns[23481] = 29'b0_101101110111_001_0_110111101101;
      patterns[23482] = 29'b0_101101110111_010_1_011011101110;
      patterns[23483] = 29'b0_101101110111_011_0_110111011101;
      patterns[23484] = 29'b0_101101110111_100_1_010110111011;
      patterns[23485] = 29'b0_101101110111_101_1_101011011101;
      patterns[23486] = 29'b0_101101110111_110_0_101101110111;
      patterns[23487] = 29'b0_101101110111_111_0_101101110111;
      patterns[23488] = 29'b0_101101111000_000_0_101101111000;
      patterns[23489] = 29'b0_101101111000_001_0_111000101101;
      patterns[23490] = 29'b0_101101111000_010_1_011011110000;
      patterns[23491] = 29'b0_101101111000_011_0_110111100001;
      patterns[23492] = 29'b0_101101111000_100_0_010110111100;
      patterns[23493] = 29'b0_101101111000_101_0_001011011110;
      patterns[23494] = 29'b0_101101111000_110_0_101101111000;
      patterns[23495] = 29'b0_101101111000_111_0_101101111000;
      patterns[23496] = 29'b0_101101111001_000_0_101101111001;
      patterns[23497] = 29'b0_101101111001_001_0_111001101101;
      patterns[23498] = 29'b0_101101111001_010_1_011011110010;
      patterns[23499] = 29'b0_101101111001_011_0_110111100101;
      patterns[23500] = 29'b0_101101111001_100_1_010110111100;
      patterns[23501] = 29'b0_101101111001_101_0_101011011110;
      patterns[23502] = 29'b0_101101111001_110_0_101101111001;
      patterns[23503] = 29'b0_101101111001_111_0_101101111001;
      patterns[23504] = 29'b0_101101111010_000_0_101101111010;
      patterns[23505] = 29'b0_101101111010_001_0_111010101101;
      patterns[23506] = 29'b0_101101111010_010_1_011011110100;
      patterns[23507] = 29'b0_101101111010_011_0_110111101001;
      patterns[23508] = 29'b0_101101111010_100_0_010110111101;
      patterns[23509] = 29'b0_101101111010_101_1_001011011110;
      patterns[23510] = 29'b0_101101111010_110_0_101101111010;
      patterns[23511] = 29'b0_101101111010_111_0_101101111010;
      patterns[23512] = 29'b0_101101111011_000_0_101101111011;
      patterns[23513] = 29'b0_101101111011_001_0_111011101101;
      patterns[23514] = 29'b0_101101111011_010_1_011011110110;
      patterns[23515] = 29'b0_101101111011_011_0_110111101101;
      patterns[23516] = 29'b0_101101111011_100_1_010110111101;
      patterns[23517] = 29'b0_101101111011_101_1_101011011110;
      patterns[23518] = 29'b0_101101111011_110_0_101101111011;
      patterns[23519] = 29'b0_101101111011_111_0_101101111011;
      patterns[23520] = 29'b0_101101111100_000_0_101101111100;
      patterns[23521] = 29'b0_101101111100_001_0_111100101101;
      patterns[23522] = 29'b0_101101111100_010_1_011011111000;
      patterns[23523] = 29'b0_101101111100_011_0_110111110001;
      patterns[23524] = 29'b0_101101111100_100_0_010110111110;
      patterns[23525] = 29'b0_101101111100_101_0_001011011111;
      patterns[23526] = 29'b0_101101111100_110_0_101101111100;
      patterns[23527] = 29'b0_101101111100_111_0_101101111100;
      patterns[23528] = 29'b0_101101111101_000_0_101101111101;
      patterns[23529] = 29'b0_101101111101_001_0_111101101101;
      patterns[23530] = 29'b0_101101111101_010_1_011011111010;
      patterns[23531] = 29'b0_101101111101_011_0_110111110101;
      patterns[23532] = 29'b0_101101111101_100_1_010110111110;
      patterns[23533] = 29'b0_101101111101_101_0_101011011111;
      patterns[23534] = 29'b0_101101111101_110_0_101101111101;
      patterns[23535] = 29'b0_101101111101_111_0_101101111101;
      patterns[23536] = 29'b0_101101111110_000_0_101101111110;
      patterns[23537] = 29'b0_101101111110_001_0_111110101101;
      patterns[23538] = 29'b0_101101111110_010_1_011011111100;
      patterns[23539] = 29'b0_101101111110_011_0_110111111001;
      patterns[23540] = 29'b0_101101111110_100_0_010110111111;
      patterns[23541] = 29'b0_101101111110_101_1_001011011111;
      patterns[23542] = 29'b0_101101111110_110_0_101101111110;
      patterns[23543] = 29'b0_101101111110_111_0_101101111110;
      patterns[23544] = 29'b0_101101111111_000_0_101101111111;
      patterns[23545] = 29'b0_101101111111_001_0_111111101101;
      patterns[23546] = 29'b0_101101111111_010_1_011011111110;
      patterns[23547] = 29'b0_101101111111_011_0_110111111101;
      patterns[23548] = 29'b0_101101111111_100_1_010110111111;
      patterns[23549] = 29'b0_101101111111_101_1_101011011111;
      patterns[23550] = 29'b0_101101111111_110_0_101101111111;
      patterns[23551] = 29'b0_101101111111_111_0_101101111111;
      patterns[23552] = 29'b0_101110000000_000_0_101110000000;
      patterns[23553] = 29'b0_101110000000_001_0_000000101110;
      patterns[23554] = 29'b0_101110000000_010_1_011100000000;
      patterns[23555] = 29'b0_101110000000_011_0_111000000001;
      patterns[23556] = 29'b0_101110000000_100_0_010111000000;
      patterns[23557] = 29'b0_101110000000_101_0_001011100000;
      patterns[23558] = 29'b0_101110000000_110_0_101110000000;
      patterns[23559] = 29'b0_101110000000_111_0_101110000000;
      patterns[23560] = 29'b0_101110000001_000_0_101110000001;
      patterns[23561] = 29'b0_101110000001_001_0_000001101110;
      patterns[23562] = 29'b0_101110000001_010_1_011100000010;
      patterns[23563] = 29'b0_101110000001_011_0_111000000101;
      patterns[23564] = 29'b0_101110000001_100_1_010111000000;
      patterns[23565] = 29'b0_101110000001_101_0_101011100000;
      patterns[23566] = 29'b0_101110000001_110_0_101110000001;
      patterns[23567] = 29'b0_101110000001_111_0_101110000001;
      patterns[23568] = 29'b0_101110000010_000_0_101110000010;
      patterns[23569] = 29'b0_101110000010_001_0_000010101110;
      patterns[23570] = 29'b0_101110000010_010_1_011100000100;
      patterns[23571] = 29'b0_101110000010_011_0_111000001001;
      patterns[23572] = 29'b0_101110000010_100_0_010111000001;
      patterns[23573] = 29'b0_101110000010_101_1_001011100000;
      patterns[23574] = 29'b0_101110000010_110_0_101110000010;
      patterns[23575] = 29'b0_101110000010_111_0_101110000010;
      patterns[23576] = 29'b0_101110000011_000_0_101110000011;
      patterns[23577] = 29'b0_101110000011_001_0_000011101110;
      patterns[23578] = 29'b0_101110000011_010_1_011100000110;
      patterns[23579] = 29'b0_101110000011_011_0_111000001101;
      patterns[23580] = 29'b0_101110000011_100_1_010111000001;
      patterns[23581] = 29'b0_101110000011_101_1_101011100000;
      patterns[23582] = 29'b0_101110000011_110_0_101110000011;
      patterns[23583] = 29'b0_101110000011_111_0_101110000011;
      patterns[23584] = 29'b0_101110000100_000_0_101110000100;
      patterns[23585] = 29'b0_101110000100_001_0_000100101110;
      patterns[23586] = 29'b0_101110000100_010_1_011100001000;
      patterns[23587] = 29'b0_101110000100_011_0_111000010001;
      patterns[23588] = 29'b0_101110000100_100_0_010111000010;
      patterns[23589] = 29'b0_101110000100_101_0_001011100001;
      patterns[23590] = 29'b0_101110000100_110_0_101110000100;
      patterns[23591] = 29'b0_101110000100_111_0_101110000100;
      patterns[23592] = 29'b0_101110000101_000_0_101110000101;
      patterns[23593] = 29'b0_101110000101_001_0_000101101110;
      patterns[23594] = 29'b0_101110000101_010_1_011100001010;
      patterns[23595] = 29'b0_101110000101_011_0_111000010101;
      patterns[23596] = 29'b0_101110000101_100_1_010111000010;
      patterns[23597] = 29'b0_101110000101_101_0_101011100001;
      patterns[23598] = 29'b0_101110000101_110_0_101110000101;
      patterns[23599] = 29'b0_101110000101_111_0_101110000101;
      patterns[23600] = 29'b0_101110000110_000_0_101110000110;
      patterns[23601] = 29'b0_101110000110_001_0_000110101110;
      patterns[23602] = 29'b0_101110000110_010_1_011100001100;
      patterns[23603] = 29'b0_101110000110_011_0_111000011001;
      patterns[23604] = 29'b0_101110000110_100_0_010111000011;
      patterns[23605] = 29'b0_101110000110_101_1_001011100001;
      patterns[23606] = 29'b0_101110000110_110_0_101110000110;
      patterns[23607] = 29'b0_101110000110_111_0_101110000110;
      patterns[23608] = 29'b0_101110000111_000_0_101110000111;
      patterns[23609] = 29'b0_101110000111_001_0_000111101110;
      patterns[23610] = 29'b0_101110000111_010_1_011100001110;
      patterns[23611] = 29'b0_101110000111_011_0_111000011101;
      patterns[23612] = 29'b0_101110000111_100_1_010111000011;
      patterns[23613] = 29'b0_101110000111_101_1_101011100001;
      patterns[23614] = 29'b0_101110000111_110_0_101110000111;
      patterns[23615] = 29'b0_101110000111_111_0_101110000111;
      patterns[23616] = 29'b0_101110001000_000_0_101110001000;
      patterns[23617] = 29'b0_101110001000_001_0_001000101110;
      patterns[23618] = 29'b0_101110001000_010_1_011100010000;
      patterns[23619] = 29'b0_101110001000_011_0_111000100001;
      patterns[23620] = 29'b0_101110001000_100_0_010111000100;
      patterns[23621] = 29'b0_101110001000_101_0_001011100010;
      patterns[23622] = 29'b0_101110001000_110_0_101110001000;
      patterns[23623] = 29'b0_101110001000_111_0_101110001000;
      patterns[23624] = 29'b0_101110001001_000_0_101110001001;
      patterns[23625] = 29'b0_101110001001_001_0_001001101110;
      patterns[23626] = 29'b0_101110001001_010_1_011100010010;
      patterns[23627] = 29'b0_101110001001_011_0_111000100101;
      patterns[23628] = 29'b0_101110001001_100_1_010111000100;
      patterns[23629] = 29'b0_101110001001_101_0_101011100010;
      patterns[23630] = 29'b0_101110001001_110_0_101110001001;
      patterns[23631] = 29'b0_101110001001_111_0_101110001001;
      patterns[23632] = 29'b0_101110001010_000_0_101110001010;
      patterns[23633] = 29'b0_101110001010_001_0_001010101110;
      patterns[23634] = 29'b0_101110001010_010_1_011100010100;
      patterns[23635] = 29'b0_101110001010_011_0_111000101001;
      patterns[23636] = 29'b0_101110001010_100_0_010111000101;
      patterns[23637] = 29'b0_101110001010_101_1_001011100010;
      patterns[23638] = 29'b0_101110001010_110_0_101110001010;
      patterns[23639] = 29'b0_101110001010_111_0_101110001010;
      patterns[23640] = 29'b0_101110001011_000_0_101110001011;
      patterns[23641] = 29'b0_101110001011_001_0_001011101110;
      patterns[23642] = 29'b0_101110001011_010_1_011100010110;
      patterns[23643] = 29'b0_101110001011_011_0_111000101101;
      patterns[23644] = 29'b0_101110001011_100_1_010111000101;
      patterns[23645] = 29'b0_101110001011_101_1_101011100010;
      patterns[23646] = 29'b0_101110001011_110_0_101110001011;
      patterns[23647] = 29'b0_101110001011_111_0_101110001011;
      patterns[23648] = 29'b0_101110001100_000_0_101110001100;
      patterns[23649] = 29'b0_101110001100_001_0_001100101110;
      patterns[23650] = 29'b0_101110001100_010_1_011100011000;
      patterns[23651] = 29'b0_101110001100_011_0_111000110001;
      patterns[23652] = 29'b0_101110001100_100_0_010111000110;
      patterns[23653] = 29'b0_101110001100_101_0_001011100011;
      patterns[23654] = 29'b0_101110001100_110_0_101110001100;
      patterns[23655] = 29'b0_101110001100_111_0_101110001100;
      patterns[23656] = 29'b0_101110001101_000_0_101110001101;
      patterns[23657] = 29'b0_101110001101_001_0_001101101110;
      patterns[23658] = 29'b0_101110001101_010_1_011100011010;
      patterns[23659] = 29'b0_101110001101_011_0_111000110101;
      patterns[23660] = 29'b0_101110001101_100_1_010111000110;
      patterns[23661] = 29'b0_101110001101_101_0_101011100011;
      patterns[23662] = 29'b0_101110001101_110_0_101110001101;
      patterns[23663] = 29'b0_101110001101_111_0_101110001101;
      patterns[23664] = 29'b0_101110001110_000_0_101110001110;
      patterns[23665] = 29'b0_101110001110_001_0_001110101110;
      patterns[23666] = 29'b0_101110001110_010_1_011100011100;
      patterns[23667] = 29'b0_101110001110_011_0_111000111001;
      patterns[23668] = 29'b0_101110001110_100_0_010111000111;
      patterns[23669] = 29'b0_101110001110_101_1_001011100011;
      patterns[23670] = 29'b0_101110001110_110_0_101110001110;
      patterns[23671] = 29'b0_101110001110_111_0_101110001110;
      patterns[23672] = 29'b0_101110001111_000_0_101110001111;
      patterns[23673] = 29'b0_101110001111_001_0_001111101110;
      patterns[23674] = 29'b0_101110001111_010_1_011100011110;
      patterns[23675] = 29'b0_101110001111_011_0_111000111101;
      patterns[23676] = 29'b0_101110001111_100_1_010111000111;
      patterns[23677] = 29'b0_101110001111_101_1_101011100011;
      patterns[23678] = 29'b0_101110001111_110_0_101110001111;
      patterns[23679] = 29'b0_101110001111_111_0_101110001111;
      patterns[23680] = 29'b0_101110010000_000_0_101110010000;
      patterns[23681] = 29'b0_101110010000_001_0_010000101110;
      patterns[23682] = 29'b0_101110010000_010_1_011100100000;
      patterns[23683] = 29'b0_101110010000_011_0_111001000001;
      patterns[23684] = 29'b0_101110010000_100_0_010111001000;
      patterns[23685] = 29'b0_101110010000_101_0_001011100100;
      patterns[23686] = 29'b0_101110010000_110_0_101110010000;
      patterns[23687] = 29'b0_101110010000_111_0_101110010000;
      patterns[23688] = 29'b0_101110010001_000_0_101110010001;
      patterns[23689] = 29'b0_101110010001_001_0_010001101110;
      patterns[23690] = 29'b0_101110010001_010_1_011100100010;
      patterns[23691] = 29'b0_101110010001_011_0_111001000101;
      patterns[23692] = 29'b0_101110010001_100_1_010111001000;
      patterns[23693] = 29'b0_101110010001_101_0_101011100100;
      patterns[23694] = 29'b0_101110010001_110_0_101110010001;
      patterns[23695] = 29'b0_101110010001_111_0_101110010001;
      patterns[23696] = 29'b0_101110010010_000_0_101110010010;
      patterns[23697] = 29'b0_101110010010_001_0_010010101110;
      patterns[23698] = 29'b0_101110010010_010_1_011100100100;
      patterns[23699] = 29'b0_101110010010_011_0_111001001001;
      patterns[23700] = 29'b0_101110010010_100_0_010111001001;
      patterns[23701] = 29'b0_101110010010_101_1_001011100100;
      patterns[23702] = 29'b0_101110010010_110_0_101110010010;
      patterns[23703] = 29'b0_101110010010_111_0_101110010010;
      patterns[23704] = 29'b0_101110010011_000_0_101110010011;
      patterns[23705] = 29'b0_101110010011_001_0_010011101110;
      patterns[23706] = 29'b0_101110010011_010_1_011100100110;
      patterns[23707] = 29'b0_101110010011_011_0_111001001101;
      patterns[23708] = 29'b0_101110010011_100_1_010111001001;
      patterns[23709] = 29'b0_101110010011_101_1_101011100100;
      patterns[23710] = 29'b0_101110010011_110_0_101110010011;
      patterns[23711] = 29'b0_101110010011_111_0_101110010011;
      patterns[23712] = 29'b0_101110010100_000_0_101110010100;
      patterns[23713] = 29'b0_101110010100_001_0_010100101110;
      patterns[23714] = 29'b0_101110010100_010_1_011100101000;
      patterns[23715] = 29'b0_101110010100_011_0_111001010001;
      patterns[23716] = 29'b0_101110010100_100_0_010111001010;
      patterns[23717] = 29'b0_101110010100_101_0_001011100101;
      patterns[23718] = 29'b0_101110010100_110_0_101110010100;
      patterns[23719] = 29'b0_101110010100_111_0_101110010100;
      patterns[23720] = 29'b0_101110010101_000_0_101110010101;
      patterns[23721] = 29'b0_101110010101_001_0_010101101110;
      patterns[23722] = 29'b0_101110010101_010_1_011100101010;
      patterns[23723] = 29'b0_101110010101_011_0_111001010101;
      patterns[23724] = 29'b0_101110010101_100_1_010111001010;
      patterns[23725] = 29'b0_101110010101_101_0_101011100101;
      patterns[23726] = 29'b0_101110010101_110_0_101110010101;
      patterns[23727] = 29'b0_101110010101_111_0_101110010101;
      patterns[23728] = 29'b0_101110010110_000_0_101110010110;
      patterns[23729] = 29'b0_101110010110_001_0_010110101110;
      patterns[23730] = 29'b0_101110010110_010_1_011100101100;
      patterns[23731] = 29'b0_101110010110_011_0_111001011001;
      patterns[23732] = 29'b0_101110010110_100_0_010111001011;
      patterns[23733] = 29'b0_101110010110_101_1_001011100101;
      patterns[23734] = 29'b0_101110010110_110_0_101110010110;
      patterns[23735] = 29'b0_101110010110_111_0_101110010110;
      patterns[23736] = 29'b0_101110010111_000_0_101110010111;
      patterns[23737] = 29'b0_101110010111_001_0_010111101110;
      patterns[23738] = 29'b0_101110010111_010_1_011100101110;
      patterns[23739] = 29'b0_101110010111_011_0_111001011101;
      patterns[23740] = 29'b0_101110010111_100_1_010111001011;
      patterns[23741] = 29'b0_101110010111_101_1_101011100101;
      patterns[23742] = 29'b0_101110010111_110_0_101110010111;
      patterns[23743] = 29'b0_101110010111_111_0_101110010111;
      patterns[23744] = 29'b0_101110011000_000_0_101110011000;
      patterns[23745] = 29'b0_101110011000_001_0_011000101110;
      patterns[23746] = 29'b0_101110011000_010_1_011100110000;
      patterns[23747] = 29'b0_101110011000_011_0_111001100001;
      patterns[23748] = 29'b0_101110011000_100_0_010111001100;
      patterns[23749] = 29'b0_101110011000_101_0_001011100110;
      patterns[23750] = 29'b0_101110011000_110_0_101110011000;
      patterns[23751] = 29'b0_101110011000_111_0_101110011000;
      patterns[23752] = 29'b0_101110011001_000_0_101110011001;
      patterns[23753] = 29'b0_101110011001_001_0_011001101110;
      patterns[23754] = 29'b0_101110011001_010_1_011100110010;
      patterns[23755] = 29'b0_101110011001_011_0_111001100101;
      patterns[23756] = 29'b0_101110011001_100_1_010111001100;
      patterns[23757] = 29'b0_101110011001_101_0_101011100110;
      patterns[23758] = 29'b0_101110011001_110_0_101110011001;
      patterns[23759] = 29'b0_101110011001_111_0_101110011001;
      patterns[23760] = 29'b0_101110011010_000_0_101110011010;
      patterns[23761] = 29'b0_101110011010_001_0_011010101110;
      patterns[23762] = 29'b0_101110011010_010_1_011100110100;
      patterns[23763] = 29'b0_101110011010_011_0_111001101001;
      patterns[23764] = 29'b0_101110011010_100_0_010111001101;
      patterns[23765] = 29'b0_101110011010_101_1_001011100110;
      patterns[23766] = 29'b0_101110011010_110_0_101110011010;
      patterns[23767] = 29'b0_101110011010_111_0_101110011010;
      patterns[23768] = 29'b0_101110011011_000_0_101110011011;
      patterns[23769] = 29'b0_101110011011_001_0_011011101110;
      patterns[23770] = 29'b0_101110011011_010_1_011100110110;
      patterns[23771] = 29'b0_101110011011_011_0_111001101101;
      patterns[23772] = 29'b0_101110011011_100_1_010111001101;
      patterns[23773] = 29'b0_101110011011_101_1_101011100110;
      patterns[23774] = 29'b0_101110011011_110_0_101110011011;
      patterns[23775] = 29'b0_101110011011_111_0_101110011011;
      patterns[23776] = 29'b0_101110011100_000_0_101110011100;
      patterns[23777] = 29'b0_101110011100_001_0_011100101110;
      patterns[23778] = 29'b0_101110011100_010_1_011100111000;
      patterns[23779] = 29'b0_101110011100_011_0_111001110001;
      patterns[23780] = 29'b0_101110011100_100_0_010111001110;
      patterns[23781] = 29'b0_101110011100_101_0_001011100111;
      patterns[23782] = 29'b0_101110011100_110_0_101110011100;
      patterns[23783] = 29'b0_101110011100_111_0_101110011100;
      patterns[23784] = 29'b0_101110011101_000_0_101110011101;
      patterns[23785] = 29'b0_101110011101_001_0_011101101110;
      patterns[23786] = 29'b0_101110011101_010_1_011100111010;
      patterns[23787] = 29'b0_101110011101_011_0_111001110101;
      patterns[23788] = 29'b0_101110011101_100_1_010111001110;
      patterns[23789] = 29'b0_101110011101_101_0_101011100111;
      patterns[23790] = 29'b0_101110011101_110_0_101110011101;
      patterns[23791] = 29'b0_101110011101_111_0_101110011101;
      patterns[23792] = 29'b0_101110011110_000_0_101110011110;
      patterns[23793] = 29'b0_101110011110_001_0_011110101110;
      patterns[23794] = 29'b0_101110011110_010_1_011100111100;
      patterns[23795] = 29'b0_101110011110_011_0_111001111001;
      patterns[23796] = 29'b0_101110011110_100_0_010111001111;
      patterns[23797] = 29'b0_101110011110_101_1_001011100111;
      patterns[23798] = 29'b0_101110011110_110_0_101110011110;
      patterns[23799] = 29'b0_101110011110_111_0_101110011110;
      patterns[23800] = 29'b0_101110011111_000_0_101110011111;
      patterns[23801] = 29'b0_101110011111_001_0_011111101110;
      patterns[23802] = 29'b0_101110011111_010_1_011100111110;
      patterns[23803] = 29'b0_101110011111_011_0_111001111101;
      patterns[23804] = 29'b0_101110011111_100_1_010111001111;
      patterns[23805] = 29'b0_101110011111_101_1_101011100111;
      patterns[23806] = 29'b0_101110011111_110_0_101110011111;
      patterns[23807] = 29'b0_101110011111_111_0_101110011111;
      patterns[23808] = 29'b0_101110100000_000_0_101110100000;
      patterns[23809] = 29'b0_101110100000_001_0_100000101110;
      patterns[23810] = 29'b0_101110100000_010_1_011101000000;
      patterns[23811] = 29'b0_101110100000_011_0_111010000001;
      patterns[23812] = 29'b0_101110100000_100_0_010111010000;
      patterns[23813] = 29'b0_101110100000_101_0_001011101000;
      patterns[23814] = 29'b0_101110100000_110_0_101110100000;
      patterns[23815] = 29'b0_101110100000_111_0_101110100000;
      patterns[23816] = 29'b0_101110100001_000_0_101110100001;
      patterns[23817] = 29'b0_101110100001_001_0_100001101110;
      patterns[23818] = 29'b0_101110100001_010_1_011101000010;
      patterns[23819] = 29'b0_101110100001_011_0_111010000101;
      patterns[23820] = 29'b0_101110100001_100_1_010111010000;
      patterns[23821] = 29'b0_101110100001_101_0_101011101000;
      patterns[23822] = 29'b0_101110100001_110_0_101110100001;
      patterns[23823] = 29'b0_101110100001_111_0_101110100001;
      patterns[23824] = 29'b0_101110100010_000_0_101110100010;
      patterns[23825] = 29'b0_101110100010_001_0_100010101110;
      patterns[23826] = 29'b0_101110100010_010_1_011101000100;
      patterns[23827] = 29'b0_101110100010_011_0_111010001001;
      patterns[23828] = 29'b0_101110100010_100_0_010111010001;
      patterns[23829] = 29'b0_101110100010_101_1_001011101000;
      patterns[23830] = 29'b0_101110100010_110_0_101110100010;
      patterns[23831] = 29'b0_101110100010_111_0_101110100010;
      patterns[23832] = 29'b0_101110100011_000_0_101110100011;
      patterns[23833] = 29'b0_101110100011_001_0_100011101110;
      patterns[23834] = 29'b0_101110100011_010_1_011101000110;
      patterns[23835] = 29'b0_101110100011_011_0_111010001101;
      patterns[23836] = 29'b0_101110100011_100_1_010111010001;
      patterns[23837] = 29'b0_101110100011_101_1_101011101000;
      patterns[23838] = 29'b0_101110100011_110_0_101110100011;
      patterns[23839] = 29'b0_101110100011_111_0_101110100011;
      patterns[23840] = 29'b0_101110100100_000_0_101110100100;
      patterns[23841] = 29'b0_101110100100_001_0_100100101110;
      patterns[23842] = 29'b0_101110100100_010_1_011101001000;
      patterns[23843] = 29'b0_101110100100_011_0_111010010001;
      patterns[23844] = 29'b0_101110100100_100_0_010111010010;
      patterns[23845] = 29'b0_101110100100_101_0_001011101001;
      patterns[23846] = 29'b0_101110100100_110_0_101110100100;
      patterns[23847] = 29'b0_101110100100_111_0_101110100100;
      patterns[23848] = 29'b0_101110100101_000_0_101110100101;
      patterns[23849] = 29'b0_101110100101_001_0_100101101110;
      patterns[23850] = 29'b0_101110100101_010_1_011101001010;
      patterns[23851] = 29'b0_101110100101_011_0_111010010101;
      patterns[23852] = 29'b0_101110100101_100_1_010111010010;
      patterns[23853] = 29'b0_101110100101_101_0_101011101001;
      patterns[23854] = 29'b0_101110100101_110_0_101110100101;
      patterns[23855] = 29'b0_101110100101_111_0_101110100101;
      patterns[23856] = 29'b0_101110100110_000_0_101110100110;
      patterns[23857] = 29'b0_101110100110_001_0_100110101110;
      patterns[23858] = 29'b0_101110100110_010_1_011101001100;
      patterns[23859] = 29'b0_101110100110_011_0_111010011001;
      patterns[23860] = 29'b0_101110100110_100_0_010111010011;
      patterns[23861] = 29'b0_101110100110_101_1_001011101001;
      patterns[23862] = 29'b0_101110100110_110_0_101110100110;
      patterns[23863] = 29'b0_101110100110_111_0_101110100110;
      patterns[23864] = 29'b0_101110100111_000_0_101110100111;
      patterns[23865] = 29'b0_101110100111_001_0_100111101110;
      patterns[23866] = 29'b0_101110100111_010_1_011101001110;
      patterns[23867] = 29'b0_101110100111_011_0_111010011101;
      patterns[23868] = 29'b0_101110100111_100_1_010111010011;
      patterns[23869] = 29'b0_101110100111_101_1_101011101001;
      patterns[23870] = 29'b0_101110100111_110_0_101110100111;
      patterns[23871] = 29'b0_101110100111_111_0_101110100111;
      patterns[23872] = 29'b0_101110101000_000_0_101110101000;
      patterns[23873] = 29'b0_101110101000_001_0_101000101110;
      patterns[23874] = 29'b0_101110101000_010_1_011101010000;
      patterns[23875] = 29'b0_101110101000_011_0_111010100001;
      patterns[23876] = 29'b0_101110101000_100_0_010111010100;
      patterns[23877] = 29'b0_101110101000_101_0_001011101010;
      patterns[23878] = 29'b0_101110101000_110_0_101110101000;
      patterns[23879] = 29'b0_101110101000_111_0_101110101000;
      patterns[23880] = 29'b0_101110101001_000_0_101110101001;
      patterns[23881] = 29'b0_101110101001_001_0_101001101110;
      patterns[23882] = 29'b0_101110101001_010_1_011101010010;
      patterns[23883] = 29'b0_101110101001_011_0_111010100101;
      patterns[23884] = 29'b0_101110101001_100_1_010111010100;
      patterns[23885] = 29'b0_101110101001_101_0_101011101010;
      patterns[23886] = 29'b0_101110101001_110_0_101110101001;
      patterns[23887] = 29'b0_101110101001_111_0_101110101001;
      patterns[23888] = 29'b0_101110101010_000_0_101110101010;
      patterns[23889] = 29'b0_101110101010_001_0_101010101110;
      patterns[23890] = 29'b0_101110101010_010_1_011101010100;
      patterns[23891] = 29'b0_101110101010_011_0_111010101001;
      patterns[23892] = 29'b0_101110101010_100_0_010111010101;
      patterns[23893] = 29'b0_101110101010_101_1_001011101010;
      patterns[23894] = 29'b0_101110101010_110_0_101110101010;
      patterns[23895] = 29'b0_101110101010_111_0_101110101010;
      patterns[23896] = 29'b0_101110101011_000_0_101110101011;
      patterns[23897] = 29'b0_101110101011_001_0_101011101110;
      patterns[23898] = 29'b0_101110101011_010_1_011101010110;
      patterns[23899] = 29'b0_101110101011_011_0_111010101101;
      patterns[23900] = 29'b0_101110101011_100_1_010111010101;
      patterns[23901] = 29'b0_101110101011_101_1_101011101010;
      patterns[23902] = 29'b0_101110101011_110_0_101110101011;
      patterns[23903] = 29'b0_101110101011_111_0_101110101011;
      patterns[23904] = 29'b0_101110101100_000_0_101110101100;
      patterns[23905] = 29'b0_101110101100_001_0_101100101110;
      patterns[23906] = 29'b0_101110101100_010_1_011101011000;
      patterns[23907] = 29'b0_101110101100_011_0_111010110001;
      patterns[23908] = 29'b0_101110101100_100_0_010111010110;
      patterns[23909] = 29'b0_101110101100_101_0_001011101011;
      patterns[23910] = 29'b0_101110101100_110_0_101110101100;
      patterns[23911] = 29'b0_101110101100_111_0_101110101100;
      patterns[23912] = 29'b0_101110101101_000_0_101110101101;
      patterns[23913] = 29'b0_101110101101_001_0_101101101110;
      patterns[23914] = 29'b0_101110101101_010_1_011101011010;
      patterns[23915] = 29'b0_101110101101_011_0_111010110101;
      patterns[23916] = 29'b0_101110101101_100_1_010111010110;
      patterns[23917] = 29'b0_101110101101_101_0_101011101011;
      patterns[23918] = 29'b0_101110101101_110_0_101110101101;
      patterns[23919] = 29'b0_101110101101_111_0_101110101101;
      patterns[23920] = 29'b0_101110101110_000_0_101110101110;
      patterns[23921] = 29'b0_101110101110_001_0_101110101110;
      patterns[23922] = 29'b0_101110101110_010_1_011101011100;
      patterns[23923] = 29'b0_101110101110_011_0_111010111001;
      patterns[23924] = 29'b0_101110101110_100_0_010111010111;
      patterns[23925] = 29'b0_101110101110_101_1_001011101011;
      patterns[23926] = 29'b0_101110101110_110_0_101110101110;
      patterns[23927] = 29'b0_101110101110_111_0_101110101110;
      patterns[23928] = 29'b0_101110101111_000_0_101110101111;
      patterns[23929] = 29'b0_101110101111_001_0_101111101110;
      patterns[23930] = 29'b0_101110101111_010_1_011101011110;
      patterns[23931] = 29'b0_101110101111_011_0_111010111101;
      patterns[23932] = 29'b0_101110101111_100_1_010111010111;
      patterns[23933] = 29'b0_101110101111_101_1_101011101011;
      patterns[23934] = 29'b0_101110101111_110_0_101110101111;
      patterns[23935] = 29'b0_101110101111_111_0_101110101111;
      patterns[23936] = 29'b0_101110110000_000_0_101110110000;
      patterns[23937] = 29'b0_101110110000_001_0_110000101110;
      patterns[23938] = 29'b0_101110110000_010_1_011101100000;
      patterns[23939] = 29'b0_101110110000_011_0_111011000001;
      patterns[23940] = 29'b0_101110110000_100_0_010111011000;
      patterns[23941] = 29'b0_101110110000_101_0_001011101100;
      patterns[23942] = 29'b0_101110110000_110_0_101110110000;
      patterns[23943] = 29'b0_101110110000_111_0_101110110000;
      patterns[23944] = 29'b0_101110110001_000_0_101110110001;
      patterns[23945] = 29'b0_101110110001_001_0_110001101110;
      patterns[23946] = 29'b0_101110110001_010_1_011101100010;
      patterns[23947] = 29'b0_101110110001_011_0_111011000101;
      patterns[23948] = 29'b0_101110110001_100_1_010111011000;
      patterns[23949] = 29'b0_101110110001_101_0_101011101100;
      patterns[23950] = 29'b0_101110110001_110_0_101110110001;
      patterns[23951] = 29'b0_101110110001_111_0_101110110001;
      patterns[23952] = 29'b0_101110110010_000_0_101110110010;
      patterns[23953] = 29'b0_101110110010_001_0_110010101110;
      patterns[23954] = 29'b0_101110110010_010_1_011101100100;
      patterns[23955] = 29'b0_101110110010_011_0_111011001001;
      patterns[23956] = 29'b0_101110110010_100_0_010111011001;
      patterns[23957] = 29'b0_101110110010_101_1_001011101100;
      patterns[23958] = 29'b0_101110110010_110_0_101110110010;
      patterns[23959] = 29'b0_101110110010_111_0_101110110010;
      patterns[23960] = 29'b0_101110110011_000_0_101110110011;
      patterns[23961] = 29'b0_101110110011_001_0_110011101110;
      patterns[23962] = 29'b0_101110110011_010_1_011101100110;
      patterns[23963] = 29'b0_101110110011_011_0_111011001101;
      patterns[23964] = 29'b0_101110110011_100_1_010111011001;
      patterns[23965] = 29'b0_101110110011_101_1_101011101100;
      patterns[23966] = 29'b0_101110110011_110_0_101110110011;
      patterns[23967] = 29'b0_101110110011_111_0_101110110011;
      patterns[23968] = 29'b0_101110110100_000_0_101110110100;
      patterns[23969] = 29'b0_101110110100_001_0_110100101110;
      patterns[23970] = 29'b0_101110110100_010_1_011101101000;
      patterns[23971] = 29'b0_101110110100_011_0_111011010001;
      patterns[23972] = 29'b0_101110110100_100_0_010111011010;
      patterns[23973] = 29'b0_101110110100_101_0_001011101101;
      patterns[23974] = 29'b0_101110110100_110_0_101110110100;
      patterns[23975] = 29'b0_101110110100_111_0_101110110100;
      patterns[23976] = 29'b0_101110110101_000_0_101110110101;
      patterns[23977] = 29'b0_101110110101_001_0_110101101110;
      patterns[23978] = 29'b0_101110110101_010_1_011101101010;
      patterns[23979] = 29'b0_101110110101_011_0_111011010101;
      patterns[23980] = 29'b0_101110110101_100_1_010111011010;
      patterns[23981] = 29'b0_101110110101_101_0_101011101101;
      patterns[23982] = 29'b0_101110110101_110_0_101110110101;
      patterns[23983] = 29'b0_101110110101_111_0_101110110101;
      patterns[23984] = 29'b0_101110110110_000_0_101110110110;
      patterns[23985] = 29'b0_101110110110_001_0_110110101110;
      patterns[23986] = 29'b0_101110110110_010_1_011101101100;
      patterns[23987] = 29'b0_101110110110_011_0_111011011001;
      patterns[23988] = 29'b0_101110110110_100_0_010111011011;
      patterns[23989] = 29'b0_101110110110_101_1_001011101101;
      patterns[23990] = 29'b0_101110110110_110_0_101110110110;
      patterns[23991] = 29'b0_101110110110_111_0_101110110110;
      patterns[23992] = 29'b0_101110110111_000_0_101110110111;
      patterns[23993] = 29'b0_101110110111_001_0_110111101110;
      patterns[23994] = 29'b0_101110110111_010_1_011101101110;
      patterns[23995] = 29'b0_101110110111_011_0_111011011101;
      patterns[23996] = 29'b0_101110110111_100_1_010111011011;
      patterns[23997] = 29'b0_101110110111_101_1_101011101101;
      patterns[23998] = 29'b0_101110110111_110_0_101110110111;
      patterns[23999] = 29'b0_101110110111_111_0_101110110111;
      patterns[24000] = 29'b0_101110111000_000_0_101110111000;
      patterns[24001] = 29'b0_101110111000_001_0_111000101110;
      patterns[24002] = 29'b0_101110111000_010_1_011101110000;
      patterns[24003] = 29'b0_101110111000_011_0_111011100001;
      patterns[24004] = 29'b0_101110111000_100_0_010111011100;
      patterns[24005] = 29'b0_101110111000_101_0_001011101110;
      patterns[24006] = 29'b0_101110111000_110_0_101110111000;
      patterns[24007] = 29'b0_101110111000_111_0_101110111000;
      patterns[24008] = 29'b0_101110111001_000_0_101110111001;
      patterns[24009] = 29'b0_101110111001_001_0_111001101110;
      patterns[24010] = 29'b0_101110111001_010_1_011101110010;
      patterns[24011] = 29'b0_101110111001_011_0_111011100101;
      patterns[24012] = 29'b0_101110111001_100_1_010111011100;
      patterns[24013] = 29'b0_101110111001_101_0_101011101110;
      patterns[24014] = 29'b0_101110111001_110_0_101110111001;
      patterns[24015] = 29'b0_101110111001_111_0_101110111001;
      patterns[24016] = 29'b0_101110111010_000_0_101110111010;
      patterns[24017] = 29'b0_101110111010_001_0_111010101110;
      patterns[24018] = 29'b0_101110111010_010_1_011101110100;
      patterns[24019] = 29'b0_101110111010_011_0_111011101001;
      patterns[24020] = 29'b0_101110111010_100_0_010111011101;
      patterns[24021] = 29'b0_101110111010_101_1_001011101110;
      patterns[24022] = 29'b0_101110111010_110_0_101110111010;
      patterns[24023] = 29'b0_101110111010_111_0_101110111010;
      patterns[24024] = 29'b0_101110111011_000_0_101110111011;
      patterns[24025] = 29'b0_101110111011_001_0_111011101110;
      patterns[24026] = 29'b0_101110111011_010_1_011101110110;
      patterns[24027] = 29'b0_101110111011_011_0_111011101101;
      patterns[24028] = 29'b0_101110111011_100_1_010111011101;
      patterns[24029] = 29'b0_101110111011_101_1_101011101110;
      patterns[24030] = 29'b0_101110111011_110_0_101110111011;
      patterns[24031] = 29'b0_101110111011_111_0_101110111011;
      patterns[24032] = 29'b0_101110111100_000_0_101110111100;
      patterns[24033] = 29'b0_101110111100_001_0_111100101110;
      patterns[24034] = 29'b0_101110111100_010_1_011101111000;
      patterns[24035] = 29'b0_101110111100_011_0_111011110001;
      patterns[24036] = 29'b0_101110111100_100_0_010111011110;
      patterns[24037] = 29'b0_101110111100_101_0_001011101111;
      patterns[24038] = 29'b0_101110111100_110_0_101110111100;
      patterns[24039] = 29'b0_101110111100_111_0_101110111100;
      patterns[24040] = 29'b0_101110111101_000_0_101110111101;
      patterns[24041] = 29'b0_101110111101_001_0_111101101110;
      patterns[24042] = 29'b0_101110111101_010_1_011101111010;
      patterns[24043] = 29'b0_101110111101_011_0_111011110101;
      patterns[24044] = 29'b0_101110111101_100_1_010111011110;
      patterns[24045] = 29'b0_101110111101_101_0_101011101111;
      patterns[24046] = 29'b0_101110111101_110_0_101110111101;
      patterns[24047] = 29'b0_101110111101_111_0_101110111101;
      patterns[24048] = 29'b0_101110111110_000_0_101110111110;
      patterns[24049] = 29'b0_101110111110_001_0_111110101110;
      patterns[24050] = 29'b0_101110111110_010_1_011101111100;
      patterns[24051] = 29'b0_101110111110_011_0_111011111001;
      patterns[24052] = 29'b0_101110111110_100_0_010111011111;
      patterns[24053] = 29'b0_101110111110_101_1_001011101111;
      patterns[24054] = 29'b0_101110111110_110_0_101110111110;
      patterns[24055] = 29'b0_101110111110_111_0_101110111110;
      patterns[24056] = 29'b0_101110111111_000_0_101110111111;
      patterns[24057] = 29'b0_101110111111_001_0_111111101110;
      patterns[24058] = 29'b0_101110111111_010_1_011101111110;
      patterns[24059] = 29'b0_101110111111_011_0_111011111101;
      patterns[24060] = 29'b0_101110111111_100_1_010111011111;
      patterns[24061] = 29'b0_101110111111_101_1_101011101111;
      patterns[24062] = 29'b0_101110111111_110_0_101110111111;
      patterns[24063] = 29'b0_101110111111_111_0_101110111111;
      patterns[24064] = 29'b0_101111000000_000_0_101111000000;
      patterns[24065] = 29'b0_101111000000_001_0_000000101111;
      patterns[24066] = 29'b0_101111000000_010_1_011110000000;
      patterns[24067] = 29'b0_101111000000_011_0_111100000001;
      patterns[24068] = 29'b0_101111000000_100_0_010111100000;
      patterns[24069] = 29'b0_101111000000_101_0_001011110000;
      patterns[24070] = 29'b0_101111000000_110_0_101111000000;
      patterns[24071] = 29'b0_101111000000_111_0_101111000000;
      patterns[24072] = 29'b0_101111000001_000_0_101111000001;
      patterns[24073] = 29'b0_101111000001_001_0_000001101111;
      patterns[24074] = 29'b0_101111000001_010_1_011110000010;
      patterns[24075] = 29'b0_101111000001_011_0_111100000101;
      patterns[24076] = 29'b0_101111000001_100_1_010111100000;
      patterns[24077] = 29'b0_101111000001_101_0_101011110000;
      patterns[24078] = 29'b0_101111000001_110_0_101111000001;
      patterns[24079] = 29'b0_101111000001_111_0_101111000001;
      patterns[24080] = 29'b0_101111000010_000_0_101111000010;
      patterns[24081] = 29'b0_101111000010_001_0_000010101111;
      patterns[24082] = 29'b0_101111000010_010_1_011110000100;
      patterns[24083] = 29'b0_101111000010_011_0_111100001001;
      patterns[24084] = 29'b0_101111000010_100_0_010111100001;
      patterns[24085] = 29'b0_101111000010_101_1_001011110000;
      patterns[24086] = 29'b0_101111000010_110_0_101111000010;
      patterns[24087] = 29'b0_101111000010_111_0_101111000010;
      patterns[24088] = 29'b0_101111000011_000_0_101111000011;
      patterns[24089] = 29'b0_101111000011_001_0_000011101111;
      patterns[24090] = 29'b0_101111000011_010_1_011110000110;
      patterns[24091] = 29'b0_101111000011_011_0_111100001101;
      patterns[24092] = 29'b0_101111000011_100_1_010111100001;
      patterns[24093] = 29'b0_101111000011_101_1_101011110000;
      patterns[24094] = 29'b0_101111000011_110_0_101111000011;
      patterns[24095] = 29'b0_101111000011_111_0_101111000011;
      patterns[24096] = 29'b0_101111000100_000_0_101111000100;
      patterns[24097] = 29'b0_101111000100_001_0_000100101111;
      patterns[24098] = 29'b0_101111000100_010_1_011110001000;
      patterns[24099] = 29'b0_101111000100_011_0_111100010001;
      patterns[24100] = 29'b0_101111000100_100_0_010111100010;
      patterns[24101] = 29'b0_101111000100_101_0_001011110001;
      patterns[24102] = 29'b0_101111000100_110_0_101111000100;
      patterns[24103] = 29'b0_101111000100_111_0_101111000100;
      patterns[24104] = 29'b0_101111000101_000_0_101111000101;
      patterns[24105] = 29'b0_101111000101_001_0_000101101111;
      patterns[24106] = 29'b0_101111000101_010_1_011110001010;
      patterns[24107] = 29'b0_101111000101_011_0_111100010101;
      patterns[24108] = 29'b0_101111000101_100_1_010111100010;
      patterns[24109] = 29'b0_101111000101_101_0_101011110001;
      patterns[24110] = 29'b0_101111000101_110_0_101111000101;
      patterns[24111] = 29'b0_101111000101_111_0_101111000101;
      patterns[24112] = 29'b0_101111000110_000_0_101111000110;
      patterns[24113] = 29'b0_101111000110_001_0_000110101111;
      patterns[24114] = 29'b0_101111000110_010_1_011110001100;
      patterns[24115] = 29'b0_101111000110_011_0_111100011001;
      patterns[24116] = 29'b0_101111000110_100_0_010111100011;
      patterns[24117] = 29'b0_101111000110_101_1_001011110001;
      patterns[24118] = 29'b0_101111000110_110_0_101111000110;
      patterns[24119] = 29'b0_101111000110_111_0_101111000110;
      patterns[24120] = 29'b0_101111000111_000_0_101111000111;
      patterns[24121] = 29'b0_101111000111_001_0_000111101111;
      patterns[24122] = 29'b0_101111000111_010_1_011110001110;
      patterns[24123] = 29'b0_101111000111_011_0_111100011101;
      patterns[24124] = 29'b0_101111000111_100_1_010111100011;
      patterns[24125] = 29'b0_101111000111_101_1_101011110001;
      patterns[24126] = 29'b0_101111000111_110_0_101111000111;
      patterns[24127] = 29'b0_101111000111_111_0_101111000111;
      patterns[24128] = 29'b0_101111001000_000_0_101111001000;
      patterns[24129] = 29'b0_101111001000_001_0_001000101111;
      patterns[24130] = 29'b0_101111001000_010_1_011110010000;
      patterns[24131] = 29'b0_101111001000_011_0_111100100001;
      patterns[24132] = 29'b0_101111001000_100_0_010111100100;
      patterns[24133] = 29'b0_101111001000_101_0_001011110010;
      patterns[24134] = 29'b0_101111001000_110_0_101111001000;
      patterns[24135] = 29'b0_101111001000_111_0_101111001000;
      patterns[24136] = 29'b0_101111001001_000_0_101111001001;
      patterns[24137] = 29'b0_101111001001_001_0_001001101111;
      patterns[24138] = 29'b0_101111001001_010_1_011110010010;
      patterns[24139] = 29'b0_101111001001_011_0_111100100101;
      patterns[24140] = 29'b0_101111001001_100_1_010111100100;
      patterns[24141] = 29'b0_101111001001_101_0_101011110010;
      patterns[24142] = 29'b0_101111001001_110_0_101111001001;
      patterns[24143] = 29'b0_101111001001_111_0_101111001001;
      patterns[24144] = 29'b0_101111001010_000_0_101111001010;
      patterns[24145] = 29'b0_101111001010_001_0_001010101111;
      patterns[24146] = 29'b0_101111001010_010_1_011110010100;
      patterns[24147] = 29'b0_101111001010_011_0_111100101001;
      patterns[24148] = 29'b0_101111001010_100_0_010111100101;
      patterns[24149] = 29'b0_101111001010_101_1_001011110010;
      patterns[24150] = 29'b0_101111001010_110_0_101111001010;
      patterns[24151] = 29'b0_101111001010_111_0_101111001010;
      patterns[24152] = 29'b0_101111001011_000_0_101111001011;
      patterns[24153] = 29'b0_101111001011_001_0_001011101111;
      patterns[24154] = 29'b0_101111001011_010_1_011110010110;
      patterns[24155] = 29'b0_101111001011_011_0_111100101101;
      patterns[24156] = 29'b0_101111001011_100_1_010111100101;
      patterns[24157] = 29'b0_101111001011_101_1_101011110010;
      patterns[24158] = 29'b0_101111001011_110_0_101111001011;
      patterns[24159] = 29'b0_101111001011_111_0_101111001011;
      patterns[24160] = 29'b0_101111001100_000_0_101111001100;
      patterns[24161] = 29'b0_101111001100_001_0_001100101111;
      patterns[24162] = 29'b0_101111001100_010_1_011110011000;
      patterns[24163] = 29'b0_101111001100_011_0_111100110001;
      patterns[24164] = 29'b0_101111001100_100_0_010111100110;
      patterns[24165] = 29'b0_101111001100_101_0_001011110011;
      patterns[24166] = 29'b0_101111001100_110_0_101111001100;
      patterns[24167] = 29'b0_101111001100_111_0_101111001100;
      patterns[24168] = 29'b0_101111001101_000_0_101111001101;
      patterns[24169] = 29'b0_101111001101_001_0_001101101111;
      patterns[24170] = 29'b0_101111001101_010_1_011110011010;
      patterns[24171] = 29'b0_101111001101_011_0_111100110101;
      patterns[24172] = 29'b0_101111001101_100_1_010111100110;
      patterns[24173] = 29'b0_101111001101_101_0_101011110011;
      patterns[24174] = 29'b0_101111001101_110_0_101111001101;
      patterns[24175] = 29'b0_101111001101_111_0_101111001101;
      patterns[24176] = 29'b0_101111001110_000_0_101111001110;
      patterns[24177] = 29'b0_101111001110_001_0_001110101111;
      patterns[24178] = 29'b0_101111001110_010_1_011110011100;
      patterns[24179] = 29'b0_101111001110_011_0_111100111001;
      patterns[24180] = 29'b0_101111001110_100_0_010111100111;
      patterns[24181] = 29'b0_101111001110_101_1_001011110011;
      patterns[24182] = 29'b0_101111001110_110_0_101111001110;
      patterns[24183] = 29'b0_101111001110_111_0_101111001110;
      patterns[24184] = 29'b0_101111001111_000_0_101111001111;
      patterns[24185] = 29'b0_101111001111_001_0_001111101111;
      patterns[24186] = 29'b0_101111001111_010_1_011110011110;
      patterns[24187] = 29'b0_101111001111_011_0_111100111101;
      patterns[24188] = 29'b0_101111001111_100_1_010111100111;
      patterns[24189] = 29'b0_101111001111_101_1_101011110011;
      patterns[24190] = 29'b0_101111001111_110_0_101111001111;
      patterns[24191] = 29'b0_101111001111_111_0_101111001111;
      patterns[24192] = 29'b0_101111010000_000_0_101111010000;
      patterns[24193] = 29'b0_101111010000_001_0_010000101111;
      patterns[24194] = 29'b0_101111010000_010_1_011110100000;
      patterns[24195] = 29'b0_101111010000_011_0_111101000001;
      patterns[24196] = 29'b0_101111010000_100_0_010111101000;
      patterns[24197] = 29'b0_101111010000_101_0_001011110100;
      patterns[24198] = 29'b0_101111010000_110_0_101111010000;
      patterns[24199] = 29'b0_101111010000_111_0_101111010000;
      patterns[24200] = 29'b0_101111010001_000_0_101111010001;
      patterns[24201] = 29'b0_101111010001_001_0_010001101111;
      patterns[24202] = 29'b0_101111010001_010_1_011110100010;
      patterns[24203] = 29'b0_101111010001_011_0_111101000101;
      patterns[24204] = 29'b0_101111010001_100_1_010111101000;
      patterns[24205] = 29'b0_101111010001_101_0_101011110100;
      patterns[24206] = 29'b0_101111010001_110_0_101111010001;
      patterns[24207] = 29'b0_101111010001_111_0_101111010001;
      patterns[24208] = 29'b0_101111010010_000_0_101111010010;
      patterns[24209] = 29'b0_101111010010_001_0_010010101111;
      patterns[24210] = 29'b0_101111010010_010_1_011110100100;
      patterns[24211] = 29'b0_101111010010_011_0_111101001001;
      patterns[24212] = 29'b0_101111010010_100_0_010111101001;
      patterns[24213] = 29'b0_101111010010_101_1_001011110100;
      patterns[24214] = 29'b0_101111010010_110_0_101111010010;
      patterns[24215] = 29'b0_101111010010_111_0_101111010010;
      patterns[24216] = 29'b0_101111010011_000_0_101111010011;
      patterns[24217] = 29'b0_101111010011_001_0_010011101111;
      patterns[24218] = 29'b0_101111010011_010_1_011110100110;
      patterns[24219] = 29'b0_101111010011_011_0_111101001101;
      patterns[24220] = 29'b0_101111010011_100_1_010111101001;
      patterns[24221] = 29'b0_101111010011_101_1_101011110100;
      patterns[24222] = 29'b0_101111010011_110_0_101111010011;
      patterns[24223] = 29'b0_101111010011_111_0_101111010011;
      patterns[24224] = 29'b0_101111010100_000_0_101111010100;
      patterns[24225] = 29'b0_101111010100_001_0_010100101111;
      patterns[24226] = 29'b0_101111010100_010_1_011110101000;
      patterns[24227] = 29'b0_101111010100_011_0_111101010001;
      patterns[24228] = 29'b0_101111010100_100_0_010111101010;
      patterns[24229] = 29'b0_101111010100_101_0_001011110101;
      patterns[24230] = 29'b0_101111010100_110_0_101111010100;
      patterns[24231] = 29'b0_101111010100_111_0_101111010100;
      patterns[24232] = 29'b0_101111010101_000_0_101111010101;
      patterns[24233] = 29'b0_101111010101_001_0_010101101111;
      patterns[24234] = 29'b0_101111010101_010_1_011110101010;
      patterns[24235] = 29'b0_101111010101_011_0_111101010101;
      patterns[24236] = 29'b0_101111010101_100_1_010111101010;
      patterns[24237] = 29'b0_101111010101_101_0_101011110101;
      patterns[24238] = 29'b0_101111010101_110_0_101111010101;
      patterns[24239] = 29'b0_101111010101_111_0_101111010101;
      patterns[24240] = 29'b0_101111010110_000_0_101111010110;
      patterns[24241] = 29'b0_101111010110_001_0_010110101111;
      patterns[24242] = 29'b0_101111010110_010_1_011110101100;
      patterns[24243] = 29'b0_101111010110_011_0_111101011001;
      patterns[24244] = 29'b0_101111010110_100_0_010111101011;
      patterns[24245] = 29'b0_101111010110_101_1_001011110101;
      patterns[24246] = 29'b0_101111010110_110_0_101111010110;
      patterns[24247] = 29'b0_101111010110_111_0_101111010110;
      patterns[24248] = 29'b0_101111010111_000_0_101111010111;
      patterns[24249] = 29'b0_101111010111_001_0_010111101111;
      patterns[24250] = 29'b0_101111010111_010_1_011110101110;
      patterns[24251] = 29'b0_101111010111_011_0_111101011101;
      patterns[24252] = 29'b0_101111010111_100_1_010111101011;
      patterns[24253] = 29'b0_101111010111_101_1_101011110101;
      patterns[24254] = 29'b0_101111010111_110_0_101111010111;
      patterns[24255] = 29'b0_101111010111_111_0_101111010111;
      patterns[24256] = 29'b0_101111011000_000_0_101111011000;
      patterns[24257] = 29'b0_101111011000_001_0_011000101111;
      patterns[24258] = 29'b0_101111011000_010_1_011110110000;
      patterns[24259] = 29'b0_101111011000_011_0_111101100001;
      patterns[24260] = 29'b0_101111011000_100_0_010111101100;
      patterns[24261] = 29'b0_101111011000_101_0_001011110110;
      patterns[24262] = 29'b0_101111011000_110_0_101111011000;
      patterns[24263] = 29'b0_101111011000_111_0_101111011000;
      patterns[24264] = 29'b0_101111011001_000_0_101111011001;
      patterns[24265] = 29'b0_101111011001_001_0_011001101111;
      patterns[24266] = 29'b0_101111011001_010_1_011110110010;
      patterns[24267] = 29'b0_101111011001_011_0_111101100101;
      patterns[24268] = 29'b0_101111011001_100_1_010111101100;
      patterns[24269] = 29'b0_101111011001_101_0_101011110110;
      patterns[24270] = 29'b0_101111011001_110_0_101111011001;
      patterns[24271] = 29'b0_101111011001_111_0_101111011001;
      patterns[24272] = 29'b0_101111011010_000_0_101111011010;
      patterns[24273] = 29'b0_101111011010_001_0_011010101111;
      patterns[24274] = 29'b0_101111011010_010_1_011110110100;
      patterns[24275] = 29'b0_101111011010_011_0_111101101001;
      patterns[24276] = 29'b0_101111011010_100_0_010111101101;
      patterns[24277] = 29'b0_101111011010_101_1_001011110110;
      patterns[24278] = 29'b0_101111011010_110_0_101111011010;
      patterns[24279] = 29'b0_101111011010_111_0_101111011010;
      patterns[24280] = 29'b0_101111011011_000_0_101111011011;
      patterns[24281] = 29'b0_101111011011_001_0_011011101111;
      patterns[24282] = 29'b0_101111011011_010_1_011110110110;
      patterns[24283] = 29'b0_101111011011_011_0_111101101101;
      patterns[24284] = 29'b0_101111011011_100_1_010111101101;
      patterns[24285] = 29'b0_101111011011_101_1_101011110110;
      patterns[24286] = 29'b0_101111011011_110_0_101111011011;
      patterns[24287] = 29'b0_101111011011_111_0_101111011011;
      patterns[24288] = 29'b0_101111011100_000_0_101111011100;
      patterns[24289] = 29'b0_101111011100_001_0_011100101111;
      patterns[24290] = 29'b0_101111011100_010_1_011110111000;
      patterns[24291] = 29'b0_101111011100_011_0_111101110001;
      patterns[24292] = 29'b0_101111011100_100_0_010111101110;
      patterns[24293] = 29'b0_101111011100_101_0_001011110111;
      patterns[24294] = 29'b0_101111011100_110_0_101111011100;
      patterns[24295] = 29'b0_101111011100_111_0_101111011100;
      patterns[24296] = 29'b0_101111011101_000_0_101111011101;
      patterns[24297] = 29'b0_101111011101_001_0_011101101111;
      patterns[24298] = 29'b0_101111011101_010_1_011110111010;
      patterns[24299] = 29'b0_101111011101_011_0_111101110101;
      patterns[24300] = 29'b0_101111011101_100_1_010111101110;
      patterns[24301] = 29'b0_101111011101_101_0_101011110111;
      patterns[24302] = 29'b0_101111011101_110_0_101111011101;
      patterns[24303] = 29'b0_101111011101_111_0_101111011101;
      patterns[24304] = 29'b0_101111011110_000_0_101111011110;
      patterns[24305] = 29'b0_101111011110_001_0_011110101111;
      patterns[24306] = 29'b0_101111011110_010_1_011110111100;
      patterns[24307] = 29'b0_101111011110_011_0_111101111001;
      patterns[24308] = 29'b0_101111011110_100_0_010111101111;
      patterns[24309] = 29'b0_101111011110_101_1_001011110111;
      patterns[24310] = 29'b0_101111011110_110_0_101111011110;
      patterns[24311] = 29'b0_101111011110_111_0_101111011110;
      patterns[24312] = 29'b0_101111011111_000_0_101111011111;
      patterns[24313] = 29'b0_101111011111_001_0_011111101111;
      patterns[24314] = 29'b0_101111011111_010_1_011110111110;
      patterns[24315] = 29'b0_101111011111_011_0_111101111101;
      patterns[24316] = 29'b0_101111011111_100_1_010111101111;
      patterns[24317] = 29'b0_101111011111_101_1_101011110111;
      patterns[24318] = 29'b0_101111011111_110_0_101111011111;
      patterns[24319] = 29'b0_101111011111_111_0_101111011111;
      patterns[24320] = 29'b0_101111100000_000_0_101111100000;
      patterns[24321] = 29'b0_101111100000_001_0_100000101111;
      patterns[24322] = 29'b0_101111100000_010_1_011111000000;
      patterns[24323] = 29'b0_101111100000_011_0_111110000001;
      patterns[24324] = 29'b0_101111100000_100_0_010111110000;
      patterns[24325] = 29'b0_101111100000_101_0_001011111000;
      patterns[24326] = 29'b0_101111100000_110_0_101111100000;
      patterns[24327] = 29'b0_101111100000_111_0_101111100000;
      patterns[24328] = 29'b0_101111100001_000_0_101111100001;
      patterns[24329] = 29'b0_101111100001_001_0_100001101111;
      patterns[24330] = 29'b0_101111100001_010_1_011111000010;
      patterns[24331] = 29'b0_101111100001_011_0_111110000101;
      patterns[24332] = 29'b0_101111100001_100_1_010111110000;
      patterns[24333] = 29'b0_101111100001_101_0_101011111000;
      patterns[24334] = 29'b0_101111100001_110_0_101111100001;
      patterns[24335] = 29'b0_101111100001_111_0_101111100001;
      patterns[24336] = 29'b0_101111100010_000_0_101111100010;
      patterns[24337] = 29'b0_101111100010_001_0_100010101111;
      patterns[24338] = 29'b0_101111100010_010_1_011111000100;
      patterns[24339] = 29'b0_101111100010_011_0_111110001001;
      patterns[24340] = 29'b0_101111100010_100_0_010111110001;
      patterns[24341] = 29'b0_101111100010_101_1_001011111000;
      patterns[24342] = 29'b0_101111100010_110_0_101111100010;
      patterns[24343] = 29'b0_101111100010_111_0_101111100010;
      patterns[24344] = 29'b0_101111100011_000_0_101111100011;
      patterns[24345] = 29'b0_101111100011_001_0_100011101111;
      patterns[24346] = 29'b0_101111100011_010_1_011111000110;
      patterns[24347] = 29'b0_101111100011_011_0_111110001101;
      patterns[24348] = 29'b0_101111100011_100_1_010111110001;
      patterns[24349] = 29'b0_101111100011_101_1_101011111000;
      patterns[24350] = 29'b0_101111100011_110_0_101111100011;
      patterns[24351] = 29'b0_101111100011_111_0_101111100011;
      patterns[24352] = 29'b0_101111100100_000_0_101111100100;
      patterns[24353] = 29'b0_101111100100_001_0_100100101111;
      patterns[24354] = 29'b0_101111100100_010_1_011111001000;
      patterns[24355] = 29'b0_101111100100_011_0_111110010001;
      patterns[24356] = 29'b0_101111100100_100_0_010111110010;
      patterns[24357] = 29'b0_101111100100_101_0_001011111001;
      patterns[24358] = 29'b0_101111100100_110_0_101111100100;
      patterns[24359] = 29'b0_101111100100_111_0_101111100100;
      patterns[24360] = 29'b0_101111100101_000_0_101111100101;
      patterns[24361] = 29'b0_101111100101_001_0_100101101111;
      patterns[24362] = 29'b0_101111100101_010_1_011111001010;
      patterns[24363] = 29'b0_101111100101_011_0_111110010101;
      patterns[24364] = 29'b0_101111100101_100_1_010111110010;
      patterns[24365] = 29'b0_101111100101_101_0_101011111001;
      patterns[24366] = 29'b0_101111100101_110_0_101111100101;
      patterns[24367] = 29'b0_101111100101_111_0_101111100101;
      patterns[24368] = 29'b0_101111100110_000_0_101111100110;
      patterns[24369] = 29'b0_101111100110_001_0_100110101111;
      patterns[24370] = 29'b0_101111100110_010_1_011111001100;
      patterns[24371] = 29'b0_101111100110_011_0_111110011001;
      patterns[24372] = 29'b0_101111100110_100_0_010111110011;
      patterns[24373] = 29'b0_101111100110_101_1_001011111001;
      patterns[24374] = 29'b0_101111100110_110_0_101111100110;
      patterns[24375] = 29'b0_101111100110_111_0_101111100110;
      patterns[24376] = 29'b0_101111100111_000_0_101111100111;
      patterns[24377] = 29'b0_101111100111_001_0_100111101111;
      patterns[24378] = 29'b0_101111100111_010_1_011111001110;
      patterns[24379] = 29'b0_101111100111_011_0_111110011101;
      patterns[24380] = 29'b0_101111100111_100_1_010111110011;
      patterns[24381] = 29'b0_101111100111_101_1_101011111001;
      patterns[24382] = 29'b0_101111100111_110_0_101111100111;
      patterns[24383] = 29'b0_101111100111_111_0_101111100111;
      patterns[24384] = 29'b0_101111101000_000_0_101111101000;
      patterns[24385] = 29'b0_101111101000_001_0_101000101111;
      patterns[24386] = 29'b0_101111101000_010_1_011111010000;
      patterns[24387] = 29'b0_101111101000_011_0_111110100001;
      patterns[24388] = 29'b0_101111101000_100_0_010111110100;
      patterns[24389] = 29'b0_101111101000_101_0_001011111010;
      patterns[24390] = 29'b0_101111101000_110_0_101111101000;
      patterns[24391] = 29'b0_101111101000_111_0_101111101000;
      patterns[24392] = 29'b0_101111101001_000_0_101111101001;
      patterns[24393] = 29'b0_101111101001_001_0_101001101111;
      patterns[24394] = 29'b0_101111101001_010_1_011111010010;
      patterns[24395] = 29'b0_101111101001_011_0_111110100101;
      patterns[24396] = 29'b0_101111101001_100_1_010111110100;
      patterns[24397] = 29'b0_101111101001_101_0_101011111010;
      patterns[24398] = 29'b0_101111101001_110_0_101111101001;
      patterns[24399] = 29'b0_101111101001_111_0_101111101001;
      patterns[24400] = 29'b0_101111101010_000_0_101111101010;
      patterns[24401] = 29'b0_101111101010_001_0_101010101111;
      patterns[24402] = 29'b0_101111101010_010_1_011111010100;
      patterns[24403] = 29'b0_101111101010_011_0_111110101001;
      patterns[24404] = 29'b0_101111101010_100_0_010111110101;
      patterns[24405] = 29'b0_101111101010_101_1_001011111010;
      patterns[24406] = 29'b0_101111101010_110_0_101111101010;
      patterns[24407] = 29'b0_101111101010_111_0_101111101010;
      patterns[24408] = 29'b0_101111101011_000_0_101111101011;
      patterns[24409] = 29'b0_101111101011_001_0_101011101111;
      patterns[24410] = 29'b0_101111101011_010_1_011111010110;
      patterns[24411] = 29'b0_101111101011_011_0_111110101101;
      patterns[24412] = 29'b0_101111101011_100_1_010111110101;
      patterns[24413] = 29'b0_101111101011_101_1_101011111010;
      patterns[24414] = 29'b0_101111101011_110_0_101111101011;
      patterns[24415] = 29'b0_101111101011_111_0_101111101011;
      patterns[24416] = 29'b0_101111101100_000_0_101111101100;
      patterns[24417] = 29'b0_101111101100_001_0_101100101111;
      patterns[24418] = 29'b0_101111101100_010_1_011111011000;
      patterns[24419] = 29'b0_101111101100_011_0_111110110001;
      patterns[24420] = 29'b0_101111101100_100_0_010111110110;
      patterns[24421] = 29'b0_101111101100_101_0_001011111011;
      patterns[24422] = 29'b0_101111101100_110_0_101111101100;
      patterns[24423] = 29'b0_101111101100_111_0_101111101100;
      patterns[24424] = 29'b0_101111101101_000_0_101111101101;
      patterns[24425] = 29'b0_101111101101_001_0_101101101111;
      patterns[24426] = 29'b0_101111101101_010_1_011111011010;
      patterns[24427] = 29'b0_101111101101_011_0_111110110101;
      patterns[24428] = 29'b0_101111101101_100_1_010111110110;
      patterns[24429] = 29'b0_101111101101_101_0_101011111011;
      patterns[24430] = 29'b0_101111101101_110_0_101111101101;
      patterns[24431] = 29'b0_101111101101_111_0_101111101101;
      patterns[24432] = 29'b0_101111101110_000_0_101111101110;
      patterns[24433] = 29'b0_101111101110_001_0_101110101111;
      patterns[24434] = 29'b0_101111101110_010_1_011111011100;
      patterns[24435] = 29'b0_101111101110_011_0_111110111001;
      patterns[24436] = 29'b0_101111101110_100_0_010111110111;
      patterns[24437] = 29'b0_101111101110_101_1_001011111011;
      patterns[24438] = 29'b0_101111101110_110_0_101111101110;
      patterns[24439] = 29'b0_101111101110_111_0_101111101110;
      patterns[24440] = 29'b0_101111101111_000_0_101111101111;
      patterns[24441] = 29'b0_101111101111_001_0_101111101111;
      patterns[24442] = 29'b0_101111101111_010_1_011111011110;
      patterns[24443] = 29'b0_101111101111_011_0_111110111101;
      patterns[24444] = 29'b0_101111101111_100_1_010111110111;
      patterns[24445] = 29'b0_101111101111_101_1_101011111011;
      patterns[24446] = 29'b0_101111101111_110_0_101111101111;
      patterns[24447] = 29'b0_101111101111_111_0_101111101111;
      patterns[24448] = 29'b0_101111110000_000_0_101111110000;
      patterns[24449] = 29'b0_101111110000_001_0_110000101111;
      patterns[24450] = 29'b0_101111110000_010_1_011111100000;
      patterns[24451] = 29'b0_101111110000_011_0_111111000001;
      patterns[24452] = 29'b0_101111110000_100_0_010111111000;
      patterns[24453] = 29'b0_101111110000_101_0_001011111100;
      patterns[24454] = 29'b0_101111110000_110_0_101111110000;
      patterns[24455] = 29'b0_101111110000_111_0_101111110000;
      patterns[24456] = 29'b0_101111110001_000_0_101111110001;
      patterns[24457] = 29'b0_101111110001_001_0_110001101111;
      patterns[24458] = 29'b0_101111110001_010_1_011111100010;
      patterns[24459] = 29'b0_101111110001_011_0_111111000101;
      patterns[24460] = 29'b0_101111110001_100_1_010111111000;
      patterns[24461] = 29'b0_101111110001_101_0_101011111100;
      patterns[24462] = 29'b0_101111110001_110_0_101111110001;
      patterns[24463] = 29'b0_101111110001_111_0_101111110001;
      patterns[24464] = 29'b0_101111110010_000_0_101111110010;
      patterns[24465] = 29'b0_101111110010_001_0_110010101111;
      patterns[24466] = 29'b0_101111110010_010_1_011111100100;
      patterns[24467] = 29'b0_101111110010_011_0_111111001001;
      patterns[24468] = 29'b0_101111110010_100_0_010111111001;
      patterns[24469] = 29'b0_101111110010_101_1_001011111100;
      patterns[24470] = 29'b0_101111110010_110_0_101111110010;
      patterns[24471] = 29'b0_101111110010_111_0_101111110010;
      patterns[24472] = 29'b0_101111110011_000_0_101111110011;
      patterns[24473] = 29'b0_101111110011_001_0_110011101111;
      patterns[24474] = 29'b0_101111110011_010_1_011111100110;
      patterns[24475] = 29'b0_101111110011_011_0_111111001101;
      patterns[24476] = 29'b0_101111110011_100_1_010111111001;
      patterns[24477] = 29'b0_101111110011_101_1_101011111100;
      patterns[24478] = 29'b0_101111110011_110_0_101111110011;
      patterns[24479] = 29'b0_101111110011_111_0_101111110011;
      patterns[24480] = 29'b0_101111110100_000_0_101111110100;
      patterns[24481] = 29'b0_101111110100_001_0_110100101111;
      patterns[24482] = 29'b0_101111110100_010_1_011111101000;
      patterns[24483] = 29'b0_101111110100_011_0_111111010001;
      patterns[24484] = 29'b0_101111110100_100_0_010111111010;
      patterns[24485] = 29'b0_101111110100_101_0_001011111101;
      patterns[24486] = 29'b0_101111110100_110_0_101111110100;
      patterns[24487] = 29'b0_101111110100_111_0_101111110100;
      patterns[24488] = 29'b0_101111110101_000_0_101111110101;
      patterns[24489] = 29'b0_101111110101_001_0_110101101111;
      patterns[24490] = 29'b0_101111110101_010_1_011111101010;
      patterns[24491] = 29'b0_101111110101_011_0_111111010101;
      patterns[24492] = 29'b0_101111110101_100_1_010111111010;
      patterns[24493] = 29'b0_101111110101_101_0_101011111101;
      patterns[24494] = 29'b0_101111110101_110_0_101111110101;
      patterns[24495] = 29'b0_101111110101_111_0_101111110101;
      patterns[24496] = 29'b0_101111110110_000_0_101111110110;
      patterns[24497] = 29'b0_101111110110_001_0_110110101111;
      patterns[24498] = 29'b0_101111110110_010_1_011111101100;
      patterns[24499] = 29'b0_101111110110_011_0_111111011001;
      patterns[24500] = 29'b0_101111110110_100_0_010111111011;
      patterns[24501] = 29'b0_101111110110_101_1_001011111101;
      patterns[24502] = 29'b0_101111110110_110_0_101111110110;
      patterns[24503] = 29'b0_101111110110_111_0_101111110110;
      patterns[24504] = 29'b0_101111110111_000_0_101111110111;
      patterns[24505] = 29'b0_101111110111_001_0_110111101111;
      patterns[24506] = 29'b0_101111110111_010_1_011111101110;
      patterns[24507] = 29'b0_101111110111_011_0_111111011101;
      patterns[24508] = 29'b0_101111110111_100_1_010111111011;
      patterns[24509] = 29'b0_101111110111_101_1_101011111101;
      patterns[24510] = 29'b0_101111110111_110_0_101111110111;
      patterns[24511] = 29'b0_101111110111_111_0_101111110111;
      patterns[24512] = 29'b0_101111111000_000_0_101111111000;
      patterns[24513] = 29'b0_101111111000_001_0_111000101111;
      patterns[24514] = 29'b0_101111111000_010_1_011111110000;
      patterns[24515] = 29'b0_101111111000_011_0_111111100001;
      patterns[24516] = 29'b0_101111111000_100_0_010111111100;
      patterns[24517] = 29'b0_101111111000_101_0_001011111110;
      patterns[24518] = 29'b0_101111111000_110_0_101111111000;
      patterns[24519] = 29'b0_101111111000_111_0_101111111000;
      patterns[24520] = 29'b0_101111111001_000_0_101111111001;
      patterns[24521] = 29'b0_101111111001_001_0_111001101111;
      patterns[24522] = 29'b0_101111111001_010_1_011111110010;
      patterns[24523] = 29'b0_101111111001_011_0_111111100101;
      patterns[24524] = 29'b0_101111111001_100_1_010111111100;
      patterns[24525] = 29'b0_101111111001_101_0_101011111110;
      patterns[24526] = 29'b0_101111111001_110_0_101111111001;
      patterns[24527] = 29'b0_101111111001_111_0_101111111001;
      patterns[24528] = 29'b0_101111111010_000_0_101111111010;
      patterns[24529] = 29'b0_101111111010_001_0_111010101111;
      patterns[24530] = 29'b0_101111111010_010_1_011111110100;
      patterns[24531] = 29'b0_101111111010_011_0_111111101001;
      patterns[24532] = 29'b0_101111111010_100_0_010111111101;
      patterns[24533] = 29'b0_101111111010_101_1_001011111110;
      patterns[24534] = 29'b0_101111111010_110_0_101111111010;
      patterns[24535] = 29'b0_101111111010_111_0_101111111010;
      patterns[24536] = 29'b0_101111111011_000_0_101111111011;
      patterns[24537] = 29'b0_101111111011_001_0_111011101111;
      patterns[24538] = 29'b0_101111111011_010_1_011111110110;
      patterns[24539] = 29'b0_101111111011_011_0_111111101101;
      patterns[24540] = 29'b0_101111111011_100_1_010111111101;
      patterns[24541] = 29'b0_101111111011_101_1_101011111110;
      patterns[24542] = 29'b0_101111111011_110_0_101111111011;
      patterns[24543] = 29'b0_101111111011_111_0_101111111011;
      patterns[24544] = 29'b0_101111111100_000_0_101111111100;
      patterns[24545] = 29'b0_101111111100_001_0_111100101111;
      patterns[24546] = 29'b0_101111111100_010_1_011111111000;
      patterns[24547] = 29'b0_101111111100_011_0_111111110001;
      patterns[24548] = 29'b0_101111111100_100_0_010111111110;
      patterns[24549] = 29'b0_101111111100_101_0_001011111111;
      patterns[24550] = 29'b0_101111111100_110_0_101111111100;
      patterns[24551] = 29'b0_101111111100_111_0_101111111100;
      patterns[24552] = 29'b0_101111111101_000_0_101111111101;
      patterns[24553] = 29'b0_101111111101_001_0_111101101111;
      patterns[24554] = 29'b0_101111111101_010_1_011111111010;
      patterns[24555] = 29'b0_101111111101_011_0_111111110101;
      patterns[24556] = 29'b0_101111111101_100_1_010111111110;
      patterns[24557] = 29'b0_101111111101_101_0_101011111111;
      patterns[24558] = 29'b0_101111111101_110_0_101111111101;
      patterns[24559] = 29'b0_101111111101_111_0_101111111101;
      patterns[24560] = 29'b0_101111111110_000_0_101111111110;
      patterns[24561] = 29'b0_101111111110_001_0_111110101111;
      patterns[24562] = 29'b0_101111111110_010_1_011111111100;
      patterns[24563] = 29'b0_101111111110_011_0_111111111001;
      patterns[24564] = 29'b0_101111111110_100_0_010111111111;
      patterns[24565] = 29'b0_101111111110_101_1_001011111111;
      patterns[24566] = 29'b0_101111111110_110_0_101111111110;
      patterns[24567] = 29'b0_101111111110_111_0_101111111110;
      patterns[24568] = 29'b0_101111111111_000_0_101111111111;
      patterns[24569] = 29'b0_101111111111_001_0_111111101111;
      patterns[24570] = 29'b0_101111111111_010_1_011111111110;
      patterns[24571] = 29'b0_101111111111_011_0_111111111101;
      patterns[24572] = 29'b0_101111111111_100_1_010111111111;
      patterns[24573] = 29'b0_101111111111_101_1_101011111111;
      patterns[24574] = 29'b0_101111111111_110_0_101111111111;
      patterns[24575] = 29'b0_101111111111_111_0_101111111111;
      patterns[24576] = 29'b0_110000000000_000_0_110000000000;
      patterns[24577] = 29'b0_110000000000_001_0_000000110000;
      patterns[24578] = 29'b0_110000000000_010_1_100000000000;
      patterns[24579] = 29'b0_110000000000_011_1_000000000001;
      patterns[24580] = 29'b0_110000000000_100_0_011000000000;
      patterns[24581] = 29'b0_110000000000_101_0_001100000000;
      patterns[24582] = 29'b0_110000000000_110_0_110000000000;
      patterns[24583] = 29'b0_110000000000_111_0_110000000000;
      patterns[24584] = 29'b0_110000000001_000_0_110000000001;
      patterns[24585] = 29'b0_110000000001_001_0_000001110000;
      patterns[24586] = 29'b0_110000000001_010_1_100000000010;
      patterns[24587] = 29'b0_110000000001_011_1_000000000101;
      patterns[24588] = 29'b0_110000000001_100_1_011000000000;
      patterns[24589] = 29'b0_110000000001_101_0_101100000000;
      patterns[24590] = 29'b0_110000000001_110_0_110000000001;
      patterns[24591] = 29'b0_110000000001_111_0_110000000001;
      patterns[24592] = 29'b0_110000000010_000_0_110000000010;
      patterns[24593] = 29'b0_110000000010_001_0_000010110000;
      patterns[24594] = 29'b0_110000000010_010_1_100000000100;
      patterns[24595] = 29'b0_110000000010_011_1_000000001001;
      patterns[24596] = 29'b0_110000000010_100_0_011000000001;
      patterns[24597] = 29'b0_110000000010_101_1_001100000000;
      patterns[24598] = 29'b0_110000000010_110_0_110000000010;
      patterns[24599] = 29'b0_110000000010_111_0_110000000010;
      patterns[24600] = 29'b0_110000000011_000_0_110000000011;
      patterns[24601] = 29'b0_110000000011_001_0_000011110000;
      patterns[24602] = 29'b0_110000000011_010_1_100000000110;
      patterns[24603] = 29'b0_110000000011_011_1_000000001101;
      patterns[24604] = 29'b0_110000000011_100_1_011000000001;
      patterns[24605] = 29'b0_110000000011_101_1_101100000000;
      patterns[24606] = 29'b0_110000000011_110_0_110000000011;
      patterns[24607] = 29'b0_110000000011_111_0_110000000011;
      patterns[24608] = 29'b0_110000000100_000_0_110000000100;
      patterns[24609] = 29'b0_110000000100_001_0_000100110000;
      patterns[24610] = 29'b0_110000000100_010_1_100000001000;
      patterns[24611] = 29'b0_110000000100_011_1_000000010001;
      patterns[24612] = 29'b0_110000000100_100_0_011000000010;
      patterns[24613] = 29'b0_110000000100_101_0_001100000001;
      patterns[24614] = 29'b0_110000000100_110_0_110000000100;
      patterns[24615] = 29'b0_110000000100_111_0_110000000100;
      patterns[24616] = 29'b0_110000000101_000_0_110000000101;
      patterns[24617] = 29'b0_110000000101_001_0_000101110000;
      patterns[24618] = 29'b0_110000000101_010_1_100000001010;
      patterns[24619] = 29'b0_110000000101_011_1_000000010101;
      patterns[24620] = 29'b0_110000000101_100_1_011000000010;
      patterns[24621] = 29'b0_110000000101_101_0_101100000001;
      patterns[24622] = 29'b0_110000000101_110_0_110000000101;
      patterns[24623] = 29'b0_110000000101_111_0_110000000101;
      patterns[24624] = 29'b0_110000000110_000_0_110000000110;
      patterns[24625] = 29'b0_110000000110_001_0_000110110000;
      patterns[24626] = 29'b0_110000000110_010_1_100000001100;
      patterns[24627] = 29'b0_110000000110_011_1_000000011001;
      patterns[24628] = 29'b0_110000000110_100_0_011000000011;
      patterns[24629] = 29'b0_110000000110_101_1_001100000001;
      patterns[24630] = 29'b0_110000000110_110_0_110000000110;
      patterns[24631] = 29'b0_110000000110_111_0_110000000110;
      patterns[24632] = 29'b0_110000000111_000_0_110000000111;
      patterns[24633] = 29'b0_110000000111_001_0_000111110000;
      patterns[24634] = 29'b0_110000000111_010_1_100000001110;
      patterns[24635] = 29'b0_110000000111_011_1_000000011101;
      patterns[24636] = 29'b0_110000000111_100_1_011000000011;
      patterns[24637] = 29'b0_110000000111_101_1_101100000001;
      patterns[24638] = 29'b0_110000000111_110_0_110000000111;
      patterns[24639] = 29'b0_110000000111_111_0_110000000111;
      patterns[24640] = 29'b0_110000001000_000_0_110000001000;
      patterns[24641] = 29'b0_110000001000_001_0_001000110000;
      patterns[24642] = 29'b0_110000001000_010_1_100000010000;
      patterns[24643] = 29'b0_110000001000_011_1_000000100001;
      patterns[24644] = 29'b0_110000001000_100_0_011000000100;
      patterns[24645] = 29'b0_110000001000_101_0_001100000010;
      patterns[24646] = 29'b0_110000001000_110_0_110000001000;
      patterns[24647] = 29'b0_110000001000_111_0_110000001000;
      patterns[24648] = 29'b0_110000001001_000_0_110000001001;
      patterns[24649] = 29'b0_110000001001_001_0_001001110000;
      patterns[24650] = 29'b0_110000001001_010_1_100000010010;
      patterns[24651] = 29'b0_110000001001_011_1_000000100101;
      patterns[24652] = 29'b0_110000001001_100_1_011000000100;
      patterns[24653] = 29'b0_110000001001_101_0_101100000010;
      patterns[24654] = 29'b0_110000001001_110_0_110000001001;
      patterns[24655] = 29'b0_110000001001_111_0_110000001001;
      patterns[24656] = 29'b0_110000001010_000_0_110000001010;
      patterns[24657] = 29'b0_110000001010_001_0_001010110000;
      patterns[24658] = 29'b0_110000001010_010_1_100000010100;
      patterns[24659] = 29'b0_110000001010_011_1_000000101001;
      patterns[24660] = 29'b0_110000001010_100_0_011000000101;
      patterns[24661] = 29'b0_110000001010_101_1_001100000010;
      patterns[24662] = 29'b0_110000001010_110_0_110000001010;
      patterns[24663] = 29'b0_110000001010_111_0_110000001010;
      patterns[24664] = 29'b0_110000001011_000_0_110000001011;
      patterns[24665] = 29'b0_110000001011_001_0_001011110000;
      patterns[24666] = 29'b0_110000001011_010_1_100000010110;
      patterns[24667] = 29'b0_110000001011_011_1_000000101101;
      patterns[24668] = 29'b0_110000001011_100_1_011000000101;
      patterns[24669] = 29'b0_110000001011_101_1_101100000010;
      patterns[24670] = 29'b0_110000001011_110_0_110000001011;
      patterns[24671] = 29'b0_110000001011_111_0_110000001011;
      patterns[24672] = 29'b0_110000001100_000_0_110000001100;
      patterns[24673] = 29'b0_110000001100_001_0_001100110000;
      patterns[24674] = 29'b0_110000001100_010_1_100000011000;
      patterns[24675] = 29'b0_110000001100_011_1_000000110001;
      patterns[24676] = 29'b0_110000001100_100_0_011000000110;
      patterns[24677] = 29'b0_110000001100_101_0_001100000011;
      patterns[24678] = 29'b0_110000001100_110_0_110000001100;
      patterns[24679] = 29'b0_110000001100_111_0_110000001100;
      patterns[24680] = 29'b0_110000001101_000_0_110000001101;
      patterns[24681] = 29'b0_110000001101_001_0_001101110000;
      patterns[24682] = 29'b0_110000001101_010_1_100000011010;
      patterns[24683] = 29'b0_110000001101_011_1_000000110101;
      patterns[24684] = 29'b0_110000001101_100_1_011000000110;
      patterns[24685] = 29'b0_110000001101_101_0_101100000011;
      patterns[24686] = 29'b0_110000001101_110_0_110000001101;
      patterns[24687] = 29'b0_110000001101_111_0_110000001101;
      patterns[24688] = 29'b0_110000001110_000_0_110000001110;
      patterns[24689] = 29'b0_110000001110_001_0_001110110000;
      patterns[24690] = 29'b0_110000001110_010_1_100000011100;
      patterns[24691] = 29'b0_110000001110_011_1_000000111001;
      patterns[24692] = 29'b0_110000001110_100_0_011000000111;
      patterns[24693] = 29'b0_110000001110_101_1_001100000011;
      patterns[24694] = 29'b0_110000001110_110_0_110000001110;
      patterns[24695] = 29'b0_110000001110_111_0_110000001110;
      patterns[24696] = 29'b0_110000001111_000_0_110000001111;
      patterns[24697] = 29'b0_110000001111_001_0_001111110000;
      patterns[24698] = 29'b0_110000001111_010_1_100000011110;
      patterns[24699] = 29'b0_110000001111_011_1_000000111101;
      patterns[24700] = 29'b0_110000001111_100_1_011000000111;
      patterns[24701] = 29'b0_110000001111_101_1_101100000011;
      patterns[24702] = 29'b0_110000001111_110_0_110000001111;
      patterns[24703] = 29'b0_110000001111_111_0_110000001111;
      patterns[24704] = 29'b0_110000010000_000_0_110000010000;
      patterns[24705] = 29'b0_110000010000_001_0_010000110000;
      patterns[24706] = 29'b0_110000010000_010_1_100000100000;
      patterns[24707] = 29'b0_110000010000_011_1_000001000001;
      patterns[24708] = 29'b0_110000010000_100_0_011000001000;
      patterns[24709] = 29'b0_110000010000_101_0_001100000100;
      patterns[24710] = 29'b0_110000010000_110_0_110000010000;
      patterns[24711] = 29'b0_110000010000_111_0_110000010000;
      patterns[24712] = 29'b0_110000010001_000_0_110000010001;
      patterns[24713] = 29'b0_110000010001_001_0_010001110000;
      patterns[24714] = 29'b0_110000010001_010_1_100000100010;
      patterns[24715] = 29'b0_110000010001_011_1_000001000101;
      patterns[24716] = 29'b0_110000010001_100_1_011000001000;
      patterns[24717] = 29'b0_110000010001_101_0_101100000100;
      patterns[24718] = 29'b0_110000010001_110_0_110000010001;
      patterns[24719] = 29'b0_110000010001_111_0_110000010001;
      patterns[24720] = 29'b0_110000010010_000_0_110000010010;
      patterns[24721] = 29'b0_110000010010_001_0_010010110000;
      patterns[24722] = 29'b0_110000010010_010_1_100000100100;
      patterns[24723] = 29'b0_110000010010_011_1_000001001001;
      patterns[24724] = 29'b0_110000010010_100_0_011000001001;
      patterns[24725] = 29'b0_110000010010_101_1_001100000100;
      patterns[24726] = 29'b0_110000010010_110_0_110000010010;
      patterns[24727] = 29'b0_110000010010_111_0_110000010010;
      patterns[24728] = 29'b0_110000010011_000_0_110000010011;
      patterns[24729] = 29'b0_110000010011_001_0_010011110000;
      patterns[24730] = 29'b0_110000010011_010_1_100000100110;
      patterns[24731] = 29'b0_110000010011_011_1_000001001101;
      patterns[24732] = 29'b0_110000010011_100_1_011000001001;
      patterns[24733] = 29'b0_110000010011_101_1_101100000100;
      patterns[24734] = 29'b0_110000010011_110_0_110000010011;
      patterns[24735] = 29'b0_110000010011_111_0_110000010011;
      patterns[24736] = 29'b0_110000010100_000_0_110000010100;
      patterns[24737] = 29'b0_110000010100_001_0_010100110000;
      patterns[24738] = 29'b0_110000010100_010_1_100000101000;
      patterns[24739] = 29'b0_110000010100_011_1_000001010001;
      patterns[24740] = 29'b0_110000010100_100_0_011000001010;
      patterns[24741] = 29'b0_110000010100_101_0_001100000101;
      patterns[24742] = 29'b0_110000010100_110_0_110000010100;
      patterns[24743] = 29'b0_110000010100_111_0_110000010100;
      patterns[24744] = 29'b0_110000010101_000_0_110000010101;
      patterns[24745] = 29'b0_110000010101_001_0_010101110000;
      patterns[24746] = 29'b0_110000010101_010_1_100000101010;
      patterns[24747] = 29'b0_110000010101_011_1_000001010101;
      patterns[24748] = 29'b0_110000010101_100_1_011000001010;
      patterns[24749] = 29'b0_110000010101_101_0_101100000101;
      patterns[24750] = 29'b0_110000010101_110_0_110000010101;
      patterns[24751] = 29'b0_110000010101_111_0_110000010101;
      patterns[24752] = 29'b0_110000010110_000_0_110000010110;
      patterns[24753] = 29'b0_110000010110_001_0_010110110000;
      patterns[24754] = 29'b0_110000010110_010_1_100000101100;
      patterns[24755] = 29'b0_110000010110_011_1_000001011001;
      patterns[24756] = 29'b0_110000010110_100_0_011000001011;
      patterns[24757] = 29'b0_110000010110_101_1_001100000101;
      patterns[24758] = 29'b0_110000010110_110_0_110000010110;
      patterns[24759] = 29'b0_110000010110_111_0_110000010110;
      patterns[24760] = 29'b0_110000010111_000_0_110000010111;
      patterns[24761] = 29'b0_110000010111_001_0_010111110000;
      patterns[24762] = 29'b0_110000010111_010_1_100000101110;
      patterns[24763] = 29'b0_110000010111_011_1_000001011101;
      patterns[24764] = 29'b0_110000010111_100_1_011000001011;
      patterns[24765] = 29'b0_110000010111_101_1_101100000101;
      patterns[24766] = 29'b0_110000010111_110_0_110000010111;
      patterns[24767] = 29'b0_110000010111_111_0_110000010111;
      patterns[24768] = 29'b0_110000011000_000_0_110000011000;
      patterns[24769] = 29'b0_110000011000_001_0_011000110000;
      patterns[24770] = 29'b0_110000011000_010_1_100000110000;
      patterns[24771] = 29'b0_110000011000_011_1_000001100001;
      patterns[24772] = 29'b0_110000011000_100_0_011000001100;
      patterns[24773] = 29'b0_110000011000_101_0_001100000110;
      patterns[24774] = 29'b0_110000011000_110_0_110000011000;
      patterns[24775] = 29'b0_110000011000_111_0_110000011000;
      patterns[24776] = 29'b0_110000011001_000_0_110000011001;
      patterns[24777] = 29'b0_110000011001_001_0_011001110000;
      patterns[24778] = 29'b0_110000011001_010_1_100000110010;
      patterns[24779] = 29'b0_110000011001_011_1_000001100101;
      patterns[24780] = 29'b0_110000011001_100_1_011000001100;
      patterns[24781] = 29'b0_110000011001_101_0_101100000110;
      patterns[24782] = 29'b0_110000011001_110_0_110000011001;
      patterns[24783] = 29'b0_110000011001_111_0_110000011001;
      patterns[24784] = 29'b0_110000011010_000_0_110000011010;
      patterns[24785] = 29'b0_110000011010_001_0_011010110000;
      patterns[24786] = 29'b0_110000011010_010_1_100000110100;
      patterns[24787] = 29'b0_110000011010_011_1_000001101001;
      patterns[24788] = 29'b0_110000011010_100_0_011000001101;
      patterns[24789] = 29'b0_110000011010_101_1_001100000110;
      patterns[24790] = 29'b0_110000011010_110_0_110000011010;
      patterns[24791] = 29'b0_110000011010_111_0_110000011010;
      patterns[24792] = 29'b0_110000011011_000_0_110000011011;
      patterns[24793] = 29'b0_110000011011_001_0_011011110000;
      patterns[24794] = 29'b0_110000011011_010_1_100000110110;
      patterns[24795] = 29'b0_110000011011_011_1_000001101101;
      patterns[24796] = 29'b0_110000011011_100_1_011000001101;
      patterns[24797] = 29'b0_110000011011_101_1_101100000110;
      patterns[24798] = 29'b0_110000011011_110_0_110000011011;
      patterns[24799] = 29'b0_110000011011_111_0_110000011011;
      patterns[24800] = 29'b0_110000011100_000_0_110000011100;
      patterns[24801] = 29'b0_110000011100_001_0_011100110000;
      patterns[24802] = 29'b0_110000011100_010_1_100000111000;
      patterns[24803] = 29'b0_110000011100_011_1_000001110001;
      patterns[24804] = 29'b0_110000011100_100_0_011000001110;
      patterns[24805] = 29'b0_110000011100_101_0_001100000111;
      patterns[24806] = 29'b0_110000011100_110_0_110000011100;
      patterns[24807] = 29'b0_110000011100_111_0_110000011100;
      patterns[24808] = 29'b0_110000011101_000_0_110000011101;
      patterns[24809] = 29'b0_110000011101_001_0_011101110000;
      patterns[24810] = 29'b0_110000011101_010_1_100000111010;
      patterns[24811] = 29'b0_110000011101_011_1_000001110101;
      patterns[24812] = 29'b0_110000011101_100_1_011000001110;
      patterns[24813] = 29'b0_110000011101_101_0_101100000111;
      patterns[24814] = 29'b0_110000011101_110_0_110000011101;
      patterns[24815] = 29'b0_110000011101_111_0_110000011101;
      patterns[24816] = 29'b0_110000011110_000_0_110000011110;
      patterns[24817] = 29'b0_110000011110_001_0_011110110000;
      patterns[24818] = 29'b0_110000011110_010_1_100000111100;
      patterns[24819] = 29'b0_110000011110_011_1_000001111001;
      patterns[24820] = 29'b0_110000011110_100_0_011000001111;
      patterns[24821] = 29'b0_110000011110_101_1_001100000111;
      patterns[24822] = 29'b0_110000011110_110_0_110000011110;
      patterns[24823] = 29'b0_110000011110_111_0_110000011110;
      patterns[24824] = 29'b0_110000011111_000_0_110000011111;
      patterns[24825] = 29'b0_110000011111_001_0_011111110000;
      patterns[24826] = 29'b0_110000011111_010_1_100000111110;
      patterns[24827] = 29'b0_110000011111_011_1_000001111101;
      patterns[24828] = 29'b0_110000011111_100_1_011000001111;
      patterns[24829] = 29'b0_110000011111_101_1_101100000111;
      patterns[24830] = 29'b0_110000011111_110_0_110000011111;
      patterns[24831] = 29'b0_110000011111_111_0_110000011111;
      patterns[24832] = 29'b0_110000100000_000_0_110000100000;
      patterns[24833] = 29'b0_110000100000_001_0_100000110000;
      patterns[24834] = 29'b0_110000100000_010_1_100001000000;
      patterns[24835] = 29'b0_110000100000_011_1_000010000001;
      patterns[24836] = 29'b0_110000100000_100_0_011000010000;
      patterns[24837] = 29'b0_110000100000_101_0_001100001000;
      patterns[24838] = 29'b0_110000100000_110_0_110000100000;
      patterns[24839] = 29'b0_110000100000_111_0_110000100000;
      patterns[24840] = 29'b0_110000100001_000_0_110000100001;
      patterns[24841] = 29'b0_110000100001_001_0_100001110000;
      patterns[24842] = 29'b0_110000100001_010_1_100001000010;
      patterns[24843] = 29'b0_110000100001_011_1_000010000101;
      patterns[24844] = 29'b0_110000100001_100_1_011000010000;
      patterns[24845] = 29'b0_110000100001_101_0_101100001000;
      patterns[24846] = 29'b0_110000100001_110_0_110000100001;
      patterns[24847] = 29'b0_110000100001_111_0_110000100001;
      patterns[24848] = 29'b0_110000100010_000_0_110000100010;
      patterns[24849] = 29'b0_110000100010_001_0_100010110000;
      patterns[24850] = 29'b0_110000100010_010_1_100001000100;
      patterns[24851] = 29'b0_110000100010_011_1_000010001001;
      patterns[24852] = 29'b0_110000100010_100_0_011000010001;
      patterns[24853] = 29'b0_110000100010_101_1_001100001000;
      patterns[24854] = 29'b0_110000100010_110_0_110000100010;
      patterns[24855] = 29'b0_110000100010_111_0_110000100010;
      patterns[24856] = 29'b0_110000100011_000_0_110000100011;
      patterns[24857] = 29'b0_110000100011_001_0_100011110000;
      patterns[24858] = 29'b0_110000100011_010_1_100001000110;
      patterns[24859] = 29'b0_110000100011_011_1_000010001101;
      patterns[24860] = 29'b0_110000100011_100_1_011000010001;
      patterns[24861] = 29'b0_110000100011_101_1_101100001000;
      patterns[24862] = 29'b0_110000100011_110_0_110000100011;
      patterns[24863] = 29'b0_110000100011_111_0_110000100011;
      patterns[24864] = 29'b0_110000100100_000_0_110000100100;
      patterns[24865] = 29'b0_110000100100_001_0_100100110000;
      patterns[24866] = 29'b0_110000100100_010_1_100001001000;
      patterns[24867] = 29'b0_110000100100_011_1_000010010001;
      patterns[24868] = 29'b0_110000100100_100_0_011000010010;
      patterns[24869] = 29'b0_110000100100_101_0_001100001001;
      patterns[24870] = 29'b0_110000100100_110_0_110000100100;
      patterns[24871] = 29'b0_110000100100_111_0_110000100100;
      patterns[24872] = 29'b0_110000100101_000_0_110000100101;
      patterns[24873] = 29'b0_110000100101_001_0_100101110000;
      patterns[24874] = 29'b0_110000100101_010_1_100001001010;
      patterns[24875] = 29'b0_110000100101_011_1_000010010101;
      patterns[24876] = 29'b0_110000100101_100_1_011000010010;
      patterns[24877] = 29'b0_110000100101_101_0_101100001001;
      patterns[24878] = 29'b0_110000100101_110_0_110000100101;
      patterns[24879] = 29'b0_110000100101_111_0_110000100101;
      patterns[24880] = 29'b0_110000100110_000_0_110000100110;
      patterns[24881] = 29'b0_110000100110_001_0_100110110000;
      patterns[24882] = 29'b0_110000100110_010_1_100001001100;
      patterns[24883] = 29'b0_110000100110_011_1_000010011001;
      patterns[24884] = 29'b0_110000100110_100_0_011000010011;
      patterns[24885] = 29'b0_110000100110_101_1_001100001001;
      patterns[24886] = 29'b0_110000100110_110_0_110000100110;
      patterns[24887] = 29'b0_110000100110_111_0_110000100110;
      patterns[24888] = 29'b0_110000100111_000_0_110000100111;
      patterns[24889] = 29'b0_110000100111_001_0_100111110000;
      patterns[24890] = 29'b0_110000100111_010_1_100001001110;
      patterns[24891] = 29'b0_110000100111_011_1_000010011101;
      patterns[24892] = 29'b0_110000100111_100_1_011000010011;
      patterns[24893] = 29'b0_110000100111_101_1_101100001001;
      patterns[24894] = 29'b0_110000100111_110_0_110000100111;
      patterns[24895] = 29'b0_110000100111_111_0_110000100111;
      patterns[24896] = 29'b0_110000101000_000_0_110000101000;
      patterns[24897] = 29'b0_110000101000_001_0_101000110000;
      patterns[24898] = 29'b0_110000101000_010_1_100001010000;
      patterns[24899] = 29'b0_110000101000_011_1_000010100001;
      patterns[24900] = 29'b0_110000101000_100_0_011000010100;
      patterns[24901] = 29'b0_110000101000_101_0_001100001010;
      patterns[24902] = 29'b0_110000101000_110_0_110000101000;
      patterns[24903] = 29'b0_110000101000_111_0_110000101000;
      patterns[24904] = 29'b0_110000101001_000_0_110000101001;
      patterns[24905] = 29'b0_110000101001_001_0_101001110000;
      patterns[24906] = 29'b0_110000101001_010_1_100001010010;
      patterns[24907] = 29'b0_110000101001_011_1_000010100101;
      patterns[24908] = 29'b0_110000101001_100_1_011000010100;
      patterns[24909] = 29'b0_110000101001_101_0_101100001010;
      patterns[24910] = 29'b0_110000101001_110_0_110000101001;
      patterns[24911] = 29'b0_110000101001_111_0_110000101001;
      patterns[24912] = 29'b0_110000101010_000_0_110000101010;
      patterns[24913] = 29'b0_110000101010_001_0_101010110000;
      patterns[24914] = 29'b0_110000101010_010_1_100001010100;
      patterns[24915] = 29'b0_110000101010_011_1_000010101001;
      patterns[24916] = 29'b0_110000101010_100_0_011000010101;
      patterns[24917] = 29'b0_110000101010_101_1_001100001010;
      patterns[24918] = 29'b0_110000101010_110_0_110000101010;
      patterns[24919] = 29'b0_110000101010_111_0_110000101010;
      patterns[24920] = 29'b0_110000101011_000_0_110000101011;
      patterns[24921] = 29'b0_110000101011_001_0_101011110000;
      patterns[24922] = 29'b0_110000101011_010_1_100001010110;
      patterns[24923] = 29'b0_110000101011_011_1_000010101101;
      patterns[24924] = 29'b0_110000101011_100_1_011000010101;
      patterns[24925] = 29'b0_110000101011_101_1_101100001010;
      patterns[24926] = 29'b0_110000101011_110_0_110000101011;
      patterns[24927] = 29'b0_110000101011_111_0_110000101011;
      patterns[24928] = 29'b0_110000101100_000_0_110000101100;
      patterns[24929] = 29'b0_110000101100_001_0_101100110000;
      patterns[24930] = 29'b0_110000101100_010_1_100001011000;
      patterns[24931] = 29'b0_110000101100_011_1_000010110001;
      patterns[24932] = 29'b0_110000101100_100_0_011000010110;
      patterns[24933] = 29'b0_110000101100_101_0_001100001011;
      patterns[24934] = 29'b0_110000101100_110_0_110000101100;
      patterns[24935] = 29'b0_110000101100_111_0_110000101100;
      patterns[24936] = 29'b0_110000101101_000_0_110000101101;
      patterns[24937] = 29'b0_110000101101_001_0_101101110000;
      patterns[24938] = 29'b0_110000101101_010_1_100001011010;
      patterns[24939] = 29'b0_110000101101_011_1_000010110101;
      patterns[24940] = 29'b0_110000101101_100_1_011000010110;
      patterns[24941] = 29'b0_110000101101_101_0_101100001011;
      patterns[24942] = 29'b0_110000101101_110_0_110000101101;
      patterns[24943] = 29'b0_110000101101_111_0_110000101101;
      patterns[24944] = 29'b0_110000101110_000_0_110000101110;
      patterns[24945] = 29'b0_110000101110_001_0_101110110000;
      patterns[24946] = 29'b0_110000101110_010_1_100001011100;
      patterns[24947] = 29'b0_110000101110_011_1_000010111001;
      patterns[24948] = 29'b0_110000101110_100_0_011000010111;
      patterns[24949] = 29'b0_110000101110_101_1_001100001011;
      patterns[24950] = 29'b0_110000101110_110_0_110000101110;
      patterns[24951] = 29'b0_110000101110_111_0_110000101110;
      patterns[24952] = 29'b0_110000101111_000_0_110000101111;
      patterns[24953] = 29'b0_110000101111_001_0_101111110000;
      patterns[24954] = 29'b0_110000101111_010_1_100001011110;
      patterns[24955] = 29'b0_110000101111_011_1_000010111101;
      patterns[24956] = 29'b0_110000101111_100_1_011000010111;
      patterns[24957] = 29'b0_110000101111_101_1_101100001011;
      patterns[24958] = 29'b0_110000101111_110_0_110000101111;
      patterns[24959] = 29'b0_110000101111_111_0_110000101111;
      patterns[24960] = 29'b0_110000110000_000_0_110000110000;
      patterns[24961] = 29'b0_110000110000_001_0_110000110000;
      patterns[24962] = 29'b0_110000110000_010_1_100001100000;
      patterns[24963] = 29'b0_110000110000_011_1_000011000001;
      patterns[24964] = 29'b0_110000110000_100_0_011000011000;
      patterns[24965] = 29'b0_110000110000_101_0_001100001100;
      patterns[24966] = 29'b0_110000110000_110_0_110000110000;
      patterns[24967] = 29'b0_110000110000_111_0_110000110000;
      patterns[24968] = 29'b0_110000110001_000_0_110000110001;
      patterns[24969] = 29'b0_110000110001_001_0_110001110000;
      patterns[24970] = 29'b0_110000110001_010_1_100001100010;
      patterns[24971] = 29'b0_110000110001_011_1_000011000101;
      patterns[24972] = 29'b0_110000110001_100_1_011000011000;
      patterns[24973] = 29'b0_110000110001_101_0_101100001100;
      patterns[24974] = 29'b0_110000110001_110_0_110000110001;
      patterns[24975] = 29'b0_110000110001_111_0_110000110001;
      patterns[24976] = 29'b0_110000110010_000_0_110000110010;
      patterns[24977] = 29'b0_110000110010_001_0_110010110000;
      patterns[24978] = 29'b0_110000110010_010_1_100001100100;
      patterns[24979] = 29'b0_110000110010_011_1_000011001001;
      patterns[24980] = 29'b0_110000110010_100_0_011000011001;
      patterns[24981] = 29'b0_110000110010_101_1_001100001100;
      patterns[24982] = 29'b0_110000110010_110_0_110000110010;
      patterns[24983] = 29'b0_110000110010_111_0_110000110010;
      patterns[24984] = 29'b0_110000110011_000_0_110000110011;
      patterns[24985] = 29'b0_110000110011_001_0_110011110000;
      patterns[24986] = 29'b0_110000110011_010_1_100001100110;
      patterns[24987] = 29'b0_110000110011_011_1_000011001101;
      patterns[24988] = 29'b0_110000110011_100_1_011000011001;
      patterns[24989] = 29'b0_110000110011_101_1_101100001100;
      patterns[24990] = 29'b0_110000110011_110_0_110000110011;
      patterns[24991] = 29'b0_110000110011_111_0_110000110011;
      patterns[24992] = 29'b0_110000110100_000_0_110000110100;
      patterns[24993] = 29'b0_110000110100_001_0_110100110000;
      patterns[24994] = 29'b0_110000110100_010_1_100001101000;
      patterns[24995] = 29'b0_110000110100_011_1_000011010001;
      patterns[24996] = 29'b0_110000110100_100_0_011000011010;
      patterns[24997] = 29'b0_110000110100_101_0_001100001101;
      patterns[24998] = 29'b0_110000110100_110_0_110000110100;
      patterns[24999] = 29'b0_110000110100_111_0_110000110100;
      patterns[25000] = 29'b0_110000110101_000_0_110000110101;
      patterns[25001] = 29'b0_110000110101_001_0_110101110000;
      patterns[25002] = 29'b0_110000110101_010_1_100001101010;
      patterns[25003] = 29'b0_110000110101_011_1_000011010101;
      patterns[25004] = 29'b0_110000110101_100_1_011000011010;
      patterns[25005] = 29'b0_110000110101_101_0_101100001101;
      patterns[25006] = 29'b0_110000110101_110_0_110000110101;
      patterns[25007] = 29'b0_110000110101_111_0_110000110101;
      patterns[25008] = 29'b0_110000110110_000_0_110000110110;
      patterns[25009] = 29'b0_110000110110_001_0_110110110000;
      patterns[25010] = 29'b0_110000110110_010_1_100001101100;
      patterns[25011] = 29'b0_110000110110_011_1_000011011001;
      patterns[25012] = 29'b0_110000110110_100_0_011000011011;
      patterns[25013] = 29'b0_110000110110_101_1_001100001101;
      patterns[25014] = 29'b0_110000110110_110_0_110000110110;
      patterns[25015] = 29'b0_110000110110_111_0_110000110110;
      patterns[25016] = 29'b0_110000110111_000_0_110000110111;
      patterns[25017] = 29'b0_110000110111_001_0_110111110000;
      patterns[25018] = 29'b0_110000110111_010_1_100001101110;
      patterns[25019] = 29'b0_110000110111_011_1_000011011101;
      patterns[25020] = 29'b0_110000110111_100_1_011000011011;
      patterns[25021] = 29'b0_110000110111_101_1_101100001101;
      patterns[25022] = 29'b0_110000110111_110_0_110000110111;
      patterns[25023] = 29'b0_110000110111_111_0_110000110111;
      patterns[25024] = 29'b0_110000111000_000_0_110000111000;
      patterns[25025] = 29'b0_110000111000_001_0_111000110000;
      patterns[25026] = 29'b0_110000111000_010_1_100001110000;
      patterns[25027] = 29'b0_110000111000_011_1_000011100001;
      patterns[25028] = 29'b0_110000111000_100_0_011000011100;
      patterns[25029] = 29'b0_110000111000_101_0_001100001110;
      patterns[25030] = 29'b0_110000111000_110_0_110000111000;
      patterns[25031] = 29'b0_110000111000_111_0_110000111000;
      patterns[25032] = 29'b0_110000111001_000_0_110000111001;
      patterns[25033] = 29'b0_110000111001_001_0_111001110000;
      patterns[25034] = 29'b0_110000111001_010_1_100001110010;
      patterns[25035] = 29'b0_110000111001_011_1_000011100101;
      patterns[25036] = 29'b0_110000111001_100_1_011000011100;
      patterns[25037] = 29'b0_110000111001_101_0_101100001110;
      patterns[25038] = 29'b0_110000111001_110_0_110000111001;
      patterns[25039] = 29'b0_110000111001_111_0_110000111001;
      patterns[25040] = 29'b0_110000111010_000_0_110000111010;
      patterns[25041] = 29'b0_110000111010_001_0_111010110000;
      patterns[25042] = 29'b0_110000111010_010_1_100001110100;
      patterns[25043] = 29'b0_110000111010_011_1_000011101001;
      patterns[25044] = 29'b0_110000111010_100_0_011000011101;
      patterns[25045] = 29'b0_110000111010_101_1_001100001110;
      patterns[25046] = 29'b0_110000111010_110_0_110000111010;
      patterns[25047] = 29'b0_110000111010_111_0_110000111010;
      patterns[25048] = 29'b0_110000111011_000_0_110000111011;
      patterns[25049] = 29'b0_110000111011_001_0_111011110000;
      patterns[25050] = 29'b0_110000111011_010_1_100001110110;
      patterns[25051] = 29'b0_110000111011_011_1_000011101101;
      patterns[25052] = 29'b0_110000111011_100_1_011000011101;
      patterns[25053] = 29'b0_110000111011_101_1_101100001110;
      patterns[25054] = 29'b0_110000111011_110_0_110000111011;
      patterns[25055] = 29'b0_110000111011_111_0_110000111011;
      patterns[25056] = 29'b0_110000111100_000_0_110000111100;
      patterns[25057] = 29'b0_110000111100_001_0_111100110000;
      patterns[25058] = 29'b0_110000111100_010_1_100001111000;
      patterns[25059] = 29'b0_110000111100_011_1_000011110001;
      patterns[25060] = 29'b0_110000111100_100_0_011000011110;
      patterns[25061] = 29'b0_110000111100_101_0_001100001111;
      patterns[25062] = 29'b0_110000111100_110_0_110000111100;
      patterns[25063] = 29'b0_110000111100_111_0_110000111100;
      patterns[25064] = 29'b0_110000111101_000_0_110000111101;
      patterns[25065] = 29'b0_110000111101_001_0_111101110000;
      patterns[25066] = 29'b0_110000111101_010_1_100001111010;
      patterns[25067] = 29'b0_110000111101_011_1_000011110101;
      patterns[25068] = 29'b0_110000111101_100_1_011000011110;
      patterns[25069] = 29'b0_110000111101_101_0_101100001111;
      patterns[25070] = 29'b0_110000111101_110_0_110000111101;
      patterns[25071] = 29'b0_110000111101_111_0_110000111101;
      patterns[25072] = 29'b0_110000111110_000_0_110000111110;
      patterns[25073] = 29'b0_110000111110_001_0_111110110000;
      patterns[25074] = 29'b0_110000111110_010_1_100001111100;
      patterns[25075] = 29'b0_110000111110_011_1_000011111001;
      patterns[25076] = 29'b0_110000111110_100_0_011000011111;
      patterns[25077] = 29'b0_110000111110_101_1_001100001111;
      patterns[25078] = 29'b0_110000111110_110_0_110000111110;
      patterns[25079] = 29'b0_110000111110_111_0_110000111110;
      patterns[25080] = 29'b0_110000111111_000_0_110000111111;
      patterns[25081] = 29'b0_110000111111_001_0_111111110000;
      patterns[25082] = 29'b0_110000111111_010_1_100001111110;
      patterns[25083] = 29'b0_110000111111_011_1_000011111101;
      patterns[25084] = 29'b0_110000111111_100_1_011000011111;
      patterns[25085] = 29'b0_110000111111_101_1_101100001111;
      patterns[25086] = 29'b0_110000111111_110_0_110000111111;
      patterns[25087] = 29'b0_110000111111_111_0_110000111111;
      patterns[25088] = 29'b0_110001000000_000_0_110001000000;
      patterns[25089] = 29'b0_110001000000_001_0_000000110001;
      patterns[25090] = 29'b0_110001000000_010_1_100010000000;
      patterns[25091] = 29'b0_110001000000_011_1_000100000001;
      patterns[25092] = 29'b0_110001000000_100_0_011000100000;
      patterns[25093] = 29'b0_110001000000_101_0_001100010000;
      patterns[25094] = 29'b0_110001000000_110_0_110001000000;
      patterns[25095] = 29'b0_110001000000_111_0_110001000000;
      patterns[25096] = 29'b0_110001000001_000_0_110001000001;
      patterns[25097] = 29'b0_110001000001_001_0_000001110001;
      patterns[25098] = 29'b0_110001000001_010_1_100010000010;
      patterns[25099] = 29'b0_110001000001_011_1_000100000101;
      patterns[25100] = 29'b0_110001000001_100_1_011000100000;
      patterns[25101] = 29'b0_110001000001_101_0_101100010000;
      patterns[25102] = 29'b0_110001000001_110_0_110001000001;
      patterns[25103] = 29'b0_110001000001_111_0_110001000001;
      patterns[25104] = 29'b0_110001000010_000_0_110001000010;
      patterns[25105] = 29'b0_110001000010_001_0_000010110001;
      patterns[25106] = 29'b0_110001000010_010_1_100010000100;
      patterns[25107] = 29'b0_110001000010_011_1_000100001001;
      patterns[25108] = 29'b0_110001000010_100_0_011000100001;
      patterns[25109] = 29'b0_110001000010_101_1_001100010000;
      patterns[25110] = 29'b0_110001000010_110_0_110001000010;
      patterns[25111] = 29'b0_110001000010_111_0_110001000010;
      patterns[25112] = 29'b0_110001000011_000_0_110001000011;
      patterns[25113] = 29'b0_110001000011_001_0_000011110001;
      patterns[25114] = 29'b0_110001000011_010_1_100010000110;
      patterns[25115] = 29'b0_110001000011_011_1_000100001101;
      patterns[25116] = 29'b0_110001000011_100_1_011000100001;
      patterns[25117] = 29'b0_110001000011_101_1_101100010000;
      patterns[25118] = 29'b0_110001000011_110_0_110001000011;
      patterns[25119] = 29'b0_110001000011_111_0_110001000011;
      patterns[25120] = 29'b0_110001000100_000_0_110001000100;
      patterns[25121] = 29'b0_110001000100_001_0_000100110001;
      patterns[25122] = 29'b0_110001000100_010_1_100010001000;
      patterns[25123] = 29'b0_110001000100_011_1_000100010001;
      patterns[25124] = 29'b0_110001000100_100_0_011000100010;
      patterns[25125] = 29'b0_110001000100_101_0_001100010001;
      patterns[25126] = 29'b0_110001000100_110_0_110001000100;
      patterns[25127] = 29'b0_110001000100_111_0_110001000100;
      patterns[25128] = 29'b0_110001000101_000_0_110001000101;
      patterns[25129] = 29'b0_110001000101_001_0_000101110001;
      patterns[25130] = 29'b0_110001000101_010_1_100010001010;
      patterns[25131] = 29'b0_110001000101_011_1_000100010101;
      patterns[25132] = 29'b0_110001000101_100_1_011000100010;
      patterns[25133] = 29'b0_110001000101_101_0_101100010001;
      patterns[25134] = 29'b0_110001000101_110_0_110001000101;
      patterns[25135] = 29'b0_110001000101_111_0_110001000101;
      patterns[25136] = 29'b0_110001000110_000_0_110001000110;
      patterns[25137] = 29'b0_110001000110_001_0_000110110001;
      patterns[25138] = 29'b0_110001000110_010_1_100010001100;
      patterns[25139] = 29'b0_110001000110_011_1_000100011001;
      patterns[25140] = 29'b0_110001000110_100_0_011000100011;
      patterns[25141] = 29'b0_110001000110_101_1_001100010001;
      patterns[25142] = 29'b0_110001000110_110_0_110001000110;
      patterns[25143] = 29'b0_110001000110_111_0_110001000110;
      patterns[25144] = 29'b0_110001000111_000_0_110001000111;
      patterns[25145] = 29'b0_110001000111_001_0_000111110001;
      patterns[25146] = 29'b0_110001000111_010_1_100010001110;
      patterns[25147] = 29'b0_110001000111_011_1_000100011101;
      patterns[25148] = 29'b0_110001000111_100_1_011000100011;
      patterns[25149] = 29'b0_110001000111_101_1_101100010001;
      patterns[25150] = 29'b0_110001000111_110_0_110001000111;
      patterns[25151] = 29'b0_110001000111_111_0_110001000111;
      patterns[25152] = 29'b0_110001001000_000_0_110001001000;
      patterns[25153] = 29'b0_110001001000_001_0_001000110001;
      patterns[25154] = 29'b0_110001001000_010_1_100010010000;
      patterns[25155] = 29'b0_110001001000_011_1_000100100001;
      patterns[25156] = 29'b0_110001001000_100_0_011000100100;
      patterns[25157] = 29'b0_110001001000_101_0_001100010010;
      patterns[25158] = 29'b0_110001001000_110_0_110001001000;
      patterns[25159] = 29'b0_110001001000_111_0_110001001000;
      patterns[25160] = 29'b0_110001001001_000_0_110001001001;
      patterns[25161] = 29'b0_110001001001_001_0_001001110001;
      patterns[25162] = 29'b0_110001001001_010_1_100010010010;
      patterns[25163] = 29'b0_110001001001_011_1_000100100101;
      patterns[25164] = 29'b0_110001001001_100_1_011000100100;
      patterns[25165] = 29'b0_110001001001_101_0_101100010010;
      patterns[25166] = 29'b0_110001001001_110_0_110001001001;
      patterns[25167] = 29'b0_110001001001_111_0_110001001001;
      patterns[25168] = 29'b0_110001001010_000_0_110001001010;
      patterns[25169] = 29'b0_110001001010_001_0_001010110001;
      patterns[25170] = 29'b0_110001001010_010_1_100010010100;
      patterns[25171] = 29'b0_110001001010_011_1_000100101001;
      patterns[25172] = 29'b0_110001001010_100_0_011000100101;
      patterns[25173] = 29'b0_110001001010_101_1_001100010010;
      patterns[25174] = 29'b0_110001001010_110_0_110001001010;
      patterns[25175] = 29'b0_110001001010_111_0_110001001010;
      patterns[25176] = 29'b0_110001001011_000_0_110001001011;
      patterns[25177] = 29'b0_110001001011_001_0_001011110001;
      patterns[25178] = 29'b0_110001001011_010_1_100010010110;
      patterns[25179] = 29'b0_110001001011_011_1_000100101101;
      patterns[25180] = 29'b0_110001001011_100_1_011000100101;
      patterns[25181] = 29'b0_110001001011_101_1_101100010010;
      patterns[25182] = 29'b0_110001001011_110_0_110001001011;
      patterns[25183] = 29'b0_110001001011_111_0_110001001011;
      patterns[25184] = 29'b0_110001001100_000_0_110001001100;
      patterns[25185] = 29'b0_110001001100_001_0_001100110001;
      patterns[25186] = 29'b0_110001001100_010_1_100010011000;
      patterns[25187] = 29'b0_110001001100_011_1_000100110001;
      patterns[25188] = 29'b0_110001001100_100_0_011000100110;
      patterns[25189] = 29'b0_110001001100_101_0_001100010011;
      patterns[25190] = 29'b0_110001001100_110_0_110001001100;
      patterns[25191] = 29'b0_110001001100_111_0_110001001100;
      patterns[25192] = 29'b0_110001001101_000_0_110001001101;
      patterns[25193] = 29'b0_110001001101_001_0_001101110001;
      patterns[25194] = 29'b0_110001001101_010_1_100010011010;
      patterns[25195] = 29'b0_110001001101_011_1_000100110101;
      patterns[25196] = 29'b0_110001001101_100_1_011000100110;
      patterns[25197] = 29'b0_110001001101_101_0_101100010011;
      patterns[25198] = 29'b0_110001001101_110_0_110001001101;
      patterns[25199] = 29'b0_110001001101_111_0_110001001101;
      patterns[25200] = 29'b0_110001001110_000_0_110001001110;
      patterns[25201] = 29'b0_110001001110_001_0_001110110001;
      patterns[25202] = 29'b0_110001001110_010_1_100010011100;
      patterns[25203] = 29'b0_110001001110_011_1_000100111001;
      patterns[25204] = 29'b0_110001001110_100_0_011000100111;
      patterns[25205] = 29'b0_110001001110_101_1_001100010011;
      patterns[25206] = 29'b0_110001001110_110_0_110001001110;
      patterns[25207] = 29'b0_110001001110_111_0_110001001110;
      patterns[25208] = 29'b0_110001001111_000_0_110001001111;
      patterns[25209] = 29'b0_110001001111_001_0_001111110001;
      patterns[25210] = 29'b0_110001001111_010_1_100010011110;
      patterns[25211] = 29'b0_110001001111_011_1_000100111101;
      patterns[25212] = 29'b0_110001001111_100_1_011000100111;
      patterns[25213] = 29'b0_110001001111_101_1_101100010011;
      patterns[25214] = 29'b0_110001001111_110_0_110001001111;
      patterns[25215] = 29'b0_110001001111_111_0_110001001111;
      patterns[25216] = 29'b0_110001010000_000_0_110001010000;
      patterns[25217] = 29'b0_110001010000_001_0_010000110001;
      patterns[25218] = 29'b0_110001010000_010_1_100010100000;
      patterns[25219] = 29'b0_110001010000_011_1_000101000001;
      patterns[25220] = 29'b0_110001010000_100_0_011000101000;
      patterns[25221] = 29'b0_110001010000_101_0_001100010100;
      patterns[25222] = 29'b0_110001010000_110_0_110001010000;
      patterns[25223] = 29'b0_110001010000_111_0_110001010000;
      patterns[25224] = 29'b0_110001010001_000_0_110001010001;
      patterns[25225] = 29'b0_110001010001_001_0_010001110001;
      patterns[25226] = 29'b0_110001010001_010_1_100010100010;
      patterns[25227] = 29'b0_110001010001_011_1_000101000101;
      patterns[25228] = 29'b0_110001010001_100_1_011000101000;
      patterns[25229] = 29'b0_110001010001_101_0_101100010100;
      patterns[25230] = 29'b0_110001010001_110_0_110001010001;
      patterns[25231] = 29'b0_110001010001_111_0_110001010001;
      patterns[25232] = 29'b0_110001010010_000_0_110001010010;
      patterns[25233] = 29'b0_110001010010_001_0_010010110001;
      patterns[25234] = 29'b0_110001010010_010_1_100010100100;
      patterns[25235] = 29'b0_110001010010_011_1_000101001001;
      patterns[25236] = 29'b0_110001010010_100_0_011000101001;
      patterns[25237] = 29'b0_110001010010_101_1_001100010100;
      patterns[25238] = 29'b0_110001010010_110_0_110001010010;
      patterns[25239] = 29'b0_110001010010_111_0_110001010010;
      patterns[25240] = 29'b0_110001010011_000_0_110001010011;
      patterns[25241] = 29'b0_110001010011_001_0_010011110001;
      patterns[25242] = 29'b0_110001010011_010_1_100010100110;
      patterns[25243] = 29'b0_110001010011_011_1_000101001101;
      patterns[25244] = 29'b0_110001010011_100_1_011000101001;
      patterns[25245] = 29'b0_110001010011_101_1_101100010100;
      patterns[25246] = 29'b0_110001010011_110_0_110001010011;
      patterns[25247] = 29'b0_110001010011_111_0_110001010011;
      patterns[25248] = 29'b0_110001010100_000_0_110001010100;
      patterns[25249] = 29'b0_110001010100_001_0_010100110001;
      patterns[25250] = 29'b0_110001010100_010_1_100010101000;
      patterns[25251] = 29'b0_110001010100_011_1_000101010001;
      patterns[25252] = 29'b0_110001010100_100_0_011000101010;
      patterns[25253] = 29'b0_110001010100_101_0_001100010101;
      patterns[25254] = 29'b0_110001010100_110_0_110001010100;
      patterns[25255] = 29'b0_110001010100_111_0_110001010100;
      patterns[25256] = 29'b0_110001010101_000_0_110001010101;
      patterns[25257] = 29'b0_110001010101_001_0_010101110001;
      patterns[25258] = 29'b0_110001010101_010_1_100010101010;
      patterns[25259] = 29'b0_110001010101_011_1_000101010101;
      patterns[25260] = 29'b0_110001010101_100_1_011000101010;
      patterns[25261] = 29'b0_110001010101_101_0_101100010101;
      patterns[25262] = 29'b0_110001010101_110_0_110001010101;
      patterns[25263] = 29'b0_110001010101_111_0_110001010101;
      patterns[25264] = 29'b0_110001010110_000_0_110001010110;
      patterns[25265] = 29'b0_110001010110_001_0_010110110001;
      patterns[25266] = 29'b0_110001010110_010_1_100010101100;
      patterns[25267] = 29'b0_110001010110_011_1_000101011001;
      patterns[25268] = 29'b0_110001010110_100_0_011000101011;
      patterns[25269] = 29'b0_110001010110_101_1_001100010101;
      patterns[25270] = 29'b0_110001010110_110_0_110001010110;
      patterns[25271] = 29'b0_110001010110_111_0_110001010110;
      patterns[25272] = 29'b0_110001010111_000_0_110001010111;
      patterns[25273] = 29'b0_110001010111_001_0_010111110001;
      patterns[25274] = 29'b0_110001010111_010_1_100010101110;
      patterns[25275] = 29'b0_110001010111_011_1_000101011101;
      patterns[25276] = 29'b0_110001010111_100_1_011000101011;
      patterns[25277] = 29'b0_110001010111_101_1_101100010101;
      patterns[25278] = 29'b0_110001010111_110_0_110001010111;
      patterns[25279] = 29'b0_110001010111_111_0_110001010111;
      patterns[25280] = 29'b0_110001011000_000_0_110001011000;
      patterns[25281] = 29'b0_110001011000_001_0_011000110001;
      patterns[25282] = 29'b0_110001011000_010_1_100010110000;
      patterns[25283] = 29'b0_110001011000_011_1_000101100001;
      patterns[25284] = 29'b0_110001011000_100_0_011000101100;
      patterns[25285] = 29'b0_110001011000_101_0_001100010110;
      patterns[25286] = 29'b0_110001011000_110_0_110001011000;
      patterns[25287] = 29'b0_110001011000_111_0_110001011000;
      patterns[25288] = 29'b0_110001011001_000_0_110001011001;
      patterns[25289] = 29'b0_110001011001_001_0_011001110001;
      patterns[25290] = 29'b0_110001011001_010_1_100010110010;
      patterns[25291] = 29'b0_110001011001_011_1_000101100101;
      patterns[25292] = 29'b0_110001011001_100_1_011000101100;
      patterns[25293] = 29'b0_110001011001_101_0_101100010110;
      patterns[25294] = 29'b0_110001011001_110_0_110001011001;
      patterns[25295] = 29'b0_110001011001_111_0_110001011001;
      patterns[25296] = 29'b0_110001011010_000_0_110001011010;
      patterns[25297] = 29'b0_110001011010_001_0_011010110001;
      patterns[25298] = 29'b0_110001011010_010_1_100010110100;
      patterns[25299] = 29'b0_110001011010_011_1_000101101001;
      patterns[25300] = 29'b0_110001011010_100_0_011000101101;
      patterns[25301] = 29'b0_110001011010_101_1_001100010110;
      patterns[25302] = 29'b0_110001011010_110_0_110001011010;
      patterns[25303] = 29'b0_110001011010_111_0_110001011010;
      patterns[25304] = 29'b0_110001011011_000_0_110001011011;
      patterns[25305] = 29'b0_110001011011_001_0_011011110001;
      patterns[25306] = 29'b0_110001011011_010_1_100010110110;
      patterns[25307] = 29'b0_110001011011_011_1_000101101101;
      patterns[25308] = 29'b0_110001011011_100_1_011000101101;
      patterns[25309] = 29'b0_110001011011_101_1_101100010110;
      patterns[25310] = 29'b0_110001011011_110_0_110001011011;
      patterns[25311] = 29'b0_110001011011_111_0_110001011011;
      patterns[25312] = 29'b0_110001011100_000_0_110001011100;
      patterns[25313] = 29'b0_110001011100_001_0_011100110001;
      patterns[25314] = 29'b0_110001011100_010_1_100010111000;
      patterns[25315] = 29'b0_110001011100_011_1_000101110001;
      patterns[25316] = 29'b0_110001011100_100_0_011000101110;
      patterns[25317] = 29'b0_110001011100_101_0_001100010111;
      patterns[25318] = 29'b0_110001011100_110_0_110001011100;
      patterns[25319] = 29'b0_110001011100_111_0_110001011100;
      patterns[25320] = 29'b0_110001011101_000_0_110001011101;
      patterns[25321] = 29'b0_110001011101_001_0_011101110001;
      patterns[25322] = 29'b0_110001011101_010_1_100010111010;
      patterns[25323] = 29'b0_110001011101_011_1_000101110101;
      patterns[25324] = 29'b0_110001011101_100_1_011000101110;
      patterns[25325] = 29'b0_110001011101_101_0_101100010111;
      patterns[25326] = 29'b0_110001011101_110_0_110001011101;
      patterns[25327] = 29'b0_110001011101_111_0_110001011101;
      patterns[25328] = 29'b0_110001011110_000_0_110001011110;
      patterns[25329] = 29'b0_110001011110_001_0_011110110001;
      patterns[25330] = 29'b0_110001011110_010_1_100010111100;
      patterns[25331] = 29'b0_110001011110_011_1_000101111001;
      patterns[25332] = 29'b0_110001011110_100_0_011000101111;
      patterns[25333] = 29'b0_110001011110_101_1_001100010111;
      patterns[25334] = 29'b0_110001011110_110_0_110001011110;
      patterns[25335] = 29'b0_110001011110_111_0_110001011110;
      patterns[25336] = 29'b0_110001011111_000_0_110001011111;
      patterns[25337] = 29'b0_110001011111_001_0_011111110001;
      patterns[25338] = 29'b0_110001011111_010_1_100010111110;
      patterns[25339] = 29'b0_110001011111_011_1_000101111101;
      patterns[25340] = 29'b0_110001011111_100_1_011000101111;
      patterns[25341] = 29'b0_110001011111_101_1_101100010111;
      patterns[25342] = 29'b0_110001011111_110_0_110001011111;
      patterns[25343] = 29'b0_110001011111_111_0_110001011111;
      patterns[25344] = 29'b0_110001100000_000_0_110001100000;
      patterns[25345] = 29'b0_110001100000_001_0_100000110001;
      patterns[25346] = 29'b0_110001100000_010_1_100011000000;
      patterns[25347] = 29'b0_110001100000_011_1_000110000001;
      patterns[25348] = 29'b0_110001100000_100_0_011000110000;
      patterns[25349] = 29'b0_110001100000_101_0_001100011000;
      patterns[25350] = 29'b0_110001100000_110_0_110001100000;
      patterns[25351] = 29'b0_110001100000_111_0_110001100000;
      patterns[25352] = 29'b0_110001100001_000_0_110001100001;
      patterns[25353] = 29'b0_110001100001_001_0_100001110001;
      patterns[25354] = 29'b0_110001100001_010_1_100011000010;
      patterns[25355] = 29'b0_110001100001_011_1_000110000101;
      patterns[25356] = 29'b0_110001100001_100_1_011000110000;
      patterns[25357] = 29'b0_110001100001_101_0_101100011000;
      patterns[25358] = 29'b0_110001100001_110_0_110001100001;
      patterns[25359] = 29'b0_110001100001_111_0_110001100001;
      patterns[25360] = 29'b0_110001100010_000_0_110001100010;
      patterns[25361] = 29'b0_110001100010_001_0_100010110001;
      patterns[25362] = 29'b0_110001100010_010_1_100011000100;
      patterns[25363] = 29'b0_110001100010_011_1_000110001001;
      patterns[25364] = 29'b0_110001100010_100_0_011000110001;
      patterns[25365] = 29'b0_110001100010_101_1_001100011000;
      patterns[25366] = 29'b0_110001100010_110_0_110001100010;
      patterns[25367] = 29'b0_110001100010_111_0_110001100010;
      patterns[25368] = 29'b0_110001100011_000_0_110001100011;
      patterns[25369] = 29'b0_110001100011_001_0_100011110001;
      patterns[25370] = 29'b0_110001100011_010_1_100011000110;
      patterns[25371] = 29'b0_110001100011_011_1_000110001101;
      patterns[25372] = 29'b0_110001100011_100_1_011000110001;
      patterns[25373] = 29'b0_110001100011_101_1_101100011000;
      patterns[25374] = 29'b0_110001100011_110_0_110001100011;
      patterns[25375] = 29'b0_110001100011_111_0_110001100011;
      patterns[25376] = 29'b0_110001100100_000_0_110001100100;
      patterns[25377] = 29'b0_110001100100_001_0_100100110001;
      patterns[25378] = 29'b0_110001100100_010_1_100011001000;
      patterns[25379] = 29'b0_110001100100_011_1_000110010001;
      patterns[25380] = 29'b0_110001100100_100_0_011000110010;
      patterns[25381] = 29'b0_110001100100_101_0_001100011001;
      patterns[25382] = 29'b0_110001100100_110_0_110001100100;
      patterns[25383] = 29'b0_110001100100_111_0_110001100100;
      patterns[25384] = 29'b0_110001100101_000_0_110001100101;
      patterns[25385] = 29'b0_110001100101_001_0_100101110001;
      patterns[25386] = 29'b0_110001100101_010_1_100011001010;
      patterns[25387] = 29'b0_110001100101_011_1_000110010101;
      patterns[25388] = 29'b0_110001100101_100_1_011000110010;
      patterns[25389] = 29'b0_110001100101_101_0_101100011001;
      patterns[25390] = 29'b0_110001100101_110_0_110001100101;
      patterns[25391] = 29'b0_110001100101_111_0_110001100101;
      patterns[25392] = 29'b0_110001100110_000_0_110001100110;
      patterns[25393] = 29'b0_110001100110_001_0_100110110001;
      patterns[25394] = 29'b0_110001100110_010_1_100011001100;
      patterns[25395] = 29'b0_110001100110_011_1_000110011001;
      patterns[25396] = 29'b0_110001100110_100_0_011000110011;
      patterns[25397] = 29'b0_110001100110_101_1_001100011001;
      patterns[25398] = 29'b0_110001100110_110_0_110001100110;
      patterns[25399] = 29'b0_110001100110_111_0_110001100110;
      patterns[25400] = 29'b0_110001100111_000_0_110001100111;
      patterns[25401] = 29'b0_110001100111_001_0_100111110001;
      patterns[25402] = 29'b0_110001100111_010_1_100011001110;
      patterns[25403] = 29'b0_110001100111_011_1_000110011101;
      patterns[25404] = 29'b0_110001100111_100_1_011000110011;
      patterns[25405] = 29'b0_110001100111_101_1_101100011001;
      patterns[25406] = 29'b0_110001100111_110_0_110001100111;
      patterns[25407] = 29'b0_110001100111_111_0_110001100111;
      patterns[25408] = 29'b0_110001101000_000_0_110001101000;
      patterns[25409] = 29'b0_110001101000_001_0_101000110001;
      patterns[25410] = 29'b0_110001101000_010_1_100011010000;
      patterns[25411] = 29'b0_110001101000_011_1_000110100001;
      patterns[25412] = 29'b0_110001101000_100_0_011000110100;
      patterns[25413] = 29'b0_110001101000_101_0_001100011010;
      patterns[25414] = 29'b0_110001101000_110_0_110001101000;
      patterns[25415] = 29'b0_110001101000_111_0_110001101000;
      patterns[25416] = 29'b0_110001101001_000_0_110001101001;
      patterns[25417] = 29'b0_110001101001_001_0_101001110001;
      patterns[25418] = 29'b0_110001101001_010_1_100011010010;
      patterns[25419] = 29'b0_110001101001_011_1_000110100101;
      patterns[25420] = 29'b0_110001101001_100_1_011000110100;
      patterns[25421] = 29'b0_110001101001_101_0_101100011010;
      patterns[25422] = 29'b0_110001101001_110_0_110001101001;
      patterns[25423] = 29'b0_110001101001_111_0_110001101001;
      patterns[25424] = 29'b0_110001101010_000_0_110001101010;
      patterns[25425] = 29'b0_110001101010_001_0_101010110001;
      patterns[25426] = 29'b0_110001101010_010_1_100011010100;
      patterns[25427] = 29'b0_110001101010_011_1_000110101001;
      patterns[25428] = 29'b0_110001101010_100_0_011000110101;
      patterns[25429] = 29'b0_110001101010_101_1_001100011010;
      patterns[25430] = 29'b0_110001101010_110_0_110001101010;
      patterns[25431] = 29'b0_110001101010_111_0_110001101010;
      patterns[25432] = 29'b0_110001101011_000_0_110001101011;
      patterns[25433] = 29'b0_110001101011_001_0_101011110001;
      patterns[25434] = 29'b0_110001101011_010_1_100011010110;
      patterns[25435] = 29'b0_110001101011_011_1_000110101101;
      patterns[25436] = 29'b0_110001101011_100_1_011000110101;
      patterns[25437] = 29'b0_110001101011_101_1_101100011010;
      patterns[25438] = 29'b0_110001101011_110_0_110001101011;
      patterns[25439] = 29'b0_110001101011_111_0_110001101011;
      patterns[25440] = 29'b0_110001101100_000_0_110001101100;
      patterns[25441] = 29'b0_110001101100_001_0_101100110001;
      patterns[25442] = 29'b0_110001101100_010_1_100011011000;
      patterns[25443] = 29'b0_110001101100_011_1_000110110001;
      patterns[25444] = 29'b0_110001101100_100_0_011000110110;
      patterns[25445] = 29'b0_110001101100_101_0_001100011011;
      patterns[25446] = 29'b0_110001101100_110_0_110001101100;
      patterns[25447] = 29'b0_110001101100_111_0_110001101100;
      patterns[25448] = 29'b0_110001101101_000_0_110001101101;
      patterns[25449] = 29'b0_110001101101_001_0_101101110001;
      patterns[25450] = 29'b0_110001101101_010_1_100011011010;
      patterns[25451] = 29'b0_110001101101_011_1_000110110101;
      patterns[25452] = 29'b0_110001101101_100_1_011000110110;
      patterns[25453] = 29'b0_110001101101_101_0_101100011011;
      patterns[25454] = 29'b0_110001101101_110_0_110001101101;
      patterns[25455] = 29'b0_110001101101_111_0_110001101101;
      patterns[25456] = 29'b0_110001101110_000_0_110001101110;
      patterns[25457] = 29'b0_110001101110_001_0_101110110001;
      patterns[25458] = 29'b0_110001101110_010_1_100011011100;
      patterns[25459] = 29'b0_110001101110_011_1_000110111001;
      patterns[25460] = 29'b0_110001101110_100_0_011000110111;
      patterns[25461] = 29'b0_110001101110_101_1_001100011011;
      patterns[25462] = 29'b0_110001101110_110_0_110001101110;
      patterns[25463] = 29'b0_110001101110_111_0_110001101110;
      patterns[25464] = 29'b0_110001101111_000_0_110001101111;
      patterns[25465] = 29'b0_110001101111_001_0_101111110001;
      patterns[25466] = 29'b0_110001101111_010_1_100011011110;
      patterns[25467] = 29'b0_110001101111_011_1_000110111101;
      patterns[25468] = 29'b0_110001101111_100_1_011000110111;
      patterns[25469] = 29'b0_110001101111_101_1_101100011011;
      patterns[25470] = 29'b0_110001101111_110_0_110001101111;
      patterns[25471] = 29'b0_110001101111_111_0_110001101111;
      patterns[25472] = 29'b0_110001110000_000_0_110001110000;
      patterns[25473] = 29'b0_110001110000_001_0_110000110001;
      patterns[25474] = 29'b0_110001110000_010_1_100011100000;
      patterns[25475] = 29'b0_110001110000_011_1_000111000001;
      patterns[25476] = 29'b0_110001110000_100_0_011000111000;
      patterns[25477] = 29'b0_110001110000_101_0_001100011100;
      patterns[25478] = 29'b0_110001110000_110_0_110001110000;
      patterns[25479] = 29'b0_110001110000_111_0_110001110000;
      patterns[25480] = 29'b0_110001110001_000_0_110001110001;
      patterns[25481] = 29'b0_110001110001_001_0_110001110001;
      patterns[25482] = 29'b0_110001110001_010_1_100011100010;
      patterns[25483] = 29'b0_110001110001_011_1_000111000101;
      patterns[25484] = 29'b0_110001110001_100_1_011000111000;
      patterns[25485] = 29'b0_110001110001_101_0_101100011100;
      patterns[25486] = 29'b0_110001110001_110_0_110001110001;
      patterns[25487] = 29'b0_110001110001_111_0_110001110001;
      patterns[25488] = 29'b0_110001110010_000_0_110001110010;
      patterns[25489] = 29'b0_110001110010_001_0_110010110001;
      patterns[25490] = 29'b0_110001110010_010_1_100011100100;
      patterns[25491] = 29'b0_110001110010_011_1_000111001001;
      patterns[25492] = 29'b0_110001110010_100_0_011000111001;
      patterns[25493] = 29'b0_110001110010_101_1_001100011100;
      patterns[25494] = 29'b0_110001110010_110_0_110001110010;
      patterns[25495] = 29'b0_110001110010_111_0_110001110010;
      patterns[25496] = 29'b0_110001110011_000_0_110001110011;
      patterns[25497] = 29'b0_110001110011_001_0_110011110001;
      patterns[25498] = 29'b0_110001110011_010_1_100011100110;
      patterns[25499] = 29'b0_110001110011_011_1_000111001101;
      patterns[25500] = 29'b0_110001110011_100_1_011000111001;
      patterns[25501] = 29'b0_110001110011_101_1_101100011100;
      patterns[25502] = 29'b0_110001110011_110_0_110001110011;
      patterns[25503] = 29'b0_110001110011_111_0_110001110011;
      patterns[25504] = 29'b0_110001110100_000_0_110001110100;
      patterns[25505] = 29'b0_110001110100_001_0_110100110001;
      patterns[25506] = 29'b0_110001110100_010_1_100011101000;
      patterns[25507] = 29'b0_110001110100_011_1_000111010001;
      patterns[25508] = 29'b0_110001110100_100_0_011000111010;
      patterns[25509] = 29'b0_110001110100_101_0_001100011101;
      patterns[25510] = 29'b0_110001110100_110_0_110001110100;
      patterns[25511] = 29'b0_110001110100_111_0_110001110100;
      patterns[25512] = 29'b0_110001110101_000_0_110001110101;
      patterns[25513] = 29'b0_110001110101_001_0_110101110001;
      patterns[25514] = 29'b0_110001110101_010_1_100011101010;
      patterns[25515] = 29'b0_110001110101_011_1_000111010101;
      patterns[25516] = 29'b0_110001110101_100_1_011000111010;
      patterns[25517] = 29'b0_110001110101_101_0_101100011101;
      patterns[25518] = 29'b0_110001110101_110_0_110001110101;
      patterns[25519] = 29'b0_110001110101_111_0_110001110101;
      patterns[25520] = 29'b0_110001110110_000_0_110001110110;
      patterns[25521] = 29'b0_110001110110_001_0_110110110001;
      patterns[25522] = 29'b0_110001110110_010_1_100011101100;
      patterns[25523] = 29'b0_110001110110_011_1_000111011001;
      patterns[25524] = 29'b0_110001110110_100_0_011000111011;
      patterns[25525] = 29'b0_110001110110_101_1_001100011101;
      patterns[25526] = 29'b0_110001110110_110_0_110001110110;
      patterns[25527] = 29'b0_110001110110_111_0_110001110110;
      patterns[25528] = 29'b0_110001110111_000_0_110001110111;
      patterns[25529] = 29'b0_110001110111_001_0_110111110001;
      patterns[25530] = 29'b0_110001110111_010_1_100011101110;
      patterns[25531] = 29'b0_110001110111_011_1_000111011101;
      patterns[25532] = 29'b0_110001110111_100_1_011000111011;
      patterns[25533] = 29'b0_110001110111_101_1_101100011101;
      patterns[25534] = 29'b0_110001110111_110_0_110001110111;
      patterns[25535] = 29'b0_110001110111_111_0_110001110111;
      patterns[25536] = 29'b0_110001111000_000_0_110001111000;
      patterns[25537] = 29'b0_110001111000_001_0_111000110001;
      patterns[25538] = 29'b0_110001111000_010_1_100011110000;
      patterns[25539] = 29'b0_110001111000_011_1_000111100001;
      patterns[25540] = 29'b0_110001111000_100_0_011000111100;
      patterns[25541] = 29'b0_110001111000_101_0_001100011110;
      patterns[25542] = 29'b0_110001111000_110_0_110001111000;
      patterns[25543] = 29'b0_110001111000_111_0_110001111000;
      patterns[25544] = 29'b0_110001111001_000_0_110001111001;
      patterns[25545] = 29'b0_110001111001_001_0_111001110001;
      patterns[25546] = 29'b0_110001111001_010_1_100011110010;
      patterns[25547] = 29'b0_110001111001_011_1_000111100101;
      patterns[25548] = 29'b0_110001111001_100_1_011000111100;
      patterns[25549] = 29'b0_110001111001_101_0_101100011110;
      patterns[25550] = 29'b0_110001111001_110_0_110001111001;
      patterns[25551] = 29'b0_110001111001_111_0_110001111001;
      patterns[25552] = 29'b0_110001111010_000_0_110001111010;
      patterns[25553] = 29'b0_110001111010_001_0_111010110001;
      patterns[25554] = 29'b0_110001111010_010_1_100011110100;
      patterns[25555] = 29'b0_110001111010_011_1_000111101001;
      patterns[25556] = 29'b0_110001111010_100_0_011000111101;
      patterns[25557] = 29'b0_110001111010_101_1_001100011110;
      patterns[25558] = 29'b0_110001111010_110_0_110001111010;
      patterns[25559] = 29'b0_110001111010_111_0_110001111010;
      patterns[25560] = 29'b0_110001111011_000_0_110001111011;
      patterns[25561] = 29'b0_110001111011_001_0_111011110001;
      patterns[25562] = 29'b0_110001111011_010_1_100011110110;
      patterns[25563] = 29'b0_110001111011_011_1_000111101101;
      patterns[25564] = 29'b0_110001111011_100_1_011000111101;
      patterns[25565] = 29'b0_110001111011_101_1_101100011110;
      patterns[25566] = 29'b0_110001111011_110_0_110001111011;
      patterns[25567] = 29'b0_110001111011_111_0_110001111011;
      patterns[25568] = 29'b0_110001111100_000_0_110001111100;
      patterns[25569] = 29'b0_110001111100_001_0_111100110001;
      patterns[25570] = 29'b0_110001111100_010_1_100011111000;
      patterns[25571] = 29'b0_110001111100_011_1_000111110001;
      patterns[25572] = 29'b0_110001111100_100_0_011000111110;
      patterns[25573] = 29'b0_110001111100_101_0_001100011111;
      patterns[25574] = 29'b0_110001111100_110_0_110001111100;
      patterns[25575] = 29'b0_110001111100_111_0_110001111100;
      patterns[25576] = 29'b0_110001111101_000_0_110001111101;
      patterns[25577] = 29'b0_110001111101_001_0_111101110001;
      patterns[25578] = 29'b0_110001111101_010_1_100011111010;
      patterns[25579] = 29'b0_110001111101_011_1_000111110101;
      patterns[25580] = 29'b0_110001111101_100_1_011000111110;
      patterns[25581] = 29'b0_110001111101_101_0_101100011111;
      patterns[25582] = 29'b0_110001111101_110_0_110001111101;
      patterns[25583] = 29'b0_110001111101_111_0_110001111101;
      patterns[25584] = 29'b0_110001111110_000_0_110001111110;
      patterns[25585] = 29'b0_110001111110_001_0_111110110001;
      patterns[25586] = 29'b0_110001111110_010_1_100011111100;
      patterns[25587] = 29'b0_110001111110_011_1_000111111001;
      patterns[25588] = 29'b0_110001111110_100_0_011000111111;
      patterns[25589] = 29'b0_110001111110_101_1_001100011111;
      patterns[25590] = 29'b0_110001111110_110_0_110001111110;
      patterns[25591] = 29'b0_110001111110_111_0_110001111110;
      patterns[25592] = 29'b0_110001111111_000_0_110001111111;
      patterns[25593] = 29'b0_110001111111_001_0_111111110001;
      patterns[25594] = 29'b0_110001111111_010_1_100011111110;
      patterns[25595] = 29'b0_110001111111_011_1_000111111101;
      patterns[25596] = 29'b0_110001111111_100_1_011000111111;
      patterns[25597] = 29'b0_110001111111_101_1_101100011111;
      patterns[25598] = 29'b0_110001111111_110_0_110001111111;
      patterns[25599] = 29'b0_110001111111_111_0_110001111111;
      patterns[25600] = 29'b0_110010000000_000_0_110010000000;
      patterns[25601] = 29'b0_110010000000_001_0_000000110010;
      patterns[25602] = 29'b0_110010000000_010_1_100100000000;
      patterns[25603] = 29'b0_110010000000_011_1_001000000001;
      patterns[25604] = 29'b0_110010000000_100_0_011001000000;
      patterns[25605] = 29'b0_110010000000_101_0_001100100000;
      patterns[25606] = 29'b0_110010000000_110_0_110010000000;
      patterns[25607] = 29'b0_110010000000_111_0_110010000000;
      patterns[25608] = 29'b0_110010000001_000_0_110010000001;
      patterns[25609] = 29'b0_110010000001_001_0_000001110010;
      patterns[25610] = 29'b0_110010000001_010_1_100100000010;
      patterns[25611] = 29'b0_110010000001_011_1_001000000101;
      patterns[25612] = 29'b0_110010000001_100_1_011001000000;
      patterns[25613] = 29'b0_110010000001_101_0_101100100000;
      patterns[25614] = 29'b0_110010000001_110_0_110010000001;
      patterns[25615] = 29'b0_110010000001_111_0_110010000001;
      patterns[25616] = 29'b0_110010000010_000_0_110010000010;
      patterns[25617] = 29'b0_110010000010_001_0_000010110010;
      patterns[25618] = 29'b0_110010000010_010_1_100100000100;
      patterns[25619] = 29'b0_110010000010_011_1_001000001001;
      patterns[25620] = 29'b0_110010000010_100_0_011001000001;
      patterns[25621] = 29'b0_110010000010_101_1_001100100000;
      patterns[25622] = 29'b0_110010000010_110_0_110010000010;
      patterns[25623] = 29'b0_110010000010_111_0_110010000010;
      patterns[25624] = 29'b0_110010000011_000_0_110010000011;
      patterns[25625] = 29'b0_110010000011_001_0_000011110010;
      patterns[25626] = 29'b0_110010000011_010_1_100100000110;
      patterns[25627] = 29'b0_110010000011_011_1_001000001101;
      patterns[25628] = 29'b0_110010000011_100_1_011001000001;
      patterns[25629] = 29'b0_110010000011_101_1_101100100000;
      patterns[25630] = 29'b0_110010000011_110_0_110010000011;
      patterns[25631] = 29'b0_110010000011_111_0_110010000011;
      patterns[25632] = 29'b0_110010000100_000_0_110010000100;
      patterns[25633] = 29'b0_110010000100_001_0_000100110010;
      patterns[25634] = 29'b0_110010000100_010_1_100100001000;
      patterns[25635] = 29'b0_110010000100_011_1_001000010001;
      patterns[25636] = 29'b0_110010000100_100_0_011001000010;
      patterns[25637] = 29'b0_110010000100_101_0_001100100001;
      patterns[25638] = 29'b0_110010000100_110_0_110010000100;
      patterns[25639] = 29'b0_110010000100_111_0_110010000100;
      patterns[25640] = 29'b0_110010000101_000_0_110010000101;
      patterns[25641] = 29'b0_110010000101_001_0_000101110010;
      patterns[25642] = 29'b0_110010000101_010_1_100100001010;
      patterns[25643] = 29'b0_110010000101_011_1_001000010101;
      patterns[25644] = 29'b0_110010000101_100_1_011001000010;
      patterns[25645] = 29'b0_110010000101_101_0_101100100001;
      patterns[25646] = 29'b0_110010000101_110_0_110010000101;
      patterns[25647] = 29'b0_110010000101_111_0_110010000101;
      patterns[25648] = 29'b0_110010000110_000_0_110010000110;
      patterns[25649] = 29'b0_110010000110_001_0_000110110010;
      patterns[25650] = 29'b0_110010000110_010_1_100100001100;
      patterns[25651] = 29'b0_110010000110_011_1_001000011001;
      patterns[25652] = 29'b0_110010000110_100_0_011001000011;
      patterns[25653] = 29'b0_110010000110_101_1_001100100001;
      patterns[25654] = 29'b0_110010000110_110_0_110010000110;
      patterns[25655] = 29'b0_110010000110_111_0_110010000110;
      patterns[25656] = 29'b0_110010000111_000_0_110010000111;
      patterns[25657] = 29'b0_110010000111_001_0_000111110010;
      patterns[25658] = 29'b0_110010000111_010_1_100100001110;
      patterns[25659] = 29'b0_110010000111_011_1_001000011101;
      patterns[25660] = 29'b0_110010000111_100_1_011001000011;
      patterns[25661] = 29'b0_110010000111_101_1_101100100001;
      patterns[25662] = 29'b0_110010000111_110_0_110010000111;
      patterns[25663] = 29'b0_110010000111_111_0_110010000111;
      patterns[25664] = 29'b0_110010001000_000_0_110010001000;
      patterns[25665] = 29'b0_110010001000_001_0_001000110010;
      patterns[25666] = 29'b0_110010001000_010_1_100100010000;
      patterns[25667] = 29'b0_110010001000_011_1_001000100001;
      patterns[25668] = 29'b0_110010001000_100_0_011001000100;
      patterns[25669] = 29'b0_110010001000_101_0_001100100010;
      patterns[25670] = 29'b0_110010001000_110_0_110010001000;
      patterns[25671] = 29'b0_110010001000_111_0_110010001000;
      patterns[25672] = 29'b0_110010001001_000_0_110010001001;
      patterns[25673] = 29'b0_110010001001_001_0_001001110010;
      patterns[25674] = 29'b0_110010001001_010_1_100100010010;
      patterns[25675] = 29'b0_110010001001_011_1_001000100101;
      patterns[25676] = 29'b0_110010001001_100_1_011001000100;
      patterns[25677] = 29'b0_110010001001_101_0_101100100010;
      patterns[25678] = 29'b0_110010001001_110_0_110010001001;
      patterns[25679] = 29'b0_110010001001_111_0_110010001001;
      patterns[25680] = 29'b0_110010001010_000_0_110010001010;
      patterns[25681] = 29'b0_110010001010_001_0_001010110010;
      patterns[25682] = 29'b0_110010001010_010_1_100100010100;
      patterns[25683] = 29'b0_110010001010_011_1_001000101001;
      patterns[25684] = 29'b0_110010001010_100_0_011001000101;
      patterns[25685] = 29'b0_110010001010_101_1_001100100010;
      patterns[25686] = 29'b0_110010001010_110_0_110010001010;
      patterns[25687] = 29'b0_110010001010_111_0_110010001010;
      patterns[25688] = 29'b0_110010001011_000_0_110010001011;
      patterns[25689] = 29'b0_110010001011_001_0_001011110010;
      patterns[25690] = 29'b0_110010001011_010_1_100100010110;
      patterns[25691] = 29'b0_110010001011_011_1_001000101101;
      patterns[25692] = 29'b0_110010001011_100_1_011001000101;
      patterns[25693] = 29'b0_110010001011_101_1_101100100010;
      patterns[25694] = 29'b0_110010001011_110_0_110010001011;
      patterns[25695] = 29'b0_110010001011_111_0_110010001011;
      patterns[25696] = 29'b0_110010001100_000_0_110010001100;
      patterns[25697] = 29'b0_110010001100_001_0_001100110010;
      patterns[25698] = 29'b0_110010001100_010_1_100100011000;
      patterns[25699] = 29'b0_110010001100_011_1_001000110001;
      patterns[25700] = 29'b0_110010001100_100_0_011001000110;
      patterns[25701] = 29'b0_110010001100_101_0_001100100011;
      patterns[25702] = 29'b0_110010001100_110_0_110010001100;
      patterns[25703] = 29'b0_110010001100_111_0_110010001100;
      patterns[25704] = 29'b0_110010001101_000_0_110010001101;
      patterns[25705] = 29'b0_110010001101_001_0_001101110010;
      patterns[25706] = 29'b0_110010001101_010_1_100100011010;
      patterns[25707] = 29'b0_110010001101_011_1_001000110101;
      patterns[25708] = 29'b0_110010001101_100_1_011001000110;
      patterns[25709] = 29'b0_110010001101_101_0_101100100011;
      patterns[25710] = 29'b0_110010001101_110_0_110010001101;
      patterns[25711] = 29'b0_110010001101_111_0_110010001101;
      patterns[25712] = 29'b0_110010001110_000_0_110010001110;
      patterns[25713] = 29'b0_110010001110_001_0_001110110010;
      patterns[25714] = 29'b0_110010001110_010_1_100100011100;
      patterns[25715] = 29'b0_110010001110_011_1_001000111001;
      patterns[25716] = 29'b0_110010001110_100_0_011001000111;
      patterns[25717] = 29'b0_110010001110_101_1_001100100011;
      patterns[25718] = 29'b0_110010001110_110_0_110010001110;
      patterns[25719] = 29'b0_110010001110_111_0_110010001110;
      patterns[25720] = 29'b0_110010001111_000_0_110010001111;
      patterns[25721] = 29'b0_110010001111_001_0_001111110010;
      patterns[25722] = 29'b0_110010001111_010_1_100100011110;
      patterns[25723] = 29'b0_110010001111_011_1_001000111101;
      patterns[25724] = 29'b0_110010001111_100_1_011001000111;
      patterns[25725] = 29'b0_110010001111_101_1_101100100011;
      patterns[25726] = 29'b0_110010001111_110_0_110010001111;
      patterns[25727] = 29'b0_110010001111_111_0_110010001111;
      patterns[25728] = 29'b0_110010010000_000_0_110010010000;
      patterns[25729] = 29'b0_110010010000_001_0_010000110010;
      patterns[25730] = 29'b0_110010010000_010_1_100100100000;
      patterns[25731] = 29'b0_110010010000_011_1_001001000001;
      patterns[25732] = 29'b0_110010010000_100_0_011001001000;
      patterns[25733] = 29'b0_110010010000_101_0_001100100100;
      patterns[25734] = 29'b0_110010010000_110_0_110010010000;
      patterns[25735] = 29'b0_110010010000_111_0_110010010000;
      patterns[25736] = 29'b0_110010010001_000_0_110010010001;
      patterns[25737] = 29'b0_110010010001_001_0_010001110010;
      patterns[25738] = 29'b0_110010010001_010_1_100100100010;
      patterns[25739] = 29'b0_110010010001_011_1_001001000101;
      patterns[25740] = 29'b0_110010010001_100_1_011001001000;
      patterns[25741] = 29'b0_110010010001_101_0_101100100100;
      patterns[25742] = 29'b0_110010010001_110_0_110010010001;
      patterns[25743] = 29'b0_110010010001_111_0_110010010001;
      patterns[25744] = 29'b0_110010010010_000_0_110010010010;
      patterns[25745] = 29'b0_110010010010_001_0_010010110010;
      patterns[25746] = 29'b0_110010010010_010_1_100100100100;
      patterns[25747] = 29'b0_110010010010_011_1_001001001001;
      patterns[25748] = 29'b0_110010010010_100_0_011001001001;
      patterns[25749] = 29'b0_110010010010_101_1_001100100100;
      patterns[25750] = 29'b0_110010010010_110_0_110010010010;
      patterns[25751] = 29'b0_110010010010_111_0_110010010010;
      patterns[25752] = 29'b0_110010010011_000_0_110010010011;
      patterns[25753] = 29'b0_110010010011_001_0_010011110010;
      patterns[25754] = 29'b0_110010010011_010_1_100100100110;
      patterns[25755] = 29'b0_110010010011_011_1_001001001101;
      patterns[25756] = 29'b0_110010010011_100_1_011001001001;
      patterns[25757] = 29'b0_110010010011_101_1_101100100100;
      patterns[25758] = 29'b0_110010010011_110_0_110010010011;
      patterns[25759] = 29'b0_110010010011_111_0_110010010011;
      patterns[25760] = 29'b0_110010010100_000_0_110010010100;
      patterns[25761] = 29'b0_110010010100_001_0_010100110010;
      patterns[25762] = 29'b0_110010010100_010_1_100100101000;
      patterns[25763] = 29'b0_110010010100_011_1_001001010001;
      patterns[25764] = 29'b0_110010010100_100_0_011001001010;
      patterns[25765] = 29'b0_110010010100_101_0_001100100101;
      patterns[25766] = 29'b0_110010010100_110_0_110010010100;
      patterns[25767] = 29'b0_110010010100_111_0_110010010100;
      patterns[25768] = 29'b0_110010010101_000_0_110010010101;
      patterns[25769] = 29'b0_110010010101_001_0_010101110010;
      patterns[25770] = 29'b0_110010010101_010_1_100100101010;
      patterns[25771] = 29'b0_110010010101_011_1_001001010101;
      patterns[25772] = 29'b0_110010010101_100_1_011001001010;
      patterns[25773] = 29'b0_110010010101_101_0_101100100101;
      patterns[25774] = 29'b0_110010010101_110_0_110010010101;
      patterns[25775] = 29'b0_110010010101_111_0_110010010101;
      patterns[25776] = 29'b0_110010010110_000_0_110010010110;
      patterns[25777] = 29'b0_110010010110_001_0_010110110010;
      patterns[25778] = 29'b0_110010010110_010_1_100100101100;
      patterns[25779] = 29'b0_110010010110_011_1_001001011001;
      patterns[25780] = 29'b0_110010010110_100_0_011001001011;
      patterns[25781] = 29'b0_110010010110_101_1_001100100101;
      patterns[25782] = 29'b0_110010010110_110_0_110010010110;
      patterns[25783] = 29'b0_110010010110_111_0_110010010110;
      patterns[25784] = 29'b0_110010010111_000_0_110010010111;
      patterns[25785] = 29'b0_110010010111_001_0_010111110010;
      patterns[25786] = 29'b0_110010010111_010_1_100100101110;
      patterns[25787] = 29'b0_110010010111_011_1_001001011101;
      patterns[25788] = 29'b0_110010010111_100_1_011001001011;
      patterns[25789] = 29'b0_110010010111_101_1_101100100101;
      patterns[25790] = 29'b0_110010010111_110_0_110010010111;
      patterns[25791] = 29'b0_110010010111_111_0_110010010111;
      patterns[25792] = 29'b0_110010011000_000_0_110010011000;
      patterns[25793] = 29'b0_110010011000_001_0_011000110010;
      patterns[25794] = 29'b0_110010011000_010_1_100100110000;
      patterns[25795] = 29'b0_110010011000_011_1_001001100001;
      patterns[25796] = 29'b0_110010011000_100_0_011001001100;
      patterns[25797] = 29'b0_110010011000_101_0_001100100110;
      patterns[25798] = 29'b0_110010011000_110_0_110010011000;
      patterns[25799] = 29'b0_110010011000_111_0_110010011000;
      patterns[25800] = 29'b0_110010011001_000_0_110010011001;
      patterns[25801] = 29'b0_110010011001_001_0_011001110010;
      patterns[25802] = 29'b0_110010011001_010_1_100100110010;
      patterns[25803] = 29'b0_110010011001_011_1_001001100101;
      patterns[25804] = 29'b0_110010011001_100_1_011001001100;
      patterns[25805] = 29'b0_110010011001_101_0_101100100110;
      patterns[25806] = 29'b0_110010011001_110_0_110010011001;
      patterns[25807] = 29'b0_110010011001_111_0_110010011001;
      patterns[25808] = 29'b0_110010011010_000_0_110010011010;
      patterns[25809] = 29'b0_110010011010_001_0_011010110010;
      patterns[25810] = 29'b0_110010011010_010_1_100100110100;
      patterns[25811] = 29'b0_110010011010_011_1_001001101001;
      patterns[25812] = 29'b0_110010011010_100_0_011001001101;
      patterns[25813] = 29'b0_110010011010_101_1_001100100110;
      patterns[25814] = 29'b0_110010011010_110_0_110010011010;
      patterns[25815] = 29'b0_110010011010_111_0_110010011010;
      patterns[25816] = 29'b0_110010011011_000_0_110010011011;
      patterns[25817] = 29'b0_110010011011_001_0_011011110010;
      patterns[25818] = 29'b0_110010011011_010_1_100100110110;
      patterns[25819] = 29'b0_110010011011_011_1_001001101101;
      patterns[25820] = 29'b0_110010011011_100_1_011001001101;
      patterns[25821] = 29'b0_110010011011_101_1_101100100110;
      patterns[25822] = 29'b0_110010011011_110_0_110010011011;
      patterns[25823] = 29'b0_110010011011_111_0_110010011011;
      patterns[25824] = 29'b0_110010011100_000_0_110010011100;
      patterns[25825] = 29'b0_110010011100_001_0_011100110010;
      patterns[25826] = 29'b0_110010011100_010_1_100100111000;
      patterns[25827] = 29'b0_110010011100_011_1_001001110001;
      patterns[25828] = 29'b0_110010011100_100_0_011001001110;
      patterns[25829] = 29'b0_110010011100_101_0_001100100111;
      patterns[25830] = 29'b0_110010011100_110_0_110010011100;
      patterns[25831] = 29'b0_110010011100_111_0_110010011100;
      patterns[25832] = 29'b0_110010011101_000_0_110010011101;
      patterns[25833] = 29'b0_110010011101_001_0_011101110010;
      patterns[25834] = 29'b0_110010011101_010_1_100100111010;
      patterns[25835] = 29'b0_110010011101_011_1_001001110101;
      patterns[25836] = 29'b0_110010011101_100_1_011001001110;
      patterns[25837] = 29'b0_110010011101_101_0_101100100111;
      patterns[25838] = 29'b0_110010011101_110_0_110010011101;
      patterns[25839] = 29'b0_110010011101_111_0_110010011101;
      patterns[25840] = 29'b0_110010011110_000_0_110010011110;
      patterns[25841] = 29'b0_110010011110_001_0_011110110010;
      patterns[25842] = 29'b0_110010011110_010_1_100100111100;
      patterns[25843] = 29'b0_110010011110_011_1_001001111001;
      patterns[25844] = 29'b0_110010011110_100_0_011001001111;
      patterns[25845] = 29'b0_110010011110_101_1_001100100111;
      patterns[25846] = 29'b0_110010011110_110_0_110010011110;
      patterns[25847] = 29'b0_110010011110_111_0_110010011110;
      patterns[25848] = 29'b0_110010011111_000_0_110010011111;
      patterns[25849] = 29'b0_110010011111_001_0_011111110010;
      patterns[25850] = 29'b0_110010011111_010_1_100100111110;
      patterns[25851] = 29'b0_110010011111_011_1_001001111101;
      patterns[25852] = 29'b0_110010011111_100_1_011001001111;
      patterns[25853] = 29'b0_110010011111_101_1_101100100111;
      patterns[25854] = 29'b0_110010011111_110_0_110010011111;
      patterns[25855] = 29'b0_110010011111_111_0_110010011111;
      patterns[25856] = 29'b0_110010100000_000_0_110010100000;
      patterns[25857] = 29'b0_110010100000_001_0_100000110010;
      patterns[25858] = 29'b0_110010100000_010_1_100101000000;
      patterns[25859] = 29'b0_110010100000_011_1_001010000001;
      patterns[25860] = 29'b0_110010100000_100_0_011001010000;
      patterns[25861] = 29'b0_110010100000_101_0_001100101000;
      patterns[25862] = 29'b0_110010100000_110_0_110010100000;
      patterns[25863] = 29'b0_110010100000_111_0_110010100000;
      patterns[25864] = 29'b0_110010100001_000_0_110010100001;
      patterns[25865] = 29'b0_110010100001_001_0_100001110010;
      patterns[25866] = 29'b0_110010100001_010_1_100101000010;
      patterns[25867] = 29'b0_110010100001_011_1_001010000101;
      patterns[25868] = 29'b0_110010100001_100_1_011001010000;
      patterns[25869] = 29'b0_110010100001_101_0_101100101000;
      patterns[25870] = 29'b0_110010100001_110_0_110010100001;
      patterns[25871] = 29'b0_110010100001_111_0_110010100001;
      patterns[25872] = 29'b0_110010100010_000_0_110010100010;
      patterns[25873] = 29'b0_110010100010_001_0_100010110010;
      patterns[25874] = 29'b0_110010100010_010_1_100101000100;
      patterns[25875] = 29'b0_110010100010_011_1_001010001001;
      patterns[25876] = 29'b0_110010100010_100_0_011001010001;
      patterns[25877] = 29'b0_110010100010_101_1_001100101000;
      patterns[25878] = 29'b0_110010100010_110_0_110010100010;
      patterns[25879] = 29'b0_110010100010_111_0_110010100010;
      patterns[25880] = 29'b0_110010100011_000_0_110010100011;
      patterns[25881] = 29'b0_110010100011_001_0_100011110010;
      patterns[25882] = 29'b0_110010100011_010_1_100101000110;
      patterns[25883] = 29'b0_110010100011_011_1_001010001101;
      patterns[25884] = 29'b0_110010100011_100_1_011001010001;
      patterns[25885] = 29'b0_110010100011_101_1_101100101000;
      patterns[25886] = 29'b0_110010100011_110_0_110010100011;
      patterns[25887] = 29'b0_110010100011_111_0_110010100011;
      patterns[25888] = 29'b0_110010100100_000_0_110010100100;
      patterns[25889] = 29'b0_110010100100_001_0_100100110010;
      patterns[25890] = 29'b0_110010100100_010_1_100101001000;
      patterns[25891] = 29'b0_110010100100_011_1_001010010001;
      patterns[25892] = 29'b0_110010100100_100_0_011001010010;
      patterns[25893] = 29'b0_110010100100_101_0_001100101001;
      patterns[25894] = 29'b0_110010100100_110_0_110010100100;
      patterns[25895] = 29'b0_110010100100_111_0_110010100100;
      patterns[25896] = 29'b0_110010100101_000_0_110010100101;
      patterns[25897] = 29'b0_110010100101_001_0_100101110010;
      patterns[25898] = 29'b0_110010100101_010_1_100101001010;
      patterns[25899] = 29'b0_110010100101_011_1_001010010101;
      patterns[25900] = 29'b0_110010100101_100_1_011001010010;
      patterns[25901] = 29'b0_110010100101_101_0_101100101001;
      patterns[25902] = 29'b0_110010100101_110_0_110010100101;
      patterns[25903] = 29'b0_110010100101_111_0_110010100101;
      patterns[25904] = 29'b0_110010100110_000_0_110010100110;
      patterns[25905] = 29'b0_110010100110_001_0_100110110010;
      patterns[25906] = 29'b0_110010100110_010_1_100101001100;
      patterns[25907] = 29'b0_110010100110_011_1_001010011001;
      patterns[25908] = 29'b0_110010100110_100_0_011001010011;
      patterns[25909] = 29'b0_110010100110_101_1_001100101001;
      patterns[25910] = 29'b0_110010100110_110_0_110010100110;
      patterns[25911] = 29'b0_110010100110_111_0_110010100110;
      patterns[25912] = 29'b0_110010100111_000_0_110010100111;
      patterns[25913] = 29'b0_110010100111_001_0_100111110010;
      patterns[25914] = 29'b0_110010100111_010_1_100101001110;
      patterns[25915] = 29'b0_110010100111_011_1_001010011101;
      patterns[25916] = 29'b0_110010100111_100_1_011001010011;
      patterns[25917] = 29'b0_110010100111_101_1_101100101001;
      patterns[25918] = 29'b0_110010100111_110_0_110010100111;
      patterns[25919] = 29'b0_110010100111_111_0_110010100111;
      patterns[25920] = 29'b0_110010101000_000_0_110010101000;
      patterns[25921] = 29'b0_110010101000_001_0_101000110010;
      patterns[25922] = 29'b0_110010101000_010_1_100101010000;
      patterns[25923] = 29'b0_110010101000_011_1_001010100001;
      patterns[25924] = 29'b0_110010101000_100_0_011001010100;
      patterns[25925] = 29'b0_110010101000_101_0_001100101010;
      patterns[25926] = 29'b0_110010101000_110_0_110010101000;
      patterns[25927] = 29'b0_110010101000_111_0_110010101000;
      patterns[25928] = 29'b0_110010101001_000_0_110010101001;
      patterns[25929] = 29'b0_110010101001_001_0_101001110010;
      patterns[25930] = 29'b0_110010101001_010_1_100101010010;
      patterns[25931] = 29'b0_110010101001_011_1_001010100101;
      patterns[25932] = 29'b0_110010101001_100_1_011001010100;
      patterns[25933] = 29'b0_110010101001_101_0_101100101010;
      patterns[25934] = 29'b0_110010101001_110_0_110010101001;
      patterns[25935] = 29'b0_110010101001_111_0_110010101001;
      patterns[25936] = 29'b0_110010101010_000_0_110010101010;
      patterns[25937] = 29'b0_110010101010_001_0_101010110010;
      patterns[25938] = 29'b0_110010101010_010_1_100101010100;
      patterns[25939] = 29'b0_110010101010_011_1_001010101001;
      patterns[25940] = 29'b0_110010101010_100_0_011001010101;
      patterns[25941] = 29'b0_110010101010_101_1_001100101010;
      patterns[25942] = 29'b0_110010101010_110_0_110010101010;
      patterns[25943] = 29'b0_110010101010_111_0_110010101010;
      patterns[25944] = 29'b0_110010101011_000_0_110010101011;
      patterns[25945] = 29'b0_110010101011_001_0_101011110010;
      patterns[25946] = 29'b0_110010101011_010_1_100101010110;
      patterns[25947] = 29'b0_110010101011_011_1_001010101101;
      patterns[25948] = 29'b0_110010101011_100_1_011001010101;
      patterns[25949] = 29'b0_110010101011_101_1_101100101010;
      patterns[25950] = 29'b0_110010101011_110_0_110010101011;
      patterns[25951] = 29'b0_110010101011_111_0_110010101011;
      patterns[25952] = 29'b0_110010101100_000_0_110010101100;
      patterns[25953] = 29'b0_110010101100_001_0_101100110010;
      patterns[25954] = 29'b0_110010101100_010_1_100101011000;
      patterns[25955] = 29'b0_110010101100_011_1_001010110001;
      patterns[25956] = 29'b0_110010101100_100_0_011001010110;
      patterns[25957] = 29'b0_110010101100_101_0_001100101011;
      patterns[25958] = 29'b0_110010101100_110_0_110010101100;
      patterns[25959] = 29'b0_110010101100_111_0_110010101100;
      patterns[25960] = 29'b0_110010101101_000_0_110010101101;
      patterns[25961] = 29'b0_110010101101_001_0_101101110010;
      patterns[25962] = 29'b0_110010101101_010_1_100101011010;
      patterns[25963] = 29'b0_110010101101_011_1_001010110101;
      patterns[25964] = 29'b0_110010101101_100_1_011001010110;
      patterns[25965] = 29'b0_110010101101_101_0_101100101011;
      patterns[25966] = 29'b0_110010101101_110_0_110010101101;
      patterns[25967] = 29'b0_110010101101_111_0_110010101101;
      patterns[25968] = 29'b0_110010101110_000_0_110010101110;
      patterns[25969] = 29'b0_110010101110_001_0_101110110010;
      patterns[25970] = 29'b0_110010101110_010_1_100101011100;
      patterns[25971] = 29'b0_110010101110_011_1_001010111001;
      patterns[25972] = 29'b0_110010101110_100_0_011001010111;
      patterns[25973] = 29'b0_110010101110_101_1_001100101011;
      patterns[25974] = 29'b0_110010101110_110_0_110010101110;
      patterns[25975] = 29'b0_110010101110_111_0_110010101110;
      patterns[25976] = 29'b0_110010101111_000_0_110010101111;
      patterns[25977] = 29'b0_110010101111_001_0_101111110010;
      patterns[25978] = 29'b0_110010101111_010_1_100101011110;
      patterns[25979] = 29'b0_110010101111_011_1_001010111101;
      patterns[25980] = 29'b0_110010101111_100_1_011001010111;
      patterns[25981] = 29'b0_110010101111_101_1_101100101011;
      patterns[25982] = 29'b0_110010101111_110_0_110010101111;
      patterns[25983] = 29'b0_110010101111_111_0_110010101111;
      patterns[25984] = 29'b0_110010110000_000_0_110010110000;
      patterns[25985] = 29'b0_110010110000_001_0_110000110010;
      patterns[25986] = 29'b0_110010110000_010_1_100101100000;
      patterns[25987] = 29'b0_110010110000_011_1_001011000001;
      patterns[25988] = 29'b0_110010110000_100_0_011001011000;
      patterns[25989] = 29'b0_110010110000_101_0_001100101100;
      patterns[25990] = 29'b0_110010110000_110_0_110010110000;
      patterns[25991] = 29'b0_110010110000_111_0_110010110000;
      patterns[25992] = 29'b0_110010110001_000_0_110010110001;
      patterns[25993] = 29'b0_110010110001_001_0_110001110010;
      patterns[25994] = 29'b0_110010110001_010_1_100101100010;
      patterns[25995] = 29'b0_110010110001_011_1_001011000101;
      patterns[25996] = 29'b0_110010110001_100_1_011001011000;
      patterns[25997] = 29'b0_110010110001_101_0_101100101100;
      patterns[25998] = 29'b0_110010110001_110_0_110010110001;
      patterns[25999] = 29'b0_110010110001_111_0_110010110001;
      patterns[26000] = 29'b0_110010110010_000_0_110010110010;
      patterns[26001] = 29'b0_110010110010_001_0_110010110010;
      patterns[26002] = 29'b0_110010110010_010_1_100101100100;
      patterns[26003] = 29'b0_110010110010_011_1_001011001001;
      patterns[26004] = 29'b0_110010110010_100_0_011001011001;
      patterns[26005] = 29'b0_110010110010_101_1_001100101100;
      patterns[26006] = 29'b0_110010110010_110_0_110010110010;
      patterns[26007] = 29'b0_110010110010_111_0_110010110010;
      patterns[26008] = 29'b0_110010110011_000_0_110010110011;
      patterns[26009] = 29'b0_110010110011_001_0_110011110010;
      patterns[26010] = 29'b0_110010110011_010_1_100101100110;
      patterns[26011] = 29'b0_110010110011_011_1_001011001101;
      patterns[26012] = 29'b0_110010110011_100_1_011001011001;
      patterns[26013] = 29'b0_110010110011_101_1_101100101100;
      patterns[26014] = 29'b0_110010110011_110_0_110010110011;
      patterns[26015] = 29'b0_110010110011_111_0_110010110011;
      patterns[26016] = 29'b0_110010110100_000_0_110010110100;
      patterns[26017] = 29'b0_110010110100_001_0_110100110010;
      patterns[26018] = 29'b0_110010110100_010_1_100101101000;
      patterns[26019] = 29'b0_110010110100_011_1_001011010001;
      patterns[26020] = 29'b0_110010110100_100_0_011001011010;
      patterns[26021] = 29'b0_110010110100_101_0_001100101101;
      patterns[26022] = 29'b0_110010110100_110_0_110010110100;
      patterns[26023] = 29'b0_110010110100_111_0_110010110100;
      patterns[26024] = 29'b0_110010110101_000_0_110010110101;
      patterns[26025] = 29'b0_110010110101_001_0_110101110010;
      patterns[26026] = 29'b0_110010110101_010_1_100101101010;
      patterns[26027] = 29'b0_110010110101_011_1_001011010101;
      patterns[26028] = 29'b0_110010110101_100_1_011001011010;
      patterns[26029] = 29'b0_110010110101_101_0_101100101101;
      patterns[26030] = 29'b0_110010110101_110_0_110010110101;
      patterns[26031] = 29'b0_110010110101_111_0_110010110101;
      patterns[26032] = 29'b0_110010110110_000_0_110010110110;
      patterns[26033] = 29'b0_110010110110_001_0_110110110010;
      patterns[26034] = 29'b0_110010110110_010_1_100101101100;
      patterns[26035] = 29'b0_110010110110_011_1_001011011001;
      patterns[26036] = 29'b0_110010110110_100_0_011001011011;
      patterns[26037] = 29'b0_110010110110_101_1_001100101101;
      patterns[26038] = 29'b0_110010110110_110_0_110010110110;
      patterns[26039] = 29'b0_110010110110_111_0_110010110110;
      patterns[26040] = 29'b0_110010110111_000_0_110010110111;
      patterns[26041] = 29'b0_110010110111_001_0_110111110010;
      patterns[26042] = 29'b0_110010110111_010_1_100101101110;
      patterns[26043] = 29'b0_110010110111_011_1_001011011101;
      patterns[26044] = 29'b0_110010110111_100_1_011001011011;
      patterns[26045] = 29'b0_110010110111_101_1_101100101101;
      patterns[26046] = 29'b0_110010110111_110_0_110010110111;
      patterns[26047] = 29'b0_110010110111_111_0_110010110111;
      patterns[26048] = 29'b0_110010111000_000_0_110010111000;
      patterns[26049] = 29'b0_110010111000_001_0_111000110010;
      patterns[26050] = 29'b0_110010111000_010_1_100101110000;
      patterns[26051] = 29'b0_110010111000_011_1_001011100001;
      patterns[26052] = 29'b0_110010111000_100_0_011001011100;
      patterns[26053] = 29'b0_110010111000_101_0_001100101110;
      patterns[26054] = 29'b0_110010111000_110_0_110010111000;
      patterns[26055] = 29'b0_110010111000_111_0_110010111000;
      patterns[26056] = 29'b0_110010111001_000_0_110010111001;
      patterns[26057] = 29'b0_110010111001_001_0_111001110010;
      patterns[26058] = 29'b0_110010111001_010_1_100101110010;
      patterns[26059] = 29'b0_110010111001_011_1_001011100101;
      patterns[26060] = 29'b0_110010111001_100_1_011001011100;
      patterns[26061] = 29'b0_110010111001_101_0_101100101110;
      patterns[26062] = 29'b0_110010111001_110_0_110010111001;
      patterns[26063] = 29'b0_110010111001_111_0_110010111001;
      patterns[26064] = 29'b0_110010111010_000_0_110010111010;
      patterns[26065] = 29'b0_110010111010_001_0_111010110010;
      patterns[26066] = 29'b0_110010111010_010_1_100101110100;
      patterns[26067] = 29'b0_110010111010_011_1_001011101001;
      patterns[26068] = 29'b0_110010111010_100_0_011001011101;
      patterns[26069] = 29'b0_110010111010_101_1_001100101110;
      patterns[26070] = 29'b0_110010111010_110_0_110010111010;
      patterns[26071] = 29'b0_110010111010_111_0_110010111010;
      patterns[26072] = 29'b0_110010111011_000_0_110010111011;
      patterns[26073] = 29'b0_110010111011_001_0_111011110010;
      patterns[26074] = 29'b0_110010111011_010_1_100101110110;
      patterns[26075] = 29'b0_110010111011_011_1_001011101101;
      patterns[26076] = 29'b0_110010111011_100_1_011001011101;
      patterns[26077] = 29'b0_110010111011_101_1_101100101110;
      patterns[26078] = 29'b0_110010111011_110_0_110010111011;
      patterns[26079] = 29'b0_110010111011_111_0_110010111011;
      patterns[26080] = 29'b0_110010111100_000_0_110010111100;
      patterns[26081] = 29'b0_110010111100_001_0_111100110010;
      patterns[26082] = 29'b0_110010111100_010_1_100101111000;
      patterns[26083] = 29'b0_110010111100_011_1_001011110001;
      patterns[26084] = 29'b0_110010111100_100_0_011001011110;
      patterns[26085] = 29'b0_110010111100_101_0_001100101111;
      patterns[26086] = 29'b0_110010111100_110_0_110010111100;
      patterns[26087] = 29'b0_110010111100_111_0_110010111100;
      patterns[26088] = 29'b0_110010111101_000_0_110010111101;
      patterns[26089] = 29'b0_110010111101_001_0_111101110010;
      patterns[26090] = 29'b0_110010111101_010_1_100101111010;
      patterns[26091] = 29'b0_110010111101_011_1_001011110101;
      patterns[26092] = 29'b0_110010111101_100_1_011001011110;
      patterns[26093] = 29'b0_110010111101_101_0_101100101111;
      patterns[26094] = 29'b0_110010111101_110_0_110010111101;
      patterns[26095] = 29'b0_110010111101_111_0_110010111101;
      patterns[26096] = 29'b0_110010111110_000_0_110010111110;
      patterns[26097] = 29'b0_110010111110_001_0_111110110010;
      patterns[26098] = 29'b0_110010111110_010_1_100101111100;
      patterns[26099] = 29'b0_110010111110_011_1_001011111001;
      patterns[26100] = 29'b0_110010111110_100_0_011001011111;
      patterns[26101] = 29'b0_110010111110_101_1_001100101111;
      patterns[26102] = 29'b0_110010111110_110_0_110010111110;
      patterns[26103] = 29'b0_110010111110_111_0_110010111110;
      patterns[26104] = 29'b0_110010111111_000_0_110010111111;
      patterns[26105] = 29'b0_110010111111_001_0_111111110010;
      patterns[26106] = 29'b0_110010111111_010_1_100101111110;
      patterns[26107] = 29'b0_110010111111_011_1_001011111101;
      patterns[26108] = 29'b0_110010111111_100_1_011001011111;
      patterns[26109] = 29'b0_110010111111_101_1_101100101111;
      patterns[26110] = 29'b0_110010111111_110_0_110010111111;
      patterns[26111] = 29'b0_110010111111_111_0_110010111111;
      patterns[26112] = 29'b0_110011000000_000_0_110011000000;
      patterns[26113] = 29'b0_110011000000_001_0_000000110011;
      patterns[26114] = 29'b0_110011000000_010_1_100110000000;
      patterns[26115] = 29'b0_110011000000_011_1_001100000001;
      patterns[26116] = 29'b0_110011000000_100_0_011001100000;
      patterns[26117] = 29'b0_110011000000_101_0_001100110000;
      patterns[26118] = 29'b0_110011000000_110_0_110011000000;
      patterns[26119] = 29'b0_110011000000_111_0_110011000000;
      patterns[26120] = 29'b0_110011000001_000_0_110011000001;
      patterns[26121] = 29'b0_110011000001_001_0_000001110011;
      patterns[26122] = 29'b0_110011000001_010_1_100110000010;
      patterns[26123] = 29'b0_110011000001_011_1_001100000101;
      patterns[26124] = 29'b0_110011000001_100_1_011001100000;
      patterns[26125] = 29'b0_110011000001_101_0_101100110000;
      patterns[26126] = 29'b0_110011000001_110_0_110011000001;
      patterns[26127] = 29'b0_110011000001_111_0_110011000001;
      patterns[26128] = 29'b0_110011000010_000_0_110011000010;
      patterns[26129] = 29'b0_110011000010_001_0_000010110011;
      patterns[26130] = 29'b0_110011000010_010_1_100110000100;
      patterns[26131] = 29'b0_110011000010_011_1_001100001001;
      patterns[26132] = 29'b0_110011000010_100_0_011001100001;
      patterns[26133] = 29'b0_110011000010_101_1_001100110000;
      patterns[26134] = 29'b0_110011000010_110_0_110011000010;
      patterns[26135] = 29'b0_110011000010_111_0_110011000010;
      patterns[26136] = 29'b0_110011000011_000_0_110011000011;
      patterns[26137] = 29'b0_110011000011_001_0_000011110011;
      patterns[26138] = 29'b0_110011000011_010_1_100110000110;
      patterns[26139] = 29'b0_110011000011_011_1_001100001101;
      patterns[26140] = 29'b0_110011000011_100_1_011001100001;
      patterns[26141] = 29'b0_110011000011_101_1_101100110000;
      patterns[26142] = 29'b0_110011000011_110_0_110011000011;
      patterns[26143] = 29'b0_110011000011_111_0_110011000011;
      patterns[26144] = 29'b0_110011000100_000_0_110011000100;
      patterns[26145] = 29'b0_110011000100_001_0_000100110011;
      patterns[26146] = 29'b0_110011000100_010_1_100110001000;
      patterns[26147] = 29'b0_110011000100_011_1_001100010001;
      patterns[26148] = 29'b0_110011000100_100_0_011001100010;
      patterns[26149] = 29'b0_110011000100_101_0_001100110001;
      patterns[26150] = 29'b0_110011000100_110_0_110011000100;
      patterns[26151] = 29'b0_110011000100_111_0_110011000100;
      patterns[26152] = 29'b0_110011000101_000_0_110011000101;
      patterns[26153] = 29'b0_110011000101_001_0_000101110011;
      patterns[26154] = 29'b0_110011000101_010_1_100110001010;
      patterns[26155] = 29'b0_110011000101_011_1_001100010101;
      patterns[26156] = 29'b0_110011000101_100_1_011001100010;
      patterns[26157] = 29'b0_110011000101_101_0_101100110001;
      patterns[26158] = 29'b0_110011000101_110_0_110011000101;
      patterns[26159] = 29'b0_110011000101_111_0_110011000101;
      patterns[26160] = 29'b0_110011000110_000_0_110011000110;
      patterns[26161] = 29'b0_110011000110_001_0_000110110011;
      patterns[26162] = 29'b0_110011000110_010_1_100110001100;
      patterns[26163] = 29'b0_110011000110_011_1_001100011001;
      patterns[26164] = 29'b0_110011000110_100_0_011001100011;
      patterns[26165] = 29'b0_110011000110_101_1_001100110001;
      patterns[26166] = 29'b0_110011000110_110_0_110011000110;
      patterns[26167] = 29'b0_110011000110_111_0_110011000110;
      patterns[26168] = 29'b0_110011000111_000_0_110011000111;
      patterns[26169] = 29'b0_110011000111_001_0_000111110011;
      patterns[26170] = 29'b0_110011000111_010_1_100110001110;
      patterns[26171] = 29'b0_110011000111_011_1_001100011101;
      patterns[26172] = 29'b0_110011000111_100_1_011001100011;
      patterns[26173] = 29'b0_110011000111_101_1_101100110001;
      patterns[26174] = 29'b0_110011000111_110_0_110011000111;
      patterns[26175] = 29'b0_110011000111_111_0_110011000111;
      patterns[26176] = 29'b0_110011001000_000_0_110011001000;
      patterns[26177] = 29'b0_110011001000_001_0_001000110011;
      patterns[26178] = 29'b0_110011001000_010_1_100110010000;
      patterns[26179] = 29'b0_110011001000_011_1_001100100001;
      patterns[26180] = 29'b0_110011001000_100_0_011001100100;
      patterns[26181] = 29'b0_110011001000_101_0_001100110010;
      patterns[26182] = 29'b0_110011001000_110_0_110011001000;
      patterns[26183] = 29'b0_110011001000_111_0_110011001000;
      patterns[26184] = 29'b0_110011001001_000_0_110011001001;
      patterns[26185] = 29'b0_110011001001_001_0_001001110011;
      patterns[26186] = 29'b0_110011001001_010_1_100110010010;
      patterns[26187] = 29'b0_110011001001_011_1_001100100101;
      patterns[26188] = 29'b0_110011001001_100_1_011001100100;
      patterns[26189] = 29'b0_110011001001_101_0_101100110010;
      patterns[26190] = 29'b0_110011001001_110_0_110011001001;
      patterns[26191] = 29'b0_110011001001_111_0_110011001001;
      patterns[26192] = 29'b0_110011001010_000_0_110011001010;
      patterns[26193] = 29'b0_110011001010_001_0_001010110011;
      patterns[26194] = 29'b0_110011001010_010_1_100110010100;
      patterns[26195] = 29'b0_110011001010_011_1_001100101001;
      patterns[26196] = 29'b0_110011001010_100_0_011001100101;
      patterns[26197] = 29'b0_110011001010_101_1_001100110010;
      patterns[26198] = 29'b0_110011001010_110_0_110011001010;
      patterns[26199] = 29'b0_110011001010_111_0_110011001010;
      patterns[26200] = 29'b0_110011001011_000_0_110011001011;
      patterns[26201] = 29'b0_110011001011_001_0_001011110011;
      patterns[26202] = 29'b0_110011001011_010_1_100110010110;
      patterns[26203] = 29'b0_110011001011_011_1_001100101101;
      patterns[26204] = 29'b0_110011001011_100_1_011001100101;
      patterns[26205] = 29'b0_110011001011_101_1_101100110010;
      patterns[26206] = 29'b0_110011001011_110_0_110011001011;
      patterns[26207] = 29'b0_110011001011_111_0_110011001011;
      patterns[26208] = 29'b0_110011001100_000_0_110011001100;
      patterns[26209] = 29'b0_110011001100_001_0_001100110011;
      patterns[26210] = 29'b0_110011001100_010_1_100110011000;
      patterns[26211] = 29'b0_110011001100_011_1_001100110001;
      patterns[26212] = 29'b0_110011001100_100_0_011001100110;
      patterns[26213] = 29'b0_110011001100_101_0_001100110011;
      patterns[26214] = 29'b0_110011001100_110_0_110011001100;
      patterns[26215] = 29'b0_110011001100_111_0_110011001100;
      patterns[26216] = 29'b0_110011001101_000_0_110011001101;
      patterns[26217] = 29'b0_110011001101_001_0_001101110011;
      patterns[26218] = 29'b0_110011001101_010_1_100110011010;
      patterns[26219] = 29'b0_110011001101_011_1_001100110101;
      patterns[26220] = 29'b0_110011001101_100_1_011001100110;
      patterns[26221] = 29'b0_110011001101_101_0_101100110011;
      patterns[26222] = 29'b0_110011001101_110_0_110011001101;
      patterns[26223] = 29'b0_110011001101_111_0_110011001101;
      patterns[26224] = 29'b0_110011001110_000_0_110011001110;
      patterns[26225] = 29'b0_110011001110_001_0_001110110011;
      patterns[26226] = 29'b0_110011001110_010_1_100110011100;
      patterns[26227] = 29'b0_110011001110_011_1_001100111001;
      patterns[26228] = 29'b0_110011001110_100_0_011001100111;
      patterns[26229] = 29'b0_110011001110_101_1_001100110011;
      patterns[26230] = 29'b0_110011001110_110_0_110011001110;
      patterns[26231] = 29'b0_110011001110_111_0_110011001110;
      patterns[26232] = 29'b0_110011001111_000_0_110011001111;
      patterns[26233] = 29'b0_110011001111_001_0_001111110011;
      patterns[26234] = 29'b0_110011001111_010_1_100110011110;
      patterns[26235] = 29'b0_110011001111_011_1_001100111101;
      patterns[26236] = 29'b0_110011001111_100_1_011001100111;
      patterns[26237] = 29'b0_110011001111_101_1_101100110011;
      patterns[26238] = 29'b0_110011001111_110_0_110011001111;
      patterns[26239] = 29'b0_110011001111_111_0_110011001111;
      patterns[26240] = 29'b0_110011010000_000_0_110011010000;
      patterns[26241] = 29'b0_110011010000_001_0_010000110011;
      patterns[26242] = 29'b0_110011010000_010_1_100110100000;
      patterns[26243] = 29'b0_110011010000_011_1_001101000001;
      patterns[26244] = 29'b0_110011010000_100_0_011001101000;
      patterns[26245] = 29'b0_110011010000_101_0_001100110100;
      patterns[26246] = 29'b0_110011010000_110_0_110011010000;
      patterns[26247] = 29'b0_110011010000_111_0_110011010000;
      patterns[26248] = 29'b0_110011010001_000_0_110011010001;
      patterns[26249] = 29'b0_110011010001_001_0_010001110011;
      patterns[26250] = 29'b0_110011010001_010_1_100110100010;
      patterns[26251] = 29'b0_110011010001_011_1_001101000101;
      patterns[26252] = 29'b0_110011010001_100_1_011001101000;
      patterns[26253] = 29'b0_110011010001_101_0_101100110100;
      patterns[26254] = 29'b0_110011010001_110_0_110011010001;
      patterns[26255] = 29'b0_110011010001_111_0_110011010001;
      patterns[26256] = 29'b0_110011010010_000_0_110011010010;
      patterns[26257] = 29'b0_110011010010_001_0_010010110011;
      patterns[26258] = 29'b0_110011010010_010_1_100110100100;
      patterns[26259] = 29'b0_110011010010_011_1_001101001001;
      patterns[26260] = 29'b0_110011010010_100_0_011001101001;
      patterns[26261] = 29'b0_110011010010_101_1_001100110100;
      patterns[26262] = 29'b0_110011010010_110_0_110011010010;
      patterns[26263] = 29'b0_110011010010_111_0_110011010010;
      patterns[26264] = 29'b0_110011010011_000_0_110011010011;
      patterns[26265] = 29'b0_110011010011_001_0_010011110011;
      patterns[26266] = 29'b0_110011010011_010_1_100110100110;
      patterns[26267] = 29'b0_110011010011_011_1_001101001101;
      patterns[26268] = 29'b0_110011010011_100_1_011001101001;
      patterns[26269] = 29'b0_110011010011_101_1_101100110100;
      patterns[26270] = 29'b0_110011010011_110_0_110011010011;
      patterns[26271] = 29'b0_110011010011_111_0_110011010011;
      patterns[26272] = 29'b0_110011010100_000_0_110011010100;
      patterns[26273] = 29'b0_110011010100_001_0_010100110011;
      patterns[26274] = 29'b0_110011010100_010_1_100110101000;
      patterns[26275] = 29'b0_110011010100_011_1_001101010001;
      patterns[26276] = 29'b0_110011010100_100_0_011001101010;
      patterns[26277] = 29'b0_110011010100_101_0_001100110101;
      patterns[26278] = 29'b0_110011010100_110_0_110011010100;
      patterns[26279] = 29'b0_110011010100_111_0_110011010100;
      patterns[26280] = 29'b0_110011010101_000_0_110011010101;
      patterns[26281] = 29'b0_110011010101_001_0_010101110011;
      patterns[26282] = 29'b0_110011010101_010_1_100110101010;
      patterns[26283] = 29'b0_110011010101_011_1_001101010101;
      patterns[26284] = 29'b0_110011010101_100_1_011001101010;
      patterns[26285] = 29'b0_110011010101_101_0_101100110101;
      patterns[26286] = 29'b0_110011010101_110_0_110011010101;
      patterns[26287] = 29'b0_110011010101_111_0_110011010101;
      patterns[26288] = 29'b0_110011010110_000_0_110011010110;
      patterns[26289] = 29'b0_110011010110_001_0_010110110011;
      patterns[26290] = 29'b0_110011010110_010_1_100110101100;
      patterns[26291] = 29'b0_110011010110_011_1_001101011001;
      patterns[26292] = 29'b0_110011010110_100_0_011001101011;
      patterns[26293] = 29'b0_110011010110_101_1_001100110101;
      patterns[26294] = 29'b0_110011010110_110_0_110011010110;
      patterns[26295] = 29'b0_110011010110_111_0_110011010110;
      patterns[26296] = 29'b0_110011010111_000_0_110011010111;
      patterns[26297] = 29'b0_110011010111_001_0_010111110011;
      patterns[26298] = 29'b0_110011010111_010_1_100110101110;
      patterns[26299] = 29'b0_110011010111_011_1_001101011101;
      patterns[26300] = 29'b0_110011010111_100_1_011001101011;
      patterns[26301] = 29'b0_110011010111_101_1_101100110101;
      patterns[26302] = 29'b0_110011010111_110_0_110011010111;
      patterns[26303] = 29'b0_110011010111_111_0_110011010111;
      patterns[26304] = 29'b0_110011011000_000_0_110011011000;
      patterns[26305] = 29'b0_110011011000_001_0_011000110011;
      patterns[26306] = 29'b0_110011011000_010_1_100110110000;
      patterns[26307] = 29'b0_110011011000_011_1_001101100001;
      patterns[26308] = 29'b0_110011011000_100_0_011001101100;
      patterns[26309] = 29'b0_110011011000_101_0_001100110110;
      patterns[26310] = 29'b0_110011011000_110_0_110011011000;
      patterns[26311] = 29'b0_110011011000_111_0_110011011000;
      patterns[26312] = 29'b0_110011011001_000_0_110011011001;
      patterns[26313] = 29'b0_110011011001_001_0_011001110011;
      patterns[26314] = 29'b0_110011011001_010_1_100110110010;
      patterns[26315] = 29'b0_110011011001_011_1_001101100101;
      patterns[26316] = 29'b0_110011011001_100_1_011001101100;
      patterns[26317] = 29'b0_110011011001_101_0_101100110110;
      patterns[26318] = 29'b0_110011011001_110_0_110011011001;
      patterns[26319] = 29'b0_110011011001_111_0_110011011001;
      patterns[26320] = 29'b0_110011011010_000_0_110011011010;
      patterns[26321] = 29'b0_110011011010_001_0_011010110011;
      patterns[26322] = 29'b0_110011011010_010_1_100110110100;
      patterns[26323] = 29'b0_110011011010_011_1_001101101001;
      patterns[26324] = 29'b0_110011011010_100_0_011001101101;
      patterns[26325] = 29'b0_110011011010_101_1_001100110110;
      patterns[26326] = 29'b0_110011011010_110_0_110011011010;
      patterns[26327] = 29'b0_110011011010_111_0_110011011010;
      patterns[26328] = 29'b0_110011011011_000_0_110011011011;
      patterns[26329] = 29'b0_110011011011_001_0_011011110011;
      patterns[26330] = 29'b0_110011011011_010_1_100110110110;
      patterns[26331] = 29'b0_110011011011_011_1_001101101101;
      patterns[26332] = 29'b0_110011011011_100_1_011001101101;
      patterns[26333] = 29'b0_110011011011_101_1_101100110110;
      patterns[26334] = 29'b0_110011011011_110_0_110011011011;
      patterns[26335] = 29'b0_110011011011_111_0_110011011011;
      patterns[26336] = 29'b0_110011011100_000_0_110011011100;
      patterns[26337] = 29'b0_110011011100_001_0_011100110011;
      patterns[26338] = 29'b0_110011011100_010_1_100110111000;
      patterns[26339] = 29'b0_110011011100_011_1_001101110001;
      patterns[26340] = 29'b0_110011011100_100_0_011001101110;
      patterns[26341] = 29'b0_110011011100_101_0_001100110111;
      patterns[26342] = 29'b0_110011011100_110_0_110011011100;
      patterns[26343] = 29'b0_110011011100_111_0_110011011100;
      patterns[26344] = 29'b0_110011011101_000_0_110011011101;
      patterns[26345] = 29'b0_110011011101_001_0_011101110011;
      patterns[26346] = 29'b0_110011011101_010_1_100110111010;
      patterns[26347] = 29'b0_110011011101_011_1_001101110101;
      patterns[26348] = 29'b0_110011011101_100_1_011001101110;
      patterns[26349] = 29'b0_110011011101_101_0_101100110111;
      patterns[26350] = 29'b0_110011011101_110_0_110011011101;
      patterns[26351] = 29'b0_110011011101_111_0_110011011101;
      patterns[26352] = 29'b0_110011011110_000_0_110011011110;
      patterns[26353] = 29'b0_110011011110_001_0_011110110011;
      patterns[26354] = 29'b0_110011011110_010_1_100110111100;
      patterns[26355] = 29'b0_110011011110_011_1_001101111001;
      patterns[26356] = 29'b0_110011011110_100_0_011001101111;
      patterns[26357] = 29'b0_110011011110_101_1_001100110111;
      patterns[26358] = 29'b0_110011011110_110_0_110011011110;
      patterns[26359] = 29'b0_110011011110_111_0_110011011110;
      patterns[26360] = 29'b0_110011011111_000_0_110011011111;
      patterns[26361] = 29'b0_110011011111_001_0_011111110011;
      patterns[26362] = 29'b0_110011011111_010_1_100110111110;
      patterns[26363] = 29'b0_110011011111_011_1_001101111101;
      patterns[26364] = 29'b0_110011011111_100_1_011001101111;
      patterns[26365] = 29'b0_110011011111_101_1_101100110111;
      patterns[26366] = 29'b0_110011011111_110_0_110011011111;
      patterns[26367] = 29'b0_110011011111_111_0_110011011111;
      patterns[26368] = 29'b0_110011100000_000_0_110011100000;
      patterns[26369] = 29'b0_110011100000_001_0_100000110011;
      patterns[26370] = 29'b0_110011100000_010_1_100111000000;
      patterns[26371] = 29'b0_110011100000_011_1_001110000001;
      patterns[26372] = 29'b0_110011100000_100_0_011001110000;
      patterns[26373] = 29'b0_110011100000_101_0_001100111000;
      patterns[26374] = 29'b0_110011100000_110_0_110011100000;
      patterns[26375] = 29'b0_110011100000_111_0_110011100000;
      patterns[26376] = 29'b0_110011100001_000_0_110011100001;
      patterns[26377] = 29'b0_110011100001_001_0_100001110011;
      patterns[26378] = 29'b0_110011100001_010_1_100111000010;
      patterns[26379] = 29'b0_110011100001_011_1_001110000101;
      patterns[26380] = 29'b0_110011100001_100_1_011001110000;
      patterns[26381] = 29'b0_110011100001_101_0_101100111000;
      patterns[26382] = 29'b0_110011100001_110_0_110011100001;
      patterns[26383] = 29'b0_110011100001_111_0_110011100001;
      patterns[26384] = 29'b0_110011100010_000_0_110011100010;
      patterns[26385] = 29'b0_110011100010_001_0_100010110011;
      patterns[26386] = 29'b0_110011100010_010_1_100111000100;
      patterns[26387] = 29'b0_110011100010_011_1_001110001001;
      patterns[26388] = 29'b0_110011100010_100_0_011001110001;
      patterns[26389] = 29'b0_110011100010_101_1_001100111000;
      patterns[26390] = 29'b0_110011100010_110_0_110011100010;
      patterns[26391] = 29'b0_110011100010_111_0_110011100010;
      patterns[26392] = 29'b0_110011100011_000_0_110011100011;
      patterns[26393] = 29'b0_110011100011_001_0_100011110011;
      patterns[26394] = 29'b0_110011100011_010_1_100111000110;
      patterns[26395] = 29'b0_110011100011_011_1_001110001101;
      patterns[26396] = 29'b0_110011100011_100_1_011001110001;
      patterns[26397] = 29'b0_110011100011_101_1_101100111000;
      patterns[26398] = 29'b0_110011100011_110_0_110011100011;
      patterns[26399] = 29'b0_110011100011_111_0_110011100011;
      patterns[26400] = 29'b0_110011100100_000_0_110011100100;
      patterns[26401] = 29'b0_110011100100_001_0_100100110011;
      patterns[26402] = 29'b0_110011100100_010_1_100111001000;
      patterns[26403] = 29'b0_110011100100_011_1_001110010001;
      patterns[26404] = 29'b0_110011100100_100_0_011001110010;
      patterns[26405] = 29'b0_110011100100_101_0_001100111001;
      patterns[26406] = 29'b0_110011100100_110_0_110011100100;
      patterns[26407] = 29'b0_110011100100_111_0_110011100100;
      patterns[26408] = 29'b0_110011100101_000_0_110011100101;
      patterns[26409] = 29'b0_110011100101_001_0_100101110011;
      patterns[26410] = 29'b0_110011100101_010_1_100111001010;
      patterns[26411] = 29'b0_110011100101_011_1_001110010101;
      patterns[26412] = 29'b0_110011100101_100_1_011001110010;
      patterns[26413] = 29'b0_110011100101_101_0_101100111001;
      patterns[26414] = 29'b0_110011100101_110_0_110011100101;
      patterns[26415] = 29'b0_110011100101_111_0_110011100101;
      patterns[26416] = 29'b0_110011100110_000_0_110011100110;
      patterns[26417] = 29'b0_110011100110_001_0_100110110011;
      patterns[26418] = 29'b0_110011100110_010_1_100111001100;
      patterns[26419] = 29'b0_110011100110_011_1_001110011001;
      patterns[26420] = 29'b0_110011100110_100_0_011001110011;
      patterns[26421] = 29'b0_110011100110_101_1_001100111001;
      patterns[26422] = 29'b0_110011100110_110_0_110011100110;
      patterns[26423] = 29'b0_110011100110_111_0_110011100110;
      patterns[26424] = 29'b0_110011100111_000_0_110011100111;
      patterns[26425] = 29'b0_110011100111_001_0_100111110011;
      patterns[26426] = 29'b0_110011100111_010_1_100111001110;
      patterns[26427] = 29'b0_110011100111_011_1_001110011101;
      patterns[26428] = 29'b0_110011100111_100_1_011001110011;
      patterns[26429] = 29'b0_110011100111_101_1_101100111001;
      patterns[26430] = 29'b0_110011100111_110_0_110011100111;
      patterns[26431] = 29'b0_110011100111_111_0_110011100111;
      patterns[26432] = 29'b0_110011101000_000_0_110011101000;
      patterns[26433] = 29'b0_110011101000_001_0_101000110011;
      patterns[26434] = 29'b0_110011101000_010_1_100111010000;
      patterns[26435] = 29'b0_110011101000_011_1_001110100001;
      patterns[26436] = 29'b0_110011101000_100_0_011001110100;
      patterns[26437] = 29'b0_110011101000_101_0_001100111010;
      patterns[26438] = 29'b0_110011101000_110_0_110011101000;
      patterns[26439] = 29'b0_110011101000_111_0_110011101000;
      patterns[26440] = 29'b0_110011101001_000_0_110011101001;
      patterns[26441] = 29'b0_110011101001_001_0_101001110011;
      patterns[26442] = 29'b0_110011101001_010_1_100111010010;
      patterns[26443] = 29'b0_110011101001_011_1_001110100101;
      patterns[26444] = 29'b0_110011101001_100_1_011001110100;
      patterns[26445] = 29'b0_110011101001_101_0_101100111010;
      patterns[26446] = 29'b0_110011101001_110_0_110011101001;
      patterns[26447] = 29'b0_110011101001_111_0_110011101001;
      patterns[26448] = 29'b0_110011101010_000_0_110011101010;
      patterns[26449] = 29'b0_110011101010_001_0_101010110011;
      patterns[26450] = 29'b0_110011101010_010_1_100111010100;
      patterns[26451] = 29'b0_110011101010_011_1_001110101001;
      patterns[26452] = 29'b0_110011101010_100_0_011001110101;
      patterns[26453] = 29'b0_110011101010_101_1_001100111010;
      patterns[26454] = 29'b0_110011101010_110_0_110011101010;
      patterns[26455] = 29'b0_110011101010_111_0_110011101010;
      patterns[26456] = 29'b0_110011101011_000_0_110011101011;
      patterns[26457] = 29'b0_110011101011_001_0_101011110011;
      patterns[26458] = 29'b0_110011101011_010_1_100111010110;
      patterns[26459] = 29'b0_110011101011_011_1_001110101101;
      patterns[26460] = 29'b0_110011101011_100_1_011001110101;
      patterns[26461] = 29'b0_110011101011_101_1_101100111010;
      patterns[26462] = 29'b0_110011101011_110_0_110011101011;
      patterns[26463] = 29'b0_110011101011_111_0_110011101011;
      patterns[26464] = 29'b0_110011101100_000_0_110011101100;
      patterns[26465] = 29'b0_110011101100_001_0_101100110011;
      patterns[26466] = 29'b0_110011101100_010_1_100111011000;
      patterns[26467] = 29'b0_110011101100_011_1_001110110001;
      patterns[26468] = 29'b0_110011101100_100_0_011001110110;
      patterns[26469] = 29'b0_110011101100_101_0_001100111011;
      patterns[26470] = 29'b0_110011101100_110_0_110011101100;
      patterns[26471] = 29'b0_110011101100_111_0_110011101100;
      patterns[26472] = 29'b0_110011101101_000_0_110011101101;
      patterns[26473] = 29'b0_110011101101_001_0_101101110011;
      patterns[26474] = 29'b0_110011101101_010_1_100111011010;
      patterns[26475] = 29'b0_110011101101_011_1_001110110101;
      patterns[26476] = 29'b0_110011101101_100_1_011001110110;
      patterns[26477] = 29'b0_110011101101_101_0_101100111011;
      patterns[26478] = 29'b0_110011101101_110_0_110011101101;
      patterns[26479] = 29'b0_110011101101_111_0_110011101101;
      patterns[26480] = 29'b0_110011101110_000_0_110011101110;
      patterns[26481] = 29'b0_110011101110_001_0_101110110011;
      patterns[26482] = 29'b0_110011101110_010_1_100111011100;
      patterns[26483] = 29'b0_110011101110_011_1_001110111001;
      patterns[26484] = 29'b0_110011101110_100_0_011001110111;
      patterns[26485] = 29'b0_110011101110_101_1_001100111011;
      patterns[26486] = 29'b0_110011101110_110_0_110011101110;
      patterns[26487] = 29'b0_110011101110_111_0_110011101110;
      patterns[26488] = 29'b0_110011101111_000_0_110011101111;
      patterns[26489] = 29'b0_110011101111_001_0_101111110011;
      patterns[26490] = 29'b0_110011101111_010_1_100111011110;
      patterns[26491] = 29'b0_110011101111_011_1_001110111101;
      patterns[26492] = 29'b0_110011101111_100_1_011001110111;
      patterns[26493] = 29'b0_110011101111_101_1_101100111011;
      patterns[26494] = 29'b0_110011101111_110_0_110011101111;
      patterns[26495] = 29'b0_110011101111_111_0_110011101111;
      patterns[26496] = 29'b0_110011110000_000_0_110011110000;
      patterns[26497] = 29'b0_110011110000_001_0_110000110011;
      patterns[26498] = 29'b0_110011110000_010_1_100111100000;
      patterns[26499] = 29'b0_110011110000_011_1_001111000001;
      patterns[26500] = 29'b0_110011110000_100_0_011001111000;
      patterns[26501] = 29'b0_110011110000_101_0_001100111100;
      patterns[26502] = 29'b0_110011110000_110_0_110011110000;
      patterns[26503] = 29'b0_110011110000_111_0_110011110000;
      patterns[26504] = 29'b0_110011110001_000_0_110011110001;
      patterns[26505] = 29'b0_110011110001_001_0_110001110011;
      patterns[26506] = 29'b0_110011110001_010_1_100111100010;
      patterns[26507] = 29'b0_110011110001_011_1_001111000101;
      patterns[26508] = 29'b0_110011110001_100_1_011001111000;
      patterns[26509] = 29'b0_110011110001_101_0_101100111100;
      patterns[26510] = 29'b0_110011110001_110_0_110011110001;
      patterns[26511] = 29'b0_110011110001_111_0_110011110001;
      patterns[26512] = 29'b0_110011110010_000_0_110011110010;
      patterns[26513] = 29'b0_110011110010_001_0_110010110011;
      patterns[26514] = 29'b0_110011110010_010_1_100111100100;
      patterns[26515] = 29'b0_110011110010_011_1_001111001001;
      patterns[26516] = 29'b0_110011110010_100_0_011001111001;
      patterns[26517] = 29'b0_110011110010_101_1_001100111100;
      patterns[26518] = 29'b0_110011110010_110_0_110011110010;
      patterns[26519] = 29'b0_110011110010_111_0_110011110010;
      patterns[26520] = 29'b0_110011110011_000_0_110011110011;
      patterns[26521] = 29'b0_110011110011_001_0_110011110011;
      patterns[26522] = 29'b0_110011110011_010_1_100111100110;
      patterns[26523] = 29'b0_110011110011_011_1_001111001101;
      patterns[26524] = 29'b0_110011110011_100_1_011001111001;
      patterns[26525] = 29'b0_110011110011_101_1_101100111100;
      patterns[26526] = 29'b0_110011110011_110_0_110011110011;
      patterns[26527] = 29'b0_110011110011_111_0_110011110011;
      patterns[26528] = 29'b0_110011110100_000_0_110011110100;
      patterns[26529] = 29'b0_110011110100_001_0_110100110011;
      patterns[26530] = 29'b0_110011110100_010_1_100111101000;
      patterns[26531] = 29'b0_110011110100_011_1_001111010001;
      patterns[26532] = 29'b0_110011110100_100_0_011001111010;
      patterns[26533] = 29'b0_110011110100_101_0_001100111101;
      patterns[26534] = 29'b0_110011110100_110_0_110011110100;
      patterns[26535] = 29'b0_110011110100_111_0_110011110100;
      patterns[26536] = 29'b0_110011110101_000_0_110011110101;
      patterns[26537] = 29'b0_110011110101_001_0_110101110011;
      patterns[26538] = 29'b0_110011110101_010_1_100111101010;
      patterns[26539] = 29'b0_110011110101_011_1_001111010101;
      patterns[26540] = 29'b0_110011110101_100_1_011001111010;
      patterns[26541] = 29'b0_110011110101_101_0_101100111101;
      patterns[26542] = 29'b0_110011110101_110_0_110011110101;
      patterns[26543] = 29'b0_110011110101_111_0_110011110101;
      patterns[26544] = 29'b0_110011110110_000_0_110011110110;
      patterns[26545] = 29'b0_110011110110_001_0_110110110011;
      patterns[26546] = 29'b0_110011110110_010_1_100111101100;
      patterns[26547] = 29'b0_110011110110_011_1_001111011001;
      patterns[26548] = 29'b0_110011110110_100_0_011001111011;
      patterns[26549] = 29'b0_110011110110_101_1_001100111101;
      patterns[26550] = 29'b0_110011110110_110_0_110011110110;
      patterns[26551] = 29'b0_110011110110_111_0_110011110110;
      patterns[26552] = 29'b0_110011110111_000_0_110011110111;
      patterns[26553] = 29'b0_110011110111_001_0_110111110011;
      patterns[26554] = 29'b0_110011110111_010_1_100111101110;
      patterns[26555] = 29'b0_110011110111_011_1_001111011101;
      patterns[26556] = 29'b0_110011110111_100_1_011001111011;
      patterns[26557] = 29'b0_110011110111_101_1_101100111101;
      patterns[26558] = 29'b0_110011110111_110_0_110011110111;
      patterns[26559] = 29'b0_110011110111_111_0_110011110111;
      patterns[26560] = 29'b0_110011111000_000_0_110011111000;
      patterns[26561] = 29'b0_110011111000_001_0_111000110011;
      patterns[26562] = 29'b0_110011111000_010_1_100111110000;
      patterns[26563] = 29'b0_110011111000_011_1_001111100001;
      patterns[26564] = 29'b0_110011111000_100_0_011001111100;
      patterns[26565] = 29'b0_110011111000_101_0_001100111110;
      patterns[26566] = 29'b0_110011111000_110_0_110011111000;
      patterns[26567] = 29'b0_110011111000_111_0_110011111000;
      patterns[26568] = 29'b0_110011111001_000_0_110011111001;
      patterns[26569] = 29'b0_110011111001_001_0_111001110011;
      patterns[26570] = 29'b0_110011111001_010_1_100111110010;
      patterns[26571] = 29'b0_110011111001_011_1_001111100101;
      patterns[26572] = 29'b0_110011111001_100_1_011001111100;
      patterns[26573] = 29'b0_110011111001_101_0_101100111110;
      patterns[26574] = 29'b0_110011111001_110_0_110011111001;
      patterns[26575] = 29'b0_110011111001_111_0_110011111001;
      patterns[26576] = 29'b0_110011111010_000_0_110011111010;
      patterns[26577] = 29'b0_110011111010_001_0_111010110011;
      patterns[26578] = 29'b0_110011111010_010_1_100111110100;
      patterns[26579] = 29'b0_110011111010_011_1_001111101001;
      patterns[26580] = 29'b0_110011111010_100_0_011001111101;
      patterns[26581] = 29'b0_110011111010_101_1_001100111110;
      patterns[26582] = 29'b0_110011111010_110_0_110011111010;
      patterns[26583] = 29'b0_110011111010_111_0_110011111010;
      patterns[26584] = 29'b0_110011111011_000_0_110011111011;
      patterns[26585] = 29'b0_110011111011_001_0_111011110011;
      patterns[26586] = 29'b0_110011111011_010_1_100111110110;
      patterns[26587] = 29'b0_110011111011_011_1_001111101101;
      patterns[26588] = 29'b0_110011111011_100_1_011001111101;
      patterns[26589] = 29'b0_110011111011_101_1_101100111110;
      patterns[26590] = 29'b0_110011111011_110_0_110011111011;
      patterns[26591] = 29'b0_110011111011_111_0_110011111011;
      patterns[26592] = 29'b0_110011111100_000_0_110011111100;
      patterns[26593] = 29'b0_110011111100_001_0_111100110011;
      patterns[26594] = 29'b0_110011111100_010_1_100111111000;
      patterns[26595] = 29'b0_110011111100_011_1_001111110001;
      patterns[26596] = 29'b0_110011111100_100_0_011001111110;
      patterns[26597] = 29'b0_110011111100_101_0_001100111111;
      patterns[26598] = 29'b0_110011111100_110_0_110011111100;
      patterns[26599] = 29'b0_110011111100_111_0_110011111100;
      patterns[26600] = 29'b0_110011111101_000_0_110011111101;
      patterns[26601] = 29'b0_110011111101_001_0_111101110011;
      patterns[26602] = 29'b0_110011111101_010_1_100111111010;
      patterns[26603] = 29'b0_110011111101_011_1_001111110101;
      patterns[26604] = 29'b0_110011111101_100_1_011001111110;
      patterns[26605] = 29'b0_110011111101_101_0_101100111111;
      patterns[26606] = 29'b0_110011111101_110_0_110011111101;
      patterns[26607] = 29'b0_110011111101_111_0_110011111101;
      patterns[26608] = 29'b0_110011111110_000_0_110011111110;
      patterns[26609] = 29'b0_110011111110_001_0_111110110011;
      patterns[26610] = 29'b0_110011111110_010_1_100111111100;
      patterns[26611] = 29'b0_110011111110_011_1_001111111001;
      patterns[26612] = 29'b0_110011111110_100_0_011001111111;
      patterns[26613] = 29'b0_110011111110_101_1_001100111111;
      patterns[26614] = 29'b0_110011111110_110_0_110011111110;
      patterns[26615] = 29'b0_110011111110_111_0_110011111110;
      patterns[26616] = 29'b0_110011111111_000_0_110011111111;
      patterns[26617] = 29'b0_110011111111_001_0_111111110011;
      patterns[26618] = 29'b0_110011111111_010_1_100111111110;
      patterns[26619] = 29'b0_110011111111_011_1_001111111101;
      patterns[26620] = 29'b0_110011111111_100_1_011001111111;
      patterns[26621] = 29'b0_110011111111_101_1_101100111111;
      patterns[26622] = 29'b0_110011111111_110_0_110011111111;
      patterns[26623] = 29'b0_110011111111_111_0_110011111111;
      patterns[26624] = 29'b0_110100000000_000_0_110100000000;
      patterns[26625] = 29'b0_110100000000_001_0_000000110100;
      patterns[26626] = 29'b0_110100000000_010_1_101000000000;
      patterns[26627] = 29'b0_110100000000_011_1_010000000001;
      patterns[26628] = 29'b0_110100000000_100_0_011010000000;
      patterns[26629] = 29'b0_110100000000_101_0_001101000000;
      patterns[26630] = 29'b0_110100000000_110_0_110100000000;
      patterns[26631] = 29'b0_110100000000_111_0_110100000000;
      patterns[26632] = 29'b0_110100000001_000_0_110100000001;
      patterns[26633] = 29'b0_110100000001_001_0_000001110100;
      patterns[26634] = 29'b0_110100000001_010_1_101000000010;
      patterns[26635] = 29'b0_110100000001_011_1_010000000101;
      patterns[26636] = 29'b0_110100000001_100_1_011010000000;
      patterns[26637] = 29'b0_110100000001_101_0_101101000000;
      patterns[26638] = 29'b0_110100000001_110_0_110100000001;
      patterns[26639] = 29'b0_110100000001_111_0_110100000001;
      patterns[26640] = 29'b0_110100000010_000_0_110100000010;
      patterns[26641] = 29'b0_110100000010_001_0_000010110100;
      patterns[26642] = 29'b0_110100000010_010_1_101000000100;
      patterns[26643] = 29'b0_110100000010_011_1_010000001001;
      patterns[26644] = 29'b0_110100000010_100_0_011010000001;
      patterns[26645] = 29'b0_110100000010_101_1_001101000000;
      patterns[26646] = 29'b0_110100000010_110_0_110100000010;
      patterns[26647] = 29'b0_110100000010_111_0_110100000010;
      patterns[26648] = 29'b0_110100000011_000_0_110100000011;
      patterns[26649] = 29'b0_110100000011_001_0_000011110100;
      patterns[26650] = 29'b0_110100000011_010_1_101000000110;
      patterns[26651] = 29'b0_110100000011_011_1_010000001101;
      patterns[26652] = 29'b0_110100000011_100_1_011010000001;
      patterns[26653] = 29'b0_110100000011_101_1_101101000000;
      patterns[26654] = 29'b0_110100000011_110_0_110100000011;
      patterns[26655] = 29'b0_110100000011_111_0_110100000011;
      patterns[26656] = 29'b0_110100000100_000_0_110100000100;
      patterns[26657] = 29'b0_110100000100_001_0_000100110100;
      patterns[26658] = 29'b0_110100000100_010_1_101000001000;
      patterns[26659] = 29'b0_110100000100_011_1_010000010001;
      patterns[26660] = 29'b0_110100000100_100_0_011010000010;
      patterns[26661] = 29'b0_110100000100_101_0_001101000001;
      patterns[26662] = 29'b0_110100000100_110_0_110100000100;
      patterns[26663] = 29'b0_110100000100_111_0_110100000100;
      patterns[26664] = 29'b0_110100000101_000_0_110100000101;
      patterns[26665] = 29'b0_110100000101_001_0_000101110100;
      patterns[26666] = 29'b0_110100000101_010_1_101000001010;
      patterns[26667] = 29'b0_110100000101_011_1_010000010101;
      patterns[26668] = 29'b0_110100000101_100_1_011010000010;
      patterns[26669] = 29'b0_110100000101_101_0_101101000001;
      patterns[26670] = 29'b0_110100000101_110_0_110100000101;
      patterns[26671] = 29'b0_110100000101_111_0_110100000101;
      patterns[26672] = 29'b0_110100000110_000_0_110100000110;
      patterns[26673] = 29'b0_110100000110_001_0_000110110100;
      patterns[26674] = 29'b0_110100000110_010_1_101000001100;
      patterns[26675] = 29'b0_110100000110_011_1_010000011001;
      patterns[26676] = 29'b0_110100000110_100_0_011010000011;
      patterns[26677] = 29'b0_110100000110_101_1_001101000001;
      patterns[26678] = 29'b0_110100000110_110_0_110100000110;
      patterns[26679] = 29'b0_110100000110_111_0_110100000110;
      patterns[26680] = 29'b0_110100000111_000_0_110100000111;
      patterns[26681] = 29'b0_110100000111_001_0_000111110100;
      patterns[26682] = 29'b0_110100000111_010_1_101000001110;
      patterns[26683] = 29'b0_110100000111_011_1_010000011101;
      patterns[26684] = 29'b0_110100000111_100_1_011010000011;
      patterns[26685] = 29'b0_110100000111_101_1_101101000001;
      patterns[26686] = 29'b0_110100000111_110_0_110100000111;
      patterns[26687] = 29'b0_110100000111_111_0_110100000111;
      patterns[26688] = 29'b0_110100001000_000_0_110100001000;
      patterns[26689] = 29'b0_110100001000_001_0_001000110100;
      patterns[26690] = 29'b0_110100001000_010_1_101000010000;
      patterns[26691] = 29'b0_110100001000_011_1_010000100001;
      patterns[26692] = 29'b0_110100001000_100_0_011010000100;
      patterns[26693] = 29'b0_110100001000_101_0_001101000010;
      patterns[26694] = 29'b0_110100001000_110_0_110100001000;
      patterns[26695] = 29'b0_110100001000_111_0_110100001000;
      patterns[26696] = 29'b0_110100001001_000_0_110100001001;
      patterns[26697] = 29'b0_110100001001_001_0_001001110100;
      patterns[26698] = 29'b0_110100001001_010_1_101000010010;
      patterns[26699] = 29'b0_110100001001_011_1_010000100101;
      patterns[26700] = 29'b0_110100001001_100_1_011010000100;
      patterns[26701] = 29'b0_110100001001_101_0_101101000010;
      patterns[26702] = 29'b0_110100001001_110_0_110100001001;
      patterns[26703] = 29'b0_110100001001_111_0_110100001001;
      patterns[26704] = 29'b0_110100001010_000_0_110100001010;
      patterns[26705] = 29'b0_110100001010_001_0_001010110100;
      patterns[26706] = 29'b0_110100001010_010_1_101000010100;
      patterns[26707] = 29'b0_110100001010_011_1_010000101001;
      patterns[26708] = 29'b0_110100001010_100_0_011010000101;
      patterns[26709] = 29'b0_110100001010_101_1_001101000010;
      patterns[26710] = 29'b0_110100001010_110_0_110100001010;
      patterns[26711] = 29'b0_110100001010_111_0_110100001010;
      patterns[26712] = 29'b0_110100001011_000_0_110100001011;
      patterns[26713] = 29'b0_110100001011_001_0_001011110100;
      patterns[26714] = 29'b0_110100001011_010_1_101000010110;
      patterns[26715] = 29'b0_110100001011_011_1_010000101101;
      patterns[26716] = 29'b0_110100001011_100_1_011010000101;
      patterns[26717] = 29'b0_110100001011_101_1_101101000010;
      patterns[26718] = 29'b0_110100001011_110_0_110100001011;
      patterns[26719] = 29'b0_110100001011_111_0_110100001011;
      patterns[26720] = 29'b0_110100001100_000_0_110100001100;
      patterns[26721] = 29'b0_110100001100_001_0_001100110100;
      patterns[26722] = 29'b0_110100001100_010_1_101000011000;
      patterns[26723] = 29'b0_110100001100_011_1_010000110001;
      patterns[26724] = 29'b0_110100001100_100_0_011010000110;
      patterns[26725] = 29'b0_110100001100_101_0_001101000011;
      patterns[26726] = 29'b0_110100001100_110_0_110100001100;
      patterns[26727] = 29'b0_110100001100_111_0_110100001100;
      patterns[26728] = 29'b0_110100001101_000_0_110100001101;
      patterns[26729] = 29'b0_110100001101_001_0_001101110100;
      patterns[26730] = 29'b0_110100001101_010_1_101000011010;
      patterns[26731] = 29'b0_110100001101_011_1_010000110101;
      patterns[26732] = 29'b0_110100001101_100_1_011010000110;
      patterns[26733] = 29'b0_110100001101_101_0_101101000011;
      patterns[26734] = 29'b0_110100001101_110_0_110100001101;
      patterns[26735] = 29'b0_110100001101_111_0_110100001101;
      patterns[26736] = 29'b0_110100001110_000_0_110100001110;
      patterns[26737] = 29'b0_110100001110_001_0_001110110100;
      patterns[26738] = 29'b0_110100001110_010_1_101000011100;
      patterns[26739] = 29'b0_110100001110_011_1_010000111001;
      patterns[26740] = 29'b0_110100001110_100_0_011010000111;
      patterns[26741] = 29'b0_110100001110_101_1_001101000011;
      patterns[26742] = 29'b0_110100001110_110_0_110100001110;
      patterns[26743] = 29'b0_110100001110_111_0_110100001110;
      patterns[26744] = 29'b0_110100001111_000_0_110100001111;
      patterns[26745] = 29'b0_110100001111_001_0_001111110100;
      patterns[26746] = 29'b0_110100001111_010_1_101000011110;
      patterns[26747] = 29'b0_110100001111_011_1_010000111101;
      patterns[26748] = 29'b0_110100001111_100_1_011010000111;
      patterns[26749] = 29'b0_110100001111_101_1_101101000011;
      patterns[26750] = 29'b0_110100001111_110_0_110100001111;
      patterns[26751] = 29'b0_110100001111_111_0_110100001111;
      patterns[26752] = 29'b0_110100010000_000_0_110100010000;
      patterns[26753] = 29'b0_110100010000_001_0_010000110100;
      patterns[26754] = 29'b0_110100010000_010_1_101000100000;
      patterns[26755] = 29'b0_110100010000_011_1_010001000001;
      patterns[26756] = 29'b0_110100010000_100_0_011010001000;
      patterns[26757] = 29'b0_110100010000_101_0_001101000100;
      patterns[26758] = 29'b0_110100010000_110_0_110100010000;
      patterns[26759] = 29'b0_110100010000_111_0_110100010000;
      patterns[26760] = 29'b0_110100010001_000_0_110100010001;
      patterns[26761] = 29'b0_110100010001_001_0_010001110100;
      patterns[26762] = 29'b0_110100010001_010_1_101000100010;
      patterns[26763] = 29'b0_110100010001_011_1_010001000101;
      patterns[26764] = 29'b0_110100010001_100_1_011010001000;
      patterns[26765] = 29'b0_110100010001_101_0_101101000100;
      patterns[26766] = 29'b0_110100010001_110_0_110100010001;
      patterns[26767] = 29'b0_110100010001_111_0_110100010001;
      patterns[26768] = 29'b0_110100010010_000_0_110100010010;
      patterns[26769] = 29'b0_110100010010_001_0_010010110100;
      patterns[26770] = 29'b0_110100010010_010_1_101000100100;
      patterns[26771] = 29'b0_110100010010_011_1_010001001001;
      patterns[26772] = 29'b0_110100010010_100_0_011010001001;
      patterns[26773] = 29'b0_110100010010_101_1_001101000100;
      patterns[26774] = 29'b0_110100010010_110_0_110100010010;
      patterns[26775] = 29'b0_110100010010_111_0_110100010010;
      patterns[26776] = 29'b0_110100010011_000_0_110100010011;
      patterns[26777] = 29'b0_110100010011_001_0_010011110100;
      patterns[26778] = 29'b0_110100010011_010_1_101000100110;
      patterns[26779] = 29'b0_110100010011_011_1_010001001101;
      patterns[26780] = 29'b0_110100010011_100_1_011010001001;
      patterns[26781] = 29'b0_110100010011_101_1_101101000100;
      patterns[26782] = 29'b0_110100010011_110_0_110100010011;
      patterns[26783] = 29'b0_110100010011_111_0_110100010011;
      patterns[26784] = 29'b0_110100010100_000_0_110100010100;
      patterns[26785] = 29'b0_110100010100_001_0_010100110100;
      patterns[26786] = 29'b0_110100010100_010_1_101000101000;
      patterns[26787] = 29'b0_110100010100_011_1_010001010001;
      patterns[26788] = 29'b0_110100010100_100_0_011010001010;
      patterns[26789] = 29'b0_110100010100_101_0_001101000101;
      patterns[26790] = 29'b0_110100010100_110_0_110100010100;
      patterns[26791] = 29'b0_110100010100_111_0_110100010100;
      patterns[26792] = 29'b0_110100010101_000_0_110100010101;
      patterns[26793] = 29'b0_110100010101_001_0_010101110100;
      patterns[26794] = 29'b0_110100010101_010_1_101000101010;
      patterns[26795] = 29'b0_110100010101_011_1_010001010101;
      patterns[26796] = 29'b0_110100010101_100_1_011010001010;
      patterns[26797] = 29'b0_110100010101_101_0_101101000101;
      patterns[26798] = 29'b0_110100010101_110_0_110100010101;
      patterns[26799] = 29'b0_110100010101_111_0_110100010101;
      patterns[26800] = 29'b0_110100010110_000_0_110100010110;
      patterns[26801] = 29'b0_110100010110_001_0_010110110100;
      patterns[26802] = 29'b0_110100010110_010_1_101000101100;
      patterns[26803] = 29'b0_110100010110_011_1_010001011001;
      patterns[26804] = 29'b0_110100010110_100_0_011010001011;
      patterns[26805] = 29'b0_110100010110_101_1_001101000101;
      patterns[26806] = 29'b0_110100010110_110_0_110100010110;
      patterns[26807] = 29'b0_110100010110_111_0_110100010110;
      patterns[26808] = 29'b0_110100010111_000_0_110100010111;
      patterns[26809] = 29'b0_110100010111_001_0_010111110100;
      patterns[26810] = 29'b0_110100010111_010_1_101000101110;
      patterns[26811] = 29'b0_110100010111_011_1_010001011101;
      patterns[26812] = 29'b0_110100010111_100_1_011010001011;
      patterns[26813] = 29'b0_110100010111_101_1_101101000101;
      patterns[26814] = 29'b0_110100010111_110_0_110100010111;
      patterns[26815] = 29'b0_110100010111_111_0_110100010111;
      patterns[26816] = 29'b0_110100011000_000_0_110100011000;
      patterns[26817] = 29'b0_110100011000_001_0_011000110100;
      patterns[26818] = 29'b0_110100011000_010_1_101000110000;
      patterns[26819] = 29'b0_110100011000_011_1_010001100001;
      patterns[26820] = 29'b0_110100011000_100_0_011010001100;
      patterns[26821] = 29'b0_110100011000_101_0_001101000110;
      patterns[26822] = 29'b0_110100011000_110_0_110100011000;
      patterns[26823] = 29'b0_110100011000_111_0_110100011000;
      patterns[26824] = 29'b0_110100011001_000_0_110100011001;
      patterns[26825] = 29'b0_110100011001_001_0_011001110100;
      patterns[26826] = 29'b0_110100011001_010_1_101000110010;
      patterns[26827] = 29'b0_110100011001_011_1_010001100101;
      patterns[26828] = 29'b0_110100011001_100_1_011010001100;
      patterns[26829] = 29'b0_110100011001_101_0_101101000110;
      patterns[26830] = 29'b0_110100011001_110_0_110100011001;
      patterns[26831] = 29'b0_110100011001_111_0_110100011001;
      patterns[26832] = 29'b0_110100011010_000_0_110100011010;
      patterns[26833] = 29'b0_110100011010_001_0_011010110100;
      patterns[26834] = 29'b0_110100011010_010_1_101000110100;
      patterns[26835] = 29'b0_110100011010_011_1_010001101001;
      patterns[26836] = 29'b0_110100011010_100_0_011010001101;
      patterns[26837] = 29'b0_110100011010_101_1_001101000110;
      patterns[26838] = 29'b0_110100011010_110_0_110100011010;
      patterns[26839] = 29'b0_110100011010_111_0_110100011010;
      patterns[26840] = 29'b0_110100011011_000_0_110100011011;
      patterns[26841] = 29'b0_110100011011_001_0_011011110100;
      patterns[26842] = 29'b0_110100011011_010_1_101000110110;
      patterns[26843] = 29'b0_110100011011_011_1_010001101101;
      patterns[26844] = 29'b0_110100011011_100_1_011010001101;
      patterns[26845] = 29'b0_110100011011_101_1_101101000110;
      patterns[26846] = 29'b0_110100011011_110_0_110100011011;
      patterns[26847] = 29'b0_110100011011_111_0_110100011011;
      patterns[26848] = 29'b0_110100011100_000_0_110100011100;
      patterns[26849] = 29'b0_110100011100_001_0_011100110100;
      patterns[26850] = 29'b0_110100011100_010_1_101000111000;
      patterns[26851] = 29'b0_110100011100_011_1_010001110001;
      patterns[26852] = 29'b0_110100011100_100_0_011010001110;
      patterns[26853] = 29'b0_110100011100_101_0_001101000111;
      patterns[26854] = 29'b0_110100011100_110_0_110100011100;
      patterns[26855] = 29'b0_110100011100_111_0_110100011100;
      patterns[26856] = 29'b0_110100011101_000_0_110100011101;
      patterns[26857] = 29'b0_110100011101_001_0_011101110100;
      patterns[26858] = 29'b0_110100011101_010_1_101000111010;
      patterns[26859] = 29'b0_110100011101_011_1_010001110101;
      patterns[26860] = 29'b0_110100011101_100_1_011010001110;
      patterns[26861] = 29'b0_110100011101_101_0_101101000111;
      patterns[26862] = 29'b0_110100011101_110_0_110100011101;
      patterns[26863] = 29'b0_110100011101_111_0_110100011101;
      patterns[26864] = 29'b0_110100011110_000_0_110100011110;
      patterns[26865] = 29'b0_110100011110_001_0_011110110100;
      patterns[26866] = 29'b0_110100011110_010_1_101000111100;
      patterns[26867] = 29'b0_110100011110_011_1_010001111001;
      patterns[26868] = 29'b0_110100011110_100_0_011010001111;
      patterns[26869] = 29'b0_110100011110_101_1_001101000111;
      patterns[26870] = 29'b0_110100011110_110_0_110100011110;
      patterns[26871] = 29'b0_110100011110_111_0_110100011110;
      patterns[26872] = 29'b0_110100011111_000_0_110100011111;
      patterns[26873] = 29'b0_110100011111_001_0_011111110100;
      patterns[26874] = 29'b0_110100011111_010_1_101000111110;
      patterns[26875] = 29'b0_110100011111_011_1_010001111101;
      patterns[26876] = 29'b0_110100011111_100_1_011010001111;
      patterns[26877] = 29'b0_110100011111_101_1_101101000111;
      patterns[26878] = 29'b0_110100011111_110_0_110100011111;
      patterns[26879] = 29'b0_110100011111_111_0_110100011111;
      patterns[26880] = 29'b0_110100100000_000_0_110100100000;
      patterns[26881] = 29'b0_110100100000_001_0_100000110100;
      patterns[26882] = 29'b0_110100100000_010_1_101001000000;
      patterns[26883] = 29'b0_110100100000_011_1_010010000001;
      patterns[26884] = 29'b0_110100100000_100_0_011010010000;
      patterns[26885] = 29'b0_110100100000_101_0_001101001000;
      patterns[26886] = 29'b0_110100100000_110_0_110100100000;
      patterns[26887] = 29'b0_110100100000_111_0_110100100000;
      patterns[26888] = 29'b0_110100100001_000_0_110100100001;
      patterns[26889] = 29'b0_110100100001_001_0_100001110100;
      patterns[26890] = 29'b0_110100100001_010_1_101001000010;
      patterns[26891] = 29'b0_110100100001_011_1_010010000101;
      patterns[26892] = 29'b0_110100100001_100_1_011010010000;
      patterns[26893] = 29'b0_110100100001_101_0_101101001000;
      patterns[26894] = 29'b0_110100100001_110_0_110100100001;
      patterns[26895] = 29'b0_110100100001_111_0_110100100001;
      patterns[26896] = 29'b0_110100100010_000_0_110100100010;
      patterns[26897] = 29'b0_110100100010_001_0_100010110100;
      patterns[26898] = 29'b0_110100100010_010_1_101001000100;
      patterns[26899] = 29'b0_110100100010_011_1_010010001001;
      patterns[26900] = 29'b0_110100100010_100_0_011010010001;
      patterns[26901] = 29'b0_110100100010_101_1_001101001000;
      patterns[26902] = 29'b0_110100100010_110_0_110100100010;
      patterns[26903] = 29'b0_110100100010_111_0_110100100010;
      patterns[26904] = 29'b0_110100100011_000_0_110100100011;
      patterns[26905] = 29'b0_110100100011_001_0_100011110100;
      patterns[26906] = 29'b0_110100100011_010_1_101001000110;
      patterns[26907] = 29'b0_110100100011_011_1_010010001101;
      patterns[26908] = 29'b0_110100100011_100_1_011010010001;
      patterns[26909] = 29'b0_110100100011_101_1_101101001000;
      patterns[26910] = 29'b0_110100100011_110_0_110100100011;
      patterns[26911] = 29'b0_110100100011_111_0_110100100011;
      patterns[26912] = 29'b0_110100100100_000_0_110100100100;
      patterns[26913] = 29'b0_110100100100_001_0_100100110100;
      patterns[26914] = 29'b0_110100100100_010_1_101001001000;
      patterns[26915] = 29'b0_110100100100_011_1_010010010001;
      patterns[26916] = 29'b0_110100100100_100_0_011010010010;
      patterns[26917] = 29'b0_110100100100_101_0_001101001001;
      patterns[26918] = 29'b0_110100100100_110_0_110100100100;
      patterns[26919] = 29'b0_110100100100_111_0_110100100100;
      patterns[26920] = 29'b0_110100100101_000_0_110100100101;
      patterns[26921] = 29'b0_110100100101_001_0_100101110100;
      patterns[26922] = 29'b0_110100100101_010_1_101001001010;
      patterns[26923] = 29'b0_110100100101_011_1_010010010101;
      patterns[26924] = 29'b0_110100100101_100_1_011010010010;
      patterns[26925] = 29'b0_110100100101_101_0_101101001001;
      patterns[26926] = 29'b0_110100100101_110_0_110100100101;
      patterns[26927] = 29'b0_110100100101_111_0_110100100101;
      patterns[26928] = 29'b0_110100100110_000_0_110100100110;
      patterns[26929] = 29'b0_110100100110_001_0_100110110100;
      patterns[26930] = 29'b0_110100100110_010_1_101001001100;
      patterns[26931] = 29'b0_110100100110_011_1_010010011001;
      patterns[26932] = 29'b0_110100100110_100_0_011010010011;
      patterns[26933] = 29'b0_110100100110_101_1_001101001001;
      patterns[26934] = 29'b0_110100100110_110_0_110100100110;
      patterns[26935] = 29'b0_110100100110_111_0_110100100110;
      patterns[26936] = 29'b0_110100100111_000_0_110100100111;
      patterns[26937] = 29'b0_110100100111_001_0_100111110100;
      patterns[26938] = 29'b0_110100100111_010_1_101001001110;
      patterns[26939] = 29'b0_110100100111_011_1_010010011101;
      patterns[26940] = 29'b0_110100100111_100_1_011010010011;
      patterns[26941] = 29'b0_110100100111_101_1_101101001001;
      patterns[26942] = 29'b0_110100100111_110_0_110100100111;
      patterns[26943] = 29'b0_110100100111_111_0_110100100111;
      patterns[26944] = 29'b0_110100101000_000_0_110100101000;
      patterns[26945] = 29'b0_110100101000_001_0_101000110100;
      patterns[26946] = 29'b0_110100101000_010_1_101001010000;
      patterns[26947] = 29'b0_110100101000_011_1_010010100001;
      patterns[26948] = 29'b0_110100101000_100_0_011010010100;
      patterns[26949] = 29'b0_110100101000_101_0_001101001010;
      patterns[26950] = 29'b0_110100101000_110_0_110100101000;
      patterns[26951] = 29'b0_110100101000_111_0_110100101000;
      patterns[26952] = 29'b0_110100101001_000_0_110100101001;
      patterns[26953] = 29'b0_110100101001_001_0_101001110100;
      patterns[26954] = 29'b0_110100101001_010_1_101001010010;
      patterns[26955] = 29'b0_110100101001_011_1_010010100101;
      patterns[26956] = 29'b0_110100101001_100_1_011010010100;
      patterns[26957] = 29'b0_110100101001_101_0_101101001010;
      patterns[26958] = 29'b0_110100101001_110_0_110100101001;
      patterns[26959] = 29'b0_110100101001_111_0_110100101001;
      patterns[26960] = 29'b0_110100101010_000_0_110100101010;
      patterns[26961] = 29'b0_110100101010_001_0_101010110100;
      patterns[26962] = 29'b0_110100101010_010_1_101001010100;
      patterns[26963] = 29'b0_110100101010_011_1_010010101001;
      patterns[26964] = 29'b0_110100101010_100_0_011010010101;
      patterns[26965] = 29'b0_110100101010_101_1_001101001010;
      patterns[26966] = 29'b0_110100101010_110_0_110100101010;
      patterns[26967] = 29'b0_110100101010_111_0_110100101010;
      patterns[26968] = 29'b0_110100101011_000_0_110100101011;
      patterns[26969] = 29'b0_110100101011_001_0_101011110100;
      patterns[26970] = 29'b0_110100101011_010_1_101001010110;
      patterns[26971] = 29'b0_110100101011_011_1_010010101101;
      patterns[26972] = 29'b0_110100101011_100_1_011010010101;
      patterns[26973] = 29'b0_110100101011_101_1_101101001010;
      patterns[26974] = 29'b0_110100101011_110_0_110100101011;
      patterns[26975] = 29'b0_110100101011_111_0_110100101011;
      patterns[26976] = 29'b0_110100101100_000_0_110100101100;
      patterns[26977] = 29'b0_110100101100_001_0_101100110100;
      patterns[26978] = 29'b0_110100101100_010_1_101001011000;
      patterns[26979] = 29'b0_110100101100_011_1_010010110001;
      patterns[26980] = 29'b0_110100101100_100_0_011010010110;
      patterns[26981] = 29'b0_110100101100_101_0_001101001011;
      patterns[26982] = 29'b0_110100101100_110_0_110100101100;
      patterns[26983] = 29'b0_110100101100_111_0_110100101100;
      patterns[26984] = 29'b0_110100101101_000_0_110100101101;
      patterns[26985] = 29'b0_110100101101_001_0_101101110100;
      patterns[26986] = 29'b0_110100101101_010_1_101001011010;
      patterns[26987] = 29'b0_110100101101_011_1_010010110101;
      patterns[26988] = 29'b0_110100101101_100_1_011010010110;
      patterns[26989] = 29'b0_110100101101_101_0_101101001011;
      patterns[26990] = 29'b0_110100101101_110_0_110100101101;
      patterns[26991] = 29'b0_110100101101_111_0_110100101101;
      patterns[26992] = 29'b0_110100101110_000_0_110100101110;
      patterns[26993] = 29'b0_110100101110_001_0_101110110100;
      patterns[26994] = 29'b0_110100101110_010_1_101001011100;
      patterns[26995] = 29'b0_110100101110_011_1_010010111001;
      patterns[26996] = 29'b0_110100101110_100_0_011010010111;
      patterns[26997] = 29'b0_110100101110_101_1_001101001011;
      patterns[26998] = 29'b0_110100101110_110_0_110100101110;
      patterns[26999] = 29'b0_110100101110_111_0_110100101110;
      patterns[27000] = 29'b0_110100101111_000_0_110100101111;
      patterns[27001] = 29'b0_110100101111_001_0_101111110100;
      patterns[27002] = 29'b0_110100101111_010_1_101001011110;
      patterns[27003] = 29'b0_110100101111_011_1_010010111101;
      patterns[27004] = 29'b0_110100101111_100_1_011010010111;
      patterns[27005] = 29'b0_110100101111_101_1_101101001011;
      patterns[27006] = 29'b0_110100101111_110_0_110100101111;
      patterns[27007] = 29'b0_110100101111_111_0_110100101111;
      patterns[27008] = 29'b0_110100110000_000_0_110100110000;
      patterns[27009] = 29'b0_110100110000_001_0_110000110100;
      patterns[27010] = 29'b0_110100110000_010_1_101001100000;
      patterns[27011] = 29'b0_110100110000_011_1_010011000001;
      patterns[27012] = 29'b0_110100110000_100_0_011010011000;
      patterns[27013] = 29'b0_110100110000_101_0_001101001100;
      patterns[27014] = 29'b0_110100110000_110_0_110100110000;
      patterns[27015] = 29'b0_110100110000_111_0_110100110000;
      patterns[27016] = 29'b0_110100110001_000_0_110100110001;
      patterns[27017] = 29'b0_110100110001_001_0_110001110100;
      patterns[27018] = 29'b0_110100110001_010_1_101001100010;
      patterns[27019] = 29'b0_110100110001_011_1_010011000101;
      patterns[27020] = 29'b0_110100110001_100_1_011010011000;
      patterns[27021] = 29'b0_110100110001_101_0_101101001100;
      patterns[27022] = 29'b0_110100110001_110_0_110100110001;
      patterns[27023] = 29'b0_110100110001_111_0_110100110001;
      patterns[27024] = 29'b0_110100110010_000_0_110100110010;
      patterns[27025] = 29'b0_110100110010_001_0_110010110100;
      patterns[27026] = 29'b0_110100110010_010_1_101001100100;
      patterns[27027] = 29'b0_110100110010_011_1_010011001001;
      patterns[27028] = 29'b0_110100110010_100_0_011010011001;
      patterns[27029] = 29'b0_110100110010_101_1_001101001100;
      patterns[27030] = 29'b0_110100110010_110_0_110100110010;
      patterns[27031] = 29'b0_110100110010_111_0_110100110010;
      patterns[27032] = 29'b0_110100110011_000_0_110100110011;
      patterns[27033] = 29'b0_110100110011_001_0_110011110100;
      patterns[27034] = 29'b0_110100110011_010_1_101001100110;
      patterns[27035] = 29'b0_110100110011_011_1_010011001101;
      patterns[27036] = 29'b0_110100110011_100_1_011010011001;
      patterns[27037] = 29'b0_110100110011_101_1_101101001100;
      patterns[27038] = 29'b0_110100110011_110_0_110100110011;
      patterns[27039] = 29'b0_110100110011_111_0_110100110011;
      patterns[27040] = 29'b0_110100110100_000_0_110100110100;
      patterns[27041] = 29'b0_110100110100_001_0_110100110100;
      patterns[27042] = 29'b0_110100110100_010_1_101001101000;
      patterns[27043] = 29'b0_110100110100_011_1_010011010001;
      patterns[27044] = 29'b0_110100110100_100_0_011010011010;
      patterns[27045] = 29'b0_110100110100_101_0_001101001101;
      patterns[27046] = 29'b0_110100110100_110_0_110100110100;
      patterns[27047] = 29'b0_110100110100_111_0_110100110100;
      patterns[27048] = 29'b0_110100110101_000_0_110100110101;
      patterns[27049] = 29'b0_110100110101_001_0_110101110100;
      patterns[27050] = 29'b0_110100110101_010_1_101001101010;
      patterns[27051] = 29'b0_110100110101_011_1_010011010101;
      patterns[27052] = 29'b0_110100110101_100_1_011010011010;
      patterns[27053] = 29'b0_110100110101_101_0_101101001101;
      patterns[27054] = 29'b0_110100110101_110_0_110100110101;
      patterns[27055] = 29'b0_110100110101_111_0_110100110101;
      patterns[27056] = 29'b0_110100110110_000_0_110100110110;
      patterns[27057] = 29'b0_110100110110_001_0_110110110100;
      patterns[27058] = 29'b0_110100110110_010_1_101001101100;
      patterns[27059] = 29'b0_110100110110_011_1_010011011001;
      patterns[27060] = 29'b0_110100110110_100_0_011010011011;
      patterns[27061] = 29'b0_110100110110_101_1_001101001101;
      patterns[27062] = 29'b0_110100110110_110_0_110100110110;
      patterns[27063] = 29'b0_110100110110_111_0_110100110110;
      patterns[27064] = 29'b0_110100110111_000_0_110100110111;
      patterns[27065] = 29'b0_110100110111_001_0_110111110100;
      patterns[27066] = 29'b0_110100110111_010_1_101001101110;
      patterns[27067] = 29'b0_110100110111_011_1_010011011101;
      patterns[27068] = 29'b0_110100110111_100_1_011010011011;
      patterns[27069] = 29'b0_110100110111_101_1_101101001101;
      patterns[27070] = 29'b0_110100110111_110_0_110100110111;
      patterns[27071] = 29'b0_110100110111_111_0_110100110111;
      patterns[27072] = 29'b0_110100111000_000_0_110100111000;
      patterns[27073] = 29'b0_110100111000_001_0_111000110100;
      patterns[27074] = 29'b0_110100111000_010_1_101001110000;
      patterns[27075] = 29'b0_110100111000_011_1_010011100001;
      patterns[27076] = 29'b0_110100111000_100_0_011010011100;
      patterns[27077] = 29'b0_110100111000_101_0_001101001110;
      patterns[27078] = 29'b0_110100111000_110_0_110100111000;
      patterns[27079] = 29'b0_110100111000_111_0_110100111000;
      patterns[27080] = 29'b0_110100111001_000_0_110100111001;
      patterns[27081] = 29'b0_110100111001_001_0_111001110100;
      patterns[27082] = 29'b0_110100111001_010_1_101001110010;
      patterns[27083] = 29'b0_110100111001_011_1_010011100101;
      patterns[27084] = 29'b0_110100111001_100_1_011010011100;
      patterns[27085] = 29'b0_110100111001_101_0_101101001110;
      patterns[27086] = 29'b0_110100111001_110_0_110100111001;
      patterns[27087] = 29'b0_110100111001_111_0_110100111001;
      patterns[27088] = 29'b0_110100111010_000_0_110100111010;
      patterns[27089] = 29'b0_110100111010_001_0_111010110100;
      patterns[27090] = 29'b0_110100111010_010_1_101001110100;
      patterns[27091] = 29'b0_110100111010_011_1_010011101001;
      patterns[27092] = 29'b0_110100111010_100_0_011010011101;
      patterns[27093] = 29'b0_110100111010_101_1_001101001110;
      patterns[27094] = 29'b0_110100111010_110_0_110100111010;
      patterns[27095] = 29'b0_110100111010_111_0_110100111010;
      patterns[27096] = 29'b0_110100111011_000_0_110100111011;
      patterns[27097] = 29'b0_110100111011_001_0_111011110100;
      patterns[27098] = 29'b0_110100111011_010_1_101001110110;
      patterns[27099] = 29'b0_110100111011_011_1_010011101101;
      patterns[27100] = 29'b0_110100111011_100_1_011010011101;
      patterns[27101] = 29'b0_110100111011_101_1_101101001110;
      patterns[27102] = 29'b0_110100111011_110_0_110100111011;
      patterns[27103] = 29'b0_110100111011_111_0_110100111011;
      patterns[27104] = 29'b0_110100111100_000_0_110100111100;
      patterns[27105] = 29'b0_110100111100_001_0_111100110100;
      patterns[27106] = 29'b0_110100111100_010_1_101001111000;
      patterns[27107] = 29'b0_110100111100_011_1_010011110001;
      patterns[27108] = 29'b0_110100111100_100_0_011010011110;
      patterns[27109] = 29'b0_110100111100_101_0_001101001111;
      patterns[27110] = 29'b0_110100111100_110_0_110100111100;
      patterns[27111] = 29'b0_110100111100_111_0_110100111100;
      patterns[27112] = 29'b0_110100111101_000_0_110100111101;
      patterns[27113] = 29'b0_110100111101_001_0_111101110100;
      patterns[27114] = 29'b0_110100111101_010_1_101001111010;
      patterns[27115] = 29'b0_110100111101_011_1_010011110101;
      patterns[27116] = 29'b0_110100111101_100_1_011010011110;
      patterns[27117] = 29'b0_110100111101_101_0_101101001111;
      patterns[27118] = 29'b0_110100111101_110_0_110100111101;
      patterns[27119] = 29'b0_110100111101_111_0_110100111101;
      patterns[27120] = 29'b0_110100111110_000_0_110100111110;
      patterns[27121] = 29'b0_110100111110_001_0_111110110100;
      patterns[27122] = 29'b0_110100111110_010_1_101001111100;
      patterns[27123] = 29'b0_110100111110_011_1_010011111001;
      patterns[27124] = 29'b0_110100111110_100_0_011010011111;
      patterns[27125] = 29'b0_110100111110_101_1_001101001111;
      patterns[27126] = 29'b0_110100111110_110_0_110100111110;
      patterns[27127] = 29'b0_110100111110_111_0_110100111110;
      patterns[27128] = 29'b0_110100111111_000_0_110100111111;
      patterns[27129] = 29'b0_110100111111_001_0_111111110100;
      patterns[27130] = 29'b0_110100111111_010_1_101001111110;
      patterns[27131] = 29'b0_110100111111_011_1_010011111101;
      patterns[27132] = 29'b0_110100111111_100_1_011010011111;
      patterns[27133] = 29'b0_110100111111_101_1_101101001111;
      patterns[27134] = 29'b0_110100111111_110_0_110100111111;
      patterns[27135] = 29'b0_110100111111_111_0_110100111111;
      patterns[27136] = 29'b0_110101000000_000_0_110101000000;
      patterns[27137] = 29'b0_110101000000_001_0_000000110101;
      patterns[27138] = 29'b0_110101000000_010_1_101010000000;
      patterns[27139] = 29'b0_110101000000_011_1_010100000001;
      patterns[27140] = 29'b0_110101000000_100_0_011010100000;
      patterns[27141] = 29'b0_110101000000_101_0_001101010000;
      patterns[27142] = 29'b0_110101000000_110_0_110101000000;
      patterns[27143] = 29'b0_110101000000_111_0_110101000000;
      patterns[27144] = 29'b0_110101000001_000_0_110101000001;
      patterns[27145] = 29'b0_110101000001_001_0_000001110101;
      patterns[27146] = 29'b0_110101000001_010_1_101010000010;
      patterns[27147] = 29'b0_110101000001_011_1_010100000101;
      patterns[27148] = 29'b0_110101000001_100_1_011010100000;
      patterns[27149] = 29'b0_110101000001_101_0_101101010000;
      patterns[27150] = 29'b0_110101000001_110_0_110101000001;
      patterns[27151] = 29'b0_110101000001_111_0_110101000001;
      patterns[27152] = 29'b0_110101000010_000_0_110101000010;
      patterns[27153] = 29'b0_110101000010_001_0_000010110101;
      patterns[27154] = 29'b0_110101000010_010_1_101010000100;
      patterns[27155] = 29'b0_110101000010_011_1_010100001001;
      patterns[27156] = 29'b0_110101000010_100_0_011010100001;
      patterns[27157] = 29'b0_110101000010_101_1_001101010000;
      patterns[27158] = 29'b0_110101000010_110_0_110101000010;
      patterns[27159] = 29'b0_110101000010_111_0_110101000010;
      patterns[27160] = 29'b0_110101000011_000_0_110101000011;
      patterns[27161] = 29'b0_110101000011_001_0_000011110101;
      patterns[27162] = 29'b0_110101000011_010_1_101010000110;
      patterns[27163] = 29'b0_110101000011_011_1_010100001101;
      patterns[27164] = 29'b0_110101000011_100_1_011010100001;
      patterns[27165] = 29'b0_110101000011_101_1_101101010000;
      patterns[27166] = 29'b0_110101000011_110_0_110101000011;
      patterns[27167] = 29'b0_110101000011_111_0_110101000011;
      patterns[27168] = 29'b0_110101000100_000_0_110101000100;
      patterns[27169] = 29'b0_110101000100_001_0_000100110101;
      patterns[27170] = 29'b0_110101000100_010_1_101010001000;
      patterns[27171] = 29'b0_110101000100_011_1_010100010001;
      patterns[27172] = 29'b0_110101000100_100_0_011010100010;
      patterns[27173] = 29'b0_110101000100_101_0_001101010001;
      patterns[27174] = 29'b0_110101000100_110_0_110101000100;
      patterns[27175] = 29'b0_110101000100_111_0_110101000100;
      patterns[27176] = 29'b0_110101000101_000_0_110101000101;
      patterns[27177] = 29'b0_110101000101_001_0_000101110101;
      patterns[27178] = 29'b0_110101000101_010_1_101010001010;
      patterns[27179] = 29'b0_110101000101_011_1_010100010101;
      patterns[27180] = 29'b0_110101000101_100_1_011010100010;
      patterns[27181] = 29'b0_110101000101_101_0_101101010001;
      patterns[27182] = 29'b0_110101000101_110_0_110101000101;
      patterns[27183] = 29'b0_110101000101_111_0_110101000101;
      patterns[27184] = 29'b0_110101000110_000_0_110101000110;
      patterns[27185] = 29'b0_110101000110_001_0_000110110101;
      patterns[27186] = 29'b0_110101000110_010_1_101010001100;
      patterns[27187] = 29'b0_110101000110_011_1_010100011001;
      patterns[27188] = 29'b0_110101000110_100_0_011010100011;
      patterns[27189] = 29'b0_110101000110_101_1_001101010001;
      patterns[27190] = 29'b0_110101000110_110_0_110101000110;
      patterns[27191] = 29'b0_110101000110_111_0_110101000110;
      patterns[27192] = 29'b0_110101000111_000_0_110101000111;
      patterns[27193] = 29'b0_110101000111_001_0_000111110101;
      patterns[27194] = 29'b0_110101000111_010_1_101010001110;
      patterns[27195] = 29'b0_110101000111_011_1_010100011101;
      patterns[27196] = 29'b0_110101000111_100_1_011010100011;
      patterns[27197] = 29'b0_110101000111_101_1_101101010001;
      patterns[27198] = 29'b0_110101000111_110_0_110101000111;
      patterns[27199] = 29'b0_110101000111_111_0_110101000111;
      patterns[27200] = 29'b0_110101001000_000_0_110101001000;
      patterns[27201] = 29'b0_110101001000_001_0_001000110101;
      patterns[27202] = 29'b0_110101001000_010_1_101010010000;
      patterns[27203] = 29'b0_110101001000_011_1_010100100001;
      patterns[27204] = 29'b0_110101001000_100_0_011010100100;
      patterns[27205] = 29'b0_110101001000_101_0_001101010010;
      patterns[27206] = 29'b0_110101001000_110_0_110101001000;
      patterns[27207] = 29'b0_110101001000_111_0_110101001000;
      patterns[27208] = 29'b0_110101001001_000_0_110101001001;
      patterns[27209] = 29'b0_110101001001_001_0_001001110101;
      patterns[27210] = 29'b0_110101001001_010_1_101010010010;
      patterns[27211] = 29'b0_110101001001_011_1_010100100101;
      patterns[27212] = 29'b0_110101001001_100_1_011010100100;
      patterns[27213] = 29'b0_110101001001_101_0_101101010010;
      patterns[27214] = 29'b0_110101001001_110_0_110101001001;
      patterns[27215] = 29'b0_110101001001_111_0_110101001001;
      patterns[27216] = 29'b0_110101001010_000_0_110101001010;
      patterns[27217] = 29'b0_110101001010_001_0_001010110101;
      patterns[27218] = 29'b0_110101001010_010_1_101010010100;
      patterns[27219] = 29'b0_110101001010_011_1_010100101001;
      patterns[27220] = 29'b0_110101001010_100_0_011010100101;
      patterns[27221] = 29'b0_110101001010_101_1_001101010010;
      patterns[27222] = 29'b0_110101001010_110_0_110101001010;
      patterns[27223] = 29'b0_110101001010_111_0_110101001010;
      patterns[27224] = 29'b0_110101001011_000_0_110101001011;
      patterns[27225] = 29'b0_110101001011_001_0_001011110101;
      patterns[27226] = 29'b0_110101001011_010_1_101010010110;
      patterns[27227] = 29'b0_110101001011_011_1_010100101101;
      patterns[27228] = 29'b0_110101001011_100_1_011010100101;
      patterns[27229] = 29'b0_110101001011_101_1_101101010010;
      patterns[27230] = 29'b0_110101001011_110_0_110101001011;
      patterns[27231] = 29'b0_110101001011_111_0_110101001011;
      patterns[27232] = 29'b0_110101001100_000_0_110101001100;
      patterns[27233] = 29'b0_110101001100_001_0_001100110101;
      patterns[27234] = 29'b0_110101001100_010_1_101010011000;
      patterns[27235] = 29'b0_110101001100_011_1_010100110001;
      patterns[27236] = 29'b0_110101001100_100_0_011010100110;
      patterns[27237] = 29'b0_110101001100_101_0_001101010011;
      patterns[27238] = 29'b0_110101001100_110_0_110101001100;
      patterns[27239] = 29'b0_110101001100_111_0_110101001100;
      patterns[27240] = 29'b0_110101001101_000_0_110101001101;
      patterns[27241] = 29'b0_110101001101_001_0_001101110101;
      patterns[27242] = 29'b0_110101001101_010_1_101010011010;
      patterns[27243] = 29'b0_110101001101_011_1_010100110101;
      patterns[27244] = 29'b0_110101001101_100_1_011010100110;
      patterns[27245] = 29'b0_110101001101_101_0_101101010011;
      patterns[27246] = 29'b0_110101001101_110_0_110101001101;
      patterns[27247] = 29'b0_110101001101_111_0_110101001101;
      patterns[27248] = 29'b0_110101001110_000_0_110101001110;
      patterns[27249] = 29'b0_110101001110_001_0_001110110101;
      patterns[27250] = 29'b0_110101001110_010_1_101010011100;
      patterns[27251] = 29'b0_110101001110_011_1_010100111001;
      patterns[27252] = 29'b0_110101001110_100_0_011010100111;
      patterns[27253] = 29'b0_110101001110_101_1_001101010011;
      patterns[27254] = 29'b0_110101001110_110_0_110101001110;
      patterns[27255] = 29'b0_110101001110_111_0_110101001110;
      patterns[27256] = 29'b0_110101001111_000_0_110101001111;
      patterns[27257] = 29'b0_110101001111_001_0_001111110101;
      patterns[27258] = 29'b0_110101001111_010_1_101010011110;
      patterns[27259] = 29'b0_110101001111_011_1_010100111101;
      patterns[27260] = 29'b0_110101001111_100_1_011010100111;
      patterns[27261] = 29'b0_110101001111_101_1_101101010011;
      patterns[27262] = 29'b0_110101001111_110_0_110101001111;
      patterns[27263] = 29'b0_110101001111_111_0_110101001111;
      patterns[27264] = 29'b0_110101010000_000_0_110101010000;
      patterns[27265] = 29'b0_110101010000_001_0_010000110101;
      patterns[27266] = 29'b0_110101010000_010_1_101010100000;
      patterns[27267] = 29'b0_110101010000_011_1_010101000001;
      patterns[27268] = 29'b0_110101010000_100_0_011010101000;
      patterns[27269] = 29'b0_110101010000_101_0_001101010100;
      patterns[27270] = 29'b0_110101010000_110_0_110101010000;
      patterns[27271] = 29'b0_110101010000_111_0_110101010000;
      patterns[27272] = 29'b0_110101010001_000_0_110101010001;
      patterns[27273] = 29'b0_110101010001_001_0_010001110101;
      patterns[27274] = 29'b0_110101010001_010_1_101010100010;
      patterns[27275] = 29'b0_110101010001_011_1_010101000101;
      patterns[27276] = 29'b0_110101010001_100_1_011010101000;
      patterns[27277] = 29'b0_110101010001_101_0_101101010100;
      patterns[27278] = 29'b0_110101010001_110_0_110101010001;
      patterns[27279] = 29'b0_110101010001_111_0_110101010001;
      patterns[27280] = 29'b0_110101010010_000_0_110101010010;
      patterns[27281] = 29'b0_110101010010_001_0_010010110101;
      patterns[27282] = 29'b0_110101010010_010_1_101010100100;
      patterns[27283] = 29'b0_110101010010_011_1_010101001001;
      patterns[27284] = 29'b0_110101010010_100_0_011010101001;
      patterns[27285] = 29'b0_110101010010_101_1_001101010100;
      patterns[27286] = 29'b0_110101010010_110_0_110101010010;
      patterns[27287] = 29'b0_110101010010_111_0_110101010010;
      patterns[27288] = 29'b0_110101010011_000_0_110101010011;
      patterns[27289] = 29'b0_110101010011_001_0_010011110101;
      patterns[27290] = 29'b0_110101010011_010_1_101010100110;
      patterns[27291] = 29'b0_110101010011_011_1_010101001101;
      patterns[27292] = 29'b0_110101010011_100_1_011010101001;
      patterns[27293] = 29'b0_110101010011_101_1_101101010100;
      patterns[27294] = 29'b0_110101010011_110_0_110101010011;
      patterns[27295] = 29'b0_110101010011_111_0_110101010011;
      patterns[27296] = 29'b0_110101010100_000_0_110101010100;
      patterns[27297] = 29'b0_110101010100_001_0_010100110101;
      patterns[27298] = 29'b0_110101010100_010_1_101010101000;
      patterns[27299] = 29'b0_110101010100_011_1_010101010001;
      patterns[27300] = 29'b0_110101010100_100_0_011010101010;
      patterns[27301] = 29'b0_110101010100_101_0_001101010101;
      patterns[27302] = 29'b0_110101010100_110_0_110101010100;
      patterns[27303] = 29'b0_110101010100_111_0_110101010100;
      patterns[27304] = 29'b0_110101010101_000_0_110101010101;
      patterns[27305] = 29'b0_110101010101_001_0_010101110101;
      patterns[27306] = 29'b0_110101010101_010_1_101010101010;
      patterns[27307] = 29'b0_110101010101_011_1_010101010101;
      patterns[27308] = 29'b0_110101010101_100_1_011010101010;
      patterns[27309] = 29'b0_110101010101_101_0_101101010101;
      patterns[27310] = 29'b0_110101010101_110_0_110101010101;
      patterns[27311] = 29'b0_110101010101_111_0_110101010101;
      patterns[27312] = 29'b0_110101010110_000_0_110101010110;
      patterns[27313] = 29'b0_110101010110_001_0_010110110101;
      patterns[27314] = 29'b0_110101010110_010_1_101010101100;
      patterns[27315] = 29'b0_110101010110_011_1_010101011001;
      patterns[27316] = 29'b0_110101010110_100_0_011010101011;
      patterns[27317] = 29'b0_110101010110_101_1_001101010101;
      patterns[27318] = 29'b0_110101010110_110_0_110101010110;
      patterns[27319] = 29'b0_110101010110_111_0_110101010110;
      patterns[27320] = 29'b0_110101010111_000_0_110101010111;
      patterns[27321] = 29'b0_110101010111_001_0_010111110101;
      patterns[27322] = 29'b0_110101010111_010_1_101010101110;
      patterns[27323] = 29'b0_110101010111_011_1_010101011101;
      patterns[27324] = 29'b0_110101010111_100_1_011010101011;
      patterns[27325] = 29'b0_110101010111_101_1_101101010101;
      patterns[27326] = 29'b0_110101010111_110_0_110101010111;
      patterns[27327] = 29'b0_110101010111_111_0_110101010111;
      patterns[27328] = 29'b0_110101011000_000_0_110101011000;
      patterns[27329] = 29'b0_110101011000_001_0_011000110101;
      patterns[27330] = 29'b0_110101011000_010_1_101010110000;
      patterns[27331] = 29'b0_110101011000_011_1_010101100001;
      patterns[27332] = 29'b0_110101011000_100_0_011010101100;
      patterns[27333] = 29'b0_110101011000_101_0_001101010110;
      patterns[27334] = 29'b0_110101011000_110_0_110101011000;
      patterns[27335] = 29'b0_110101011000_111_0_110101011000;
      patterns[27336] = 29'b0_110101011001_000_0_110101011001;
      patterns[27337] = 29'b0_110101011001_001_0_011001110101;
      patterns[27338] = 29'b0_110101011001_010_1_101010110010;
      patterns[27339] = 29'b0_110101011001_011_1_010101100101;
      patterns[27340] = 29'b0_110101011001_100_1_011010101100;
      patterns[27341] = 29'b0_110101011001_101_0_101101010110;
      patterns[27342] = 29'b0_110101011001_110_0_110101011001;
      patterns[27343] = 29'b0_110101011001_111_0_110101011001;
      patterns[27344] = 29'b0_110101011010_000_0_110101011010;
      patterns[27345] = 29'b0_110101011010_001_0_011010110101;
      patterns[27346] = 29'b0_110101011010_010_1_101010110100;
      patterns[27347] = 29'b0_110101011010_011_1_010101101001;
      patterns[27348] = 29'b0_110101011010_100_0_011010101101;
      patterns[27349] = 29'b0_110101011010_101_1_001101010110;
      patterns[27350] = 29'b0_110101011010_110_0_110101011010;
      patterns[27351] = 29'b0_110101011010_111_0_110101011010;
      patterns[27352] = 29'b0_110101011011_000_0_110101011011;
      patterns[27353] = 29'b0_110101011011_001_0_011011110101;
      patterns[27354] = 29'b0_110101011011_010_1_101010110110;
      patterns[27355] = 29'b0_110101011011_011_1_010101101101;
      patterns[27356] = 29'b0_110101011011_100_1_011010101101;
      patterns[27357] = 29'b0_110101011011_101_1_101101010110;
      patterns[27358] = 29'b0_110101011011_110_0_110101011011;
      patterns[27359] = 29'b0_110101011011_111_0_110101011011;
      patterns[27360] = 29'b0_110101011100_000_0_110101011100;
      patterns[27361] = 29'b0_110101011100_001_0_011100110101;
      patterns[27362] = 29'b0_110101011100_010_1_101010111000;
      patterns[27363] = 29'b0_110101011100_011_1_010101110001;
      patterns[27364] = 29'b0_110101011100_100_0_011010101110;
      patterns[27365] = 29'b0_110101011100_101_0_001101010111;
      patterns[27366] = 29'b0_110101011100_110_0_110101011100;
      patterns[27367] = 29'b0_110101011100_111_0_110101011100;
      patterns[27368] = 29'b0_110101011101_000_0_110101011101;
      patterns[27369] = 29'b0_110101011101_001_0_011101110101;
      patterns[27370] = 29'b0_110101011101_010_1_101010111010;
      patterns[27371] = 29'b0_110101011101_011_1_010101110101;
      patterns[27372] = 29'b0_110101011101_100_1_011010101110;
      patterns[27373] = 29'b0_110101011101_101_0_101101010111;
      patterns[27374] = 29'b0_110101011101_110_0_110101011101;
      patterns[27375] = 29'b0_110101011101_111_0_110101011101;
      patterns[27376] = 29'b0_110101011110_000_0_110101011110;
      patterns[27377] = 29'b0_110101011110_001_0_011110110101;
      patterns[27378] = 29'b0_110101011110_010_1_101010111100;
      patterns[27379] = 29'b0_110101011110_011_1_010101111001;
      patterns[27380] = 29'b0_110101011110_100_0_011010101111;
      patterns[27381] = 29'b0_110101011110_101_1_001101010111;
      patterns[27382] = 29'b0_110101011110_110_0_110101011110;
      patterns[27383] = 29'b0_110101011110_111_0_110101011110;
      patterns[27384] = 29'b0_110101011111_000_0_110101011111;
      patterns[27385] = 29'b0_110101011111_001_0_011111110101;
      patterns[27386] = 29'b0_110101011111_010_1_101010111110;
      patterns[27387] = 29'b0_110101011111_011_1_010101111101;
      patterns[27388] = 29'b0_110101011111_100_1_011010101111;
      patterns[27389] = 29'b0_110101011111_101_1_101101010111;
      patterns[27390] = 29'b0_110101011111_110_0_110101011111;
      patterns[27391] = 29'b0_110101011111_111_0_110101011111;
      patterns[27392] = 29'b0_110101100000_000_0_110101100000;
      patterns[27393] = 29'b0_110101100000_001_0_100000110101;
      patterns[27394] = 29'b0_110101100000_010_1_101011000000;
      patterns[27395] = 29'b0_110101100000_011_1_010110000001;
      patterns[27396] = 29'b0_110101100000_100_0_011010110000;
      patterns[27397] = 29'b0_110101100000_101_0_001101011000;
      patterns[27398] = 29'b0_110101100000_110_0_110101100000;
      patterns[27399] = 29'b0_110101100000_111_0_110101100000;
      patterns[27400] = 29'b0_110101100001_000_0_110101100001;
      patterns[27401] = 29'b0_110101100001_001_0_100001110101;
      patterns[27402] = 29'b0_110101100001_010_1_101011000010;
      patterns[27403] = 29'b0_110101100001_011_1_010110000101;
      patterns[27404] = 29'b0_110101100001_100_1_011010110000;
      patterns[27405] = 29'b0_110101100001_101_0_101101011000;
      patterns[27406] = 29'b0_110101100001_110_0_110101100001;
      patterns[27407] = 29'b0_110101100001_111_0_110101100001;
      patterns[27408] = 29'b0_110101100010_000_0_110101100010;
      patterns[27409] = 29'b0_110101100010_001_0_100010110101;
      patterns[27410] = 29'b0_110101100010_010_1_101011000100;
      patterns[27411] = 29'b0_110101100010_011_1_010110001001;
      patterns[27412] = 29'b0_110101100010_100_0_011010110001;
      patterns[27413] = 29'b0_110101100010_101_1_001101011000;
      patterns[27414] = 29'b0_110101100010_110_0_110101100010;
      patterns[27415] = 29'b0_110101100010_111_0_110101100010;
      patterns[27416] = 29'b0_110101100011_000_0_110101100011;
      patterns[27417] = 29'b0_110101100011_001_0_100011110101;
      patterns[27418] = 29'b0_110101100011_010_1_101011000110;
      patterns[27419] = 29'b0_110101100011_011_1_010110001101;
      patterns[27420] = 29'b0_110101100011_100_1_011010110001;
      patterns[27421] = 29'b0_110101100011_101_1_101101011000;
      patterns[27422] = 29'b0_110101100011_110_0_110101100011;
      patterns[27423] = 29'b0_110101100011_111_0_110101100011;
      patterns[27424] = 29'b0_110101100100_000_0_110101100100;
      patterns[27425] = 29'b0_110101100100_001_0_100100110101;
      patterns[27426] = 29'b0_110101100100_010_1_101011001000;
      patterns[27427] = 29'b0_110101100100_011_1_010110010001;
      patterns[27428] = 29'b0_110101100100_100_0_011010110010;
      patterns[27429] = 29'b0_110101100100_101_0_001101011001;
      patterns[27430] = 29'b0_110101100100_110_0_110101100100;
      patterns[27431] = 29'b0_110101100100_111_0_110101100100;
      patterns[27432] = 29'b0_110101100101_000_0_110101100101;
      patterns[27433] = 29'b0_110101100101_001_0_100101110101;
      patterns[27434] = 29'b0_110101100101_010_1_101011001010;
      patterns[27435] = 29'b0_110101100101_011_1_010110010101;
      patterns[27436] = 29'b0_110101100101_100_1_011010110010;
      patterns[27437] = 29'b0_110101100101_101_0_101101011001;
      patterns[27438] = 29'b0_110101100101_110_0_110101100101;
      patterns[27439] = 29'b0_110101100101_111_0_110101100101;
      patterns[27440] = 29'b0_110101100110_000_0_110101100110;
      patterns[27441] = 29'b0_110101100110_001_0_100110110101;
      patterns[27442] = 29'b0_110101100110_010_1_101011001100;
      patterns[27443] = 29'b0_110101100110_011_1_010110011001;
      patterns[27444] = 29'b0_110101100110_100_0_011010110011;
      patterns[27445] = 29'b0_110101100110_101_1_001101011001;
      patterns[27446] = 29'b0_110101100110_110_0_110101100110;
      patterns[27447] = 29'b0_110101100110_111_0_110101100110;
      patterns[27448] = 29'b0_110101100111_000_0_110101100111;
      patterns[27449] = 29'b0_110101100111_001_0_100111110101;
      patterns[27450] = 29'b0_110101100111_010_1_101011001110;
      patterns[27451] = 29'b0_110101100111_011_1_010110011101;
      patterns[27452] = 29'b0_110101100111_100_1_011010110011;
      patterns[27453] = 29'b0_110101100111_101_1_101101011001;
      patterns[27454] = 29'b0_110101100111_110_0_110101100111;
      patterns[27455] = 29'b0_110101100111_111_0_110101100111;
      patterns[27456] = 29'b0_110101101000_000_0_110101101000;
      patterns[27457] = 29'b0_110101101000_001_0_101000110101;
      patterns[27458] = 29'b0_110101101000_010_1_101011010000;
      patterns[27459] = 29'b0_110101101000_011_1_010110100001;
      patterns[27460] = 29'b0_110101101000_100_0_011010110100;
      patterns[27461] = 29'b0_110101101000_101_0_001101011010;
      patterns[27462] = 29'b0_110101101000_110_0_110101101000;
      patterns[27463] = 29'b0_110101101000_111_0_110101101000;
      patterns[27464] = 29'b0_110101101001_000_0_110101101001;
      patterns[27465] = 29'b0_110101101001_001_0_101001110101;
      patterns[27466] = 29'b0_110101101001_010_1_101011010010;
      patterns[27467] = 29'b0_110101101001_011_1_010110100101;
      patterns[27468] = 29'b0_110101101001_100_1_011010110100;
      patterns[27469] = 29'b0_110101101001_101_0_101101011010;
      patterns[27470] = 29'b0_110101101001_110_0_110101101001;
      patterns[27471] = 29'b0_110101101001_111_0_110101101001;
      patterns[27472] = 29'b0_110101101010_000_0_110101101010;
      patterns[27473] = 29'b0_110101101010_001_0_101010110101;
      patterns[27474] = 29'b0_110101101010_010_1_101011010100;
      patterns[27475] = 29'b0_110101101010_011_1_010110101001;
      patterns[27476] = 29'b0_110101101010_100_0_011010110101;
      patterns[27477] = 29'b0_110101101010_101_1_001101011010;
      patterns[27478] = 29'b0_110101101010_110_0_110101101010;
      patterns[27479] = 29'b0_110101101010_111_0_110101101010;
      patterns[27480] = 29'b0_110101101011_000_0_110101101011;
      patterns[27481] = 29'b0_110101101011_001_0_101011110101;
      patterns[27482] = 29'b0_110101101011_010_1_101011010110;
      patterns[27483] = 29'b0_110101101011_011_1_010110101101;
      patterns[27484] = 29'b0_110101101011_100_1_011010110101;
      patterns[27485] = 29'b0_110101101011_101_1_101101011010;
      patterns[27486] = 29'b0_110101101011_110_0_110101101011;
      patterns[27487] = 29'b0_110101101011_111_0_110101101011;
      patterns[27488] = 29'b0_110101101100_000_0_110101101100;
      patterns[27489] = 29'b0_110101101100_001_0_101100110101;
      patterns[27490] = 29'b0_110101101100_010_1_101011011000;
      patterns[27491] = 29'b0_110101101100_011_1_010110110001;
      patterns[27492] = 29'b0_110101101100_100_0_011010110110;
      patterns[27493] = 29'b0_110101101100_101_0_001101011011;
      patterns[27494] = 29'b0_110101101100_110_0_110101101100;
      patterns[27495] = 29'b0_110101101100_111_0_110101101100;
      patterns[27496] = 29'b0_110101101101_000_0_110101101101;
      patterns[27497] = 29'b0_110101101101_001_0_101101110101;
      patterns[27498] = 29'b0_110101101101_010_1_101011011010;
      patterns[27499] = 29'b0_110101101101_011_1_010110110101;
      patterns[27500] = 29'b0_110101101101_100_1_011010110110;
      patterns[27501] = 29'b0_110101101101_101_0_101101011011;
      patterns[27502] = 29'b0_110101101101_110_0_110101101101;
      patterns[27503] = 29'b0_110101101101_111_0_110101101101;
      patterns[27504] = 29'b0_110101101110_000_0_110101101110;
      patterns[27505] = 29'b0_110101101110_001_0_101110110101;
      patterns[27506] = 29'b0_110101101110_010_1_101011011100;
      patterns[27507] = 29'b0_110101101110_011_1_010110111001;
      patterns[27508] = 29'b0_110101101110_100_0_011010110111;
      patterns[27509] = 29'b0_110101101110_101_1_001101011011;
      patterns[27510] = 29'b0_110101101110_110_0_110101101110;
      patterns[27511] = 29'b0_110101101110_111_0_110101101110;
      patterns[27512] = 29'b0_110101101111_000_0_110101101111;
      patterns[27513] = 29'b0_110101101111_001_0_101111110101;
      patterns[27514] = 29'b0_110101101111_010_1_101011011110;
      patterns[27515] = 29'b0_110101101111_011_1_010110111101;
      patterns[27516] = 29'b0_110101101111_100_1_011010110111;
      patterns[27517] = 29'b0_110101101111_101_1_101101011011;
      patterns[27518] = 29'b0_110101101111_110_0_110101101111;
      patterns[27519] = 29'b0_110101101111_111_0_110101101111;
      patterns[27520] = 29'b0_110101110000_000_0_110101110000;
      patterns[27521] = 29'b0_110101110000_001_0_110000110101;
      patterns[27522] = 29'b0_110101110000_010_1_101011100000;
      patterns[27523] = 29'b0_110101110000_011_1_010111000001;
      patterns[27524] = 29'b0_110101110000_100_0_011010111000;
      patterns[27525] = 29'b0_110101110000_101_0_001101011100;
      patterns[27526] = 29'b0_110101110000_110_0_110101110000;
      patterns[27527] = 29'b0_110101110000_111_0_110101110000;
      patterns[27528] = 29'b0_110101110001_000_0_110101110001;
      patterns[27529] = 29'b0_110101110001_001_0_110001110101;
      patterns[27530] = 29'b0_110101110001_010_1_101011100010;
      patterns[27531] = 29'b0_110101110001_011_1_010111000101;
      patterns[27532] = 29'b0_110101110001_100_1_011010111000;
      patterns[27533] = 29'b0_110101110001_101_0_101101011100;
      patterns[27534] = 29'b0_110101110001_110_0_110101110001;
      patterns[27535] = 29'b0_110101110001_111_0_110101110001;
      patterns[27536] = 29'b0_110101110010_000_0_110101110010;
      patterns[27537] = 29'b0_110101110010_001_0_110010110101;
      patterns[27538] = 29'b0_110101110010_010_1_101011100100;
      patterns[27539] = 29'b0_110101110010_011_1_010111001001;
      patterns[27540] = 29'b0_110101110010_100_0_011010111001;
      patterns[27541] = 29'b0_110101110010_101_1_001101011100;
      patterns[27542] = 29'b0_110101110010_110_0_110101110010;
      patterns[27543] = 29'b0_110101110010_111_0_110101110010;
      patterns[27544] = 29'b0_110101110011_000_0_110101110011;
      patterns[27545] = 29'b0_110101110011_001_0_110011110101;
      patterns[27546] = 29'b0_110101110011_010_1_101011100110;
      patterns[27547] = 29'b0_110101110011_011_1_010111001101;
      patterns[27548] = 29'b0_110101110011_100_1_011010111001;
      patterns[27549] = 29'b0_110101110011_101_1_101101011100;
      patterns[27550] = 29'b0_110101110011_110_0_110101110011;
      patterns[27551] = 29'b0_110101110011_111_0_110101110011;
      patterns[27552] = 29'b0_110101110100_000_0_110101110100;
      patterns[27553] = 29'b0_110101110100_001_0_110100110101;
      patterns[27554] = 29'b0_110101110100_010_1_101011101000;
      patterns[27555] = 29'b0_110101110100_011_1_010111010001;
      patterns[27556] = 29'b0_110101110100_100_0_011010111010;
      patterns[27557] = 29'b0_110101110100_101_0_001101011101;
      patterns[27558] = 29'b0_110101110100_110_0_110101110100;
      patterns[27559] = 29'b0_110101110100_111_0_110101110100;
      patterns[27560] = 29'b0_110101110101_000_0_110101110101;
      patterns[27561] = 29'b0_110101110101_001_0_110101110101;
      patterns[27562] = 29'b0_110101110101_010_1_101011101010;
      patterns[27563] = 29'b0_110101110101_011_1_010111010101;
      patterns[27564] = 29'b0_110101110101_100_1_011010111010;
      patterns[27565] = 29'b0_110101110101_101_0_101101011101;
      patterns[27566] = 29'b0_110101110101_110_0_110101110101;
      patterns[27567] = 29'b0_110101110101_111_0_110101110101;
      patterns[27568] = 29'b0_110101110110_000_0_110101110110;
      patterns[27569] = 29'b0_110101110110_001_0_110110110101;
      patterns[27570] = 29'b0_110101110110_010_1_101011101100;
      patterns[27571] = 29'b0_110101110110_011_1_010111011001;
      patterns[27572] = 29'b0_110101110110_100_0_011010111011;
      patterns[27573] = 29'b0_110101110110_101_1_001101011101;
      patterns[27574] = 29'b0_110101110110_110_0_110101110110;
      patterns[27575] = 29'b0_110101110110_111_0_110101110110;
      patterns[27576] = 29'b0_110101110111_000_0_110101110111;
      patterns[27577] = 29'b0_110101110111_001_0_110111110101;
      patterns[27578] = 29'b0_110101110111_010_1_101011101110;
      patterns[27579] = 29'b0_110101110111_011_1_010111011101;
      patterns[27580] = 29'b0_110101110111_100_1_011010111011;
      patterns[27581] = 29'b0_110101110111_101_1_101101011101;
      patterns[27582] = 29'b0_110101110111_110_0_110101110111;
      patterns[27583] = 29'b0_110101110111_111_0_110101110111;
      patterns[27584] = 29'b0_110101111000_000_0_110101111000;
      patterns[27585] = 29'b0_110101111000_001_0_111000110101;
      patterns[27586] = 29'b0_110101111000_010_1_101011110000;
      patterns[27587] = 29'b0_110101111000_011_1_010111100001;
      patterns[27588] = 29'b0_110101111000_100_0_011010111100;
      patterns[27589] = 29'b0_110101111000_101_0_001101011110;
      patterns[27590] = 29'b0_110101111000_110_0_110101111000;
      patterns[27591] = 29'b0_110101111000_111_0_110101111000;
      patterns[27592] = 29'b0_110101111001_000_0_110101111001;
      patterns[27593] = 29'b0_110101111001_001_0_111001110101;
      patterns[27594] = 29'b0_110101111001_010_1_101011110010;
      patterns[27595] = 29'b0_110101111001_011_1_010111100101;
      patterns[27596] = 29'b0_110101111001_100_1_011010111100;
      patterns[27597] = 29'b0_110101111001_101_0_101101011110;
      patterns[27598] = 29'b0_110101111001_110_0_110101111001;
      patterns[27599] = 29'b0_110101111001_111_0_110101111001;
      patterns[27600] = 29'b0_110101111010_000_0_110101111010;
      patterns[27601] = 29'b0_110101111010_001_0_111010110101;
      patterns[27602] = 29'b0_110101111010_010_1_101011110100;
      patterns[27603] = 29'b0_110101111010_011_1_010111101001;
      patterns[27604] = 29'b0_110101111010_100_0_011010111101;
      patterns[27605] = 29'b0_110101111010_101_1_001101011110;
      patterns[27606] = 29'b0_110101111010_110_0_110101111010;
      patterns[27607] = 29'b0_110101111010_111_0_110101111010;
      patterns[27608] = 29'b0_110101111011_000_0_110101111011;
      patterns[27609] = 29'b0_110101111011_001_0_111011110101;
      patterns[27610] = 29'b0_110101111011_010_1_101011110110;
      patterns[27611] = 29'b0_110101111011_011_1_010111101101;
      patterns[27612] = 29'b0_110101111011_100_1_011010111101;
      patterns[27613] = 29'b0_110101111011_101_1_101101011110;
      patterns[27614] = 29'b0_110101111011_110_0_110101111011;
      patterns[27615] = 29'b0_110101111011_111_0_110101111011;
      patterns[27616] = 29'b0_110101111100_000_0_110101111100;
      patterns[27617] = 29'b0_110101111100_001_0_111100110101;
      patterns[27618] = 29'b0_110101111100_010_1_101011111000;
      patterns[27619] = 29'b0_110101111100_011_1_010111110001;
      patterns[27620] = 29'b0_110101111100_100_0_011010111110;
      patterns[27621] = 29'b0_110101111100_101_0_001101011111;
      patterns[27622] = 29'b0_110101111100_110_0_110101111100;
      patterns[27623] = 29'b0_110101111100_111_0_110101111100;
      patterns[27624] = 29'b0_110101111101_000_0_110101111101;
      patterns[27625] = 29'b0_110101111101_001_0_111101110101;
      patterns[27626] = 29'b0_110101111101_010_1_101011111010;
      patterns[27627] = 29'b0_110101111101_011_1_010111110101;
      patterns[27628] = 29'b0_110101111101_100_1_011010111110;
      patterns[27629] = 29'b0_110101111101_101_0_101101011111;
      patterns[27630] = 29'b0_110101111101_110_0_110101111101;
      patterns[27631] = 29'b0_110101111101_111_0_110101111101;
      patterns[27632] = 29'b0_110101111110_000_0_110101111110;
      patterns[27633] = 29'b0_110101111110_001_0_111110110101;
      patterns[27634] = 29'b0_110101111110_010_1_101011111100;
      patterns[27635] = 29'b0_110101111110_011_1_010111111001;
      patterns[27636] = 29'b0_110101111110_100_0_011010111111;
      patterns[27637] = 29'b0_110101111110_101_1_001101011111;
      patterns[27638] = 29'b0_110101111110_110_0_110101111110;
      patterns[27639] = 29'b0_110101111110_111_0_110101111110;
      patterns[27640] = 29'b0_110101111111_000_0_110101111111;
      patterns[27641] = 29'b0_110101111111_001_0_111111110101;
      patterns[27642] = 29'b0_110101111111_010_1_101011111110;
      patterns[27643] = 29'b0_110101111111_011_1_010111111101;
      patterns[27644] = 29'b0_110101111111_100_1_011010111111;
      patterns[27645] = 29'b0_110101111111_101_1_101101011111;
      patterns[27646] = 29'b0_110101111111_110_0_110101111111;
      patterns[27647] = 29'b0_110101111111_111_0_110101111111;
      patterns[27648] = 29'b0_110110000000_000_0_110110000000;
      patterns[27649] = 29'b0_110110000000_001_0_000000110110;
      patterns[27650] = 29'b0_110110000000_010_1_101100000000;
      patterns[27651] = 29'b0_110110000000_011_1_011000000001;
      patterns[27652] = 29'b0_110110000000_100_0_011011000000;
      patterns[27653] = 29'b0_110110000000_101_0_001101100000;
      patterns[27654] = 29'b0_110110000000_110_0_110110000000;
      patterns[27655] = 29'b0_110110000000_111_0_110110000000;
      patterns[27656] = 29'b0_110110000001_000_0_110110000001;
      patterns[27657] = 29'b0_110110000001_001_0_000001110110;
      patterns[27658] = 29'b0_110110000001_010_1_101100000010;
      patterns[27659] = 29'b0_110110000001_011_1_011000000101;
      patterns[27660] = 29'b0_110110000001_100_1_011011000000;
      patterns[27661] = 29'b0_110110000001_101_0_101101100000;
      patterns[27662] = 29'b0_110110000001_110_0_110110000001;
      patterns[27663] = 29'b0_110110000001_111_0_110110000001;
      patterns[27664] = 29'b0_110110000010_000_0_110110000010;
      patterns[27665] = 29'b0_110110000010_001_0_000010110110;
      patterns[27666] = 29'b0_110110000010_010_1_101100000100;
      patterns[27667] = 29'b0_110110000010_011_1_011000001001;
      patterns[27668] = 29'b0_110110000010_100_0_011011000001;
      patterns[27669] = 29'b0_110110000010_101_1_001101100000;
      patterns[27670] = 29'b0_110110000010_110_0_110110000010;
      patterns[27671] = 29'b0_110110000010_111_0_110110000010;
      patterns[27672] = 29'b0_110110000011_000_0_110110000011;
      patterns[27673] = 29'b0_110110000011_001_0_000011110110;
      patterns[27674] = 29'b0_110110000011_010_1_101100000110;
      patterns[27675] = 29'b0_110110000011_011_1_011000001101;
      patterns[27676] = 29'b0_110110000011_100_1_011011000001;
      patterns[27677] = 29'b0_110110000011_101_1_101101100000;
      patterns[27678] = 29'b0_110110000011_110_0_110110000011;
      patterns[27679] = 29'b0_110110000011_111_0_110110000011;
      patterns[27680] = 29'b0_110110000100_000_0_110110000100;
      patterns[27681] = 29'b0_110110000100_001_0_000100110110;
      patterns[27682] = 29'b0_110110000100_010_1_101100001000;
      patterns[27683] = 29'b0_110110000100_011_1_011000010001;
      patterns[27684] = 29'b0_110110000100_100_0_011011000010;
      patterns[27685] = 29'b0_110110000100_101_0_001101100001;
      patterns[27686] = 29'b0_110110000100_110_0_110110000100;
      patterns[27687] = 29'b0_110110000100_111_0_110110000100;
      patterns[27688] = 29'b0_110110000101_000_0_110110000101;
      patterns[27689] = 29'b0_110110000101_001_0_000101110110;
      patterns[27690] = 29'b0_110110000101_010_1_101100001010;
      patterns[27691] = 29'b0_110110000101_011_1_011000010101;
      patterns[27692] = 29'b0_110110000101_100_1_011011000010;
      patterns[27693] = 29'b0_110110000101_101_0_101101100001;
      patterns[27694] = 29'b0_110110000101_110_0_110110000101;
      patterns[27695] = 29'b0_110110000101_111_0_110110000101;
      patterns[27696] = 29'b0_110110000110_000_0_110110000110;
      patterns[27697] = 29'b0_110110000110_001_0_000110110110;
      patterns[27698] = 29'b0_110110000110_010_1_101100001100;
      patterns[27699] = 29'b0_110110000110_011_1_011000011001;
      patterns[27700] = 29'b0_110110000110_100_0_011011000011;
      patterns[27701] = 29'b0_110110000110_101_1_001101100001;
      patterns[27702] = 29'b0_110110000110_110_0_110110000110;
      patterns[27703] = 29'b0_110110000110_111_0_110110000110;
      patterns[27704] = 29'b0_110110000111_000_0_110110000111;
      patterns[27705] = 29'b0_110110000111_001_0_000111110110;
      patterns[27706] = 29'b0_110110000111_010_1_101100001110;
      patterns[27707] = 29'b0_110110000111_011_1_011000011101;
      patterns[27708] = 29'b0_110110000111_100_1_011011000011;
      patterns[27709] = 29'b0_110110000111_101_1_101101100001;
      patterns[27710] = 29'b0_110110000111_110_0_110110000111;
      patterns[27711] = 29'b0_110110000111_111_0_110110000111;
      patterns[27712] = 29'b0_110110001000_000_0_110110001000;
      patterns[27713] = 29'b0_110110001000_001_0_001000110110;
      patterns[27714] = 29'b0_110110001000_010_1_101100010000;
      patterns[27715] = 29'b0_110110001000_011_1_011000100001;
      patterns[27716] = 29'b0_110110001000_100_0_011011000100;
      patterns[27717] = 29'b0_110110001000_101_0_001101100010;
      patterns[27718] = 29'b0_110110001000_110_0_110110001000;
      patterns[27719] = 29'b0_110110001000_111_0_110110001000;
      patterns[27720] = 29'b0_110110001001_000_0_110110001001;
      patterns[27721] = 29'b0_110110001001_001_0_001001110110;
      patterns[27722] = 29'b0_110110001001_010_1_101100010010;
      patterns[27723] = 29'b0_110110001001_011_1_011000100101;
      patterns[27724] = 29'b0_110110001001_100_1_011011000100;
      patterns[27725] = 29'b0_110110001001_101_0_101101100010;
      patterns[27726] = 29'b0_110110001001_110_0_110110001001;
      patterns[27727] = 29'b0_110110001001_111_0_110110001001;
      patterns[27728] = 29'b0_110110001010_000_0_110110001010;
      patterns[27729] = 29'b0_110110001010_001_0_001010110110;
      patterns[27730] = 29'b0_110110001010_010_1_101100010100;
      patterns[27731] = 29'b0_110110001010_011_1_011000101001;
      patterns[27732] = 29'b0_110110001010_100_0_011011000101;
      patterns[27733] = 29'b0_110110001010_101_1_001101100010;
      patterns[27734] = 29'b0_110110001010_110_0_110110001010;
      patterns[27735] = 29'b0_110110001010_111_0_110110001010;
      patterns[27736] = 29'b0_110110001011_000_0_110110001011;
      patterns[27737] = 29'b0_110110001011_001_0_001011110110;
      patterns[27738] = 29'b0_110110001011_010_1_101100010110;
      patterns[27739] = 29'b0_110110001011_011_1_011000101101;
      patterns[27740] = 29'b0_110110001011_100_1_011011000101;
      patterns[27741] = 29'b0_110110001011_101_1_101101100010;
      patterns[27742] = 29'b0_110110001011_110_0_110110001011;
      patterns[27743] = 29'b0_110110001011_111_0_110110001011;
      patterns[27744] = 29'b0_110110001100_000_0_110110001100;
      patterns[27745] = 29'b0_110110001100_001_0_001100110110;
      patterns[27746] = 29'b0_110110001100_010_1_101100011000;
      patterns[27747] = 29'b0_110110001100_011_1_011000110001;
      patterns[27748] = 29'b0_110110001100_100_0_011011000110;
      patterns[27749] = 29'b0_110110001100_101_0_001101100011;
      patterns[27750] = 29'b0_110110001100_110_0_110110001100;
      patterns[27751] = 29'b0_110110001100_111_0_110110001100;
      patterns[27752] = 29'b0_110110001101_000_0_110110001101;
      patterns[27753] = 29'b0_110110001101_001_0_001101110110;
      patterns[27754] = 29'b0_110110001101_010_1_101100011010;
      patterns[27755] = 29'b0_110110001101_011_1_011000110101;
      patterns[27756] = 29'b0_110110001101_100_1_011011000110;
      patterns[27757] = 29'b0_110110001101_101_0_101101100011;
      patterns[27758] = 29'b0_110110001101_110_0_110110001101;
      patterns[27759] = 29'b0_110110001101_111_0_110110001101;
      patterns[27760] = 29'b0_110110001110_000_0_110110001110;
      patterns[27761] = 29'b0_110110001110_001_0_001110110110;
      patterns[27762] = 29'b0_110110001110_010_1_101100011100;
      patterns[27763] = 29'b0_110110001110_011_1_011000111001;
      patterns[27764] = 29'b0_110110001110_100_0_011011000111;
      patterns[27765] = 29'b0_110110001110_101_1_001101100011;
      patterns[27766] = 29'b0_110110001110_110_0_110110001110;
      patterns[27767] = 29'b0_110110001110_111_0_110110001110;
      patterns[27768] = 29'b0_110110001111_000_0_110110001111;
      patterns[27769] = 29'b0_110110001111_001_0_001111110110;
      patterns[27770] = 29'b0_110110001111_010_1_101100011110;
      patterns[27771] = 29'b0_110110001111_011_1_011000111101;
      patterns[27772] = 29'b0_110110001111_100_1_011011000111;
      patterns[27773] = 29'b0_110110001111_101_1_101101100011;
      patterns[27774] = 29'b0_110110001111_110_0_110110001111;
      patterns[27775] = 29'b0_110110001111_111_0_110110001111;
      patterns[27776] = 29'b0_110110010000_000_0_110110010000;
      patterns[27777] = 29'b0_110110010000_001_0_010000110110;
      patterns[27778] = 29'b0_110110010000_010_1_101100100000;
      patterns[27779] = 29'b0_110110010000_011_1_011001000001;
      patterns[27780] = 29'b0_110110010000_100_0_011011001000;
      patterns[27781] = 29'b0_110110010000_101_0_001101100100;
      patterns[27782] = 29'b0_110110010000_110_0_110110010000;
      patterns[27783] = 29'b0_110110010000_111_0_110110010000;
      patterns[27784] = 29'b0_110110010001_000_0_110110010001;
      patterns[27785] = 29'b0_110110010001_001_0_010001110110;
      patterns[27786] = 29'b0_110110010001_010_1_101100100010;
      patterns[27787] = 29'b0_110110010001_011_1_011001000101;
      patterns[27788] = 29'b0_110110010001_100_1_011011001000;
      patterns[27789] = 29'b0_110110010001_101_0_101101100100;
      patterns[27790] = 29'b0_110110010001_110_0_110110010001;
      patterns[27791] = 29'b0_110110010001_111_0_110110010001;
      patterns[27792] = 29'b0_110110010010_000_0_110110010010;
      patterns[27793] = 29'b0_110110010010_001_0_010010110110;
      patterns[27794] = 29'b0_110110010010_010_1_101100100100;
      patterns[27795] = 29'b0_110110010010_011_1_011001001001;
      patterns[27796] = 29'b0_110110010010_100_0_011011001001;
      patterns[27797] = 29'b0_110110010010_101_1_001101100100;
      patterns[27798] = 29'b0_110110010010_110_0_110110010010;
      patterns[27799] = 29'b0_110110010010_111_0_110110010010;
      patterns[27800] = 29'b0_110110010011_000_0_110110010011;
      patterns[27801] = 29'b0_110110010011_001_0_010011110110;
      patterns[27802] = 29'b0_110110010011_010_1_101100100110;
      patterns[27803] = 29'b0_110110010011_011_1_011001001101;
      patterns[27804] = 29'b0_110110010011_100_1_011011001001;
      patterns[27805] = 29'b0_110110010011_101_1_101101100100;
      patterns[27806] = 29'b0_110110010011_110_0_110110010011;
      patterns[27807] = 29'b0_110110010011_111_0_110110010011;
      patterns[27808] = 29'b0_110110010100_000_0_110110010100;
      patterns[27809] = 29'b0_110110010100_001_0_010100110110;
      patterns[27810] = 29'b0_110110010100_010_1_101100101000;
      patterns[27811] = 29'b0_110110010100_011_1_011001010001;
      patterns[27812] = 29'b0_110110010100_100_0_011011001010;
      patterns[27813] = 29'b0_110110010100_101_0_001101100101;
      patterns[27814] = 29'b0_110110010100_110_0_110110010100;
      patterns[27815] = 29'b0_110110010100_111_0_110110010100;
      patterns[27816] = 29'b0_110110010101_000_0_110110010101;
      patterns[27817] = 29'b0_110110010101_001_0_010101110110;
      patterns[27818] = 29'b0_110110010101_010_1_101100101010;
      patterns[27819] = 29'b0_110110010101_011_1_011001010101;
      patterns[27820] = 29'b0_110110010101_100_1_011011001010;
      patterns[27821] = 29'b0_110110010101_101_0_101101100101;
      patterns[27822] = 29'b0_110110010101_110_0_110110010101;
      patterns[27823] = 29'b0_110110010101_111_0_110110010101;
      patterns[27824] = 29'b0_110110010110_000_0_110110010110;
      patterns[27825] = 29'b0_110110010110_001_0_010110110110;
      patterns[27826] = 29'b0_110110010110_010_1_101100101100;
      patterns[27827] = 29'b0_110110010110_011_1_011001011001;
      patterns[27828] = 29'b0_110110010110_100_0_011011001011;
      patterns[27829] = 29'b0_110110010110_101_1_001101100101;
      patterns[27830] = 29'b0_110110010110_110_0_110110010110;
      patterns[27831] = 29'b0_110110010110_111_0_110110010110;
      patterns[27832] = 29'b0_110110010111_000_0_110110010111;
      patterns[27833] = 29'b0_110110010111_001_0_010111110110;
      patterns[27834] = 29'b0_110110010111_010_1_101100101110;
      patterns[27835] = 29'b0_110110010111_011_1_011001011101;
      patterns[27836] = 29'b0_110110010111_100_1_011011001011;
      patterns[27837] = 29'b0_110110010111_101_1_101101100101;
      patterns[27838] = 29'b0_110110010111_110_0_110110010111;
      patterns[27839] = 29'b0_110110010111_111_0_110110010111;
      patterns[27840] = 29'b0_110110011000_000_0_110110011000;
      patterns[27841] = 29'b0_110110011000_001_0_011000110110;
      patterns[27842] = 29'b0_110110011000_010_1_101100110000;
      patterns[27843] = 29'b0_110110011000_011_1_011001100001;
      patterns[27844] = 29'b0_110110011000_100_0_011011001100;
      patterns[27845] = 29'b0_110110011000_101_0_001101100110;
      patterns[27846] = 29'b0_110110011000_110_0_110110011000;
      patterns[27847] = 29'b0_110110011000_111_0_110110011000;
      patterns[27848] = 29'b0_110110011001_000_0_110110011001;
      patterns[27849] = 29'b0_110110011001_001_0_011001110110;
      patterns[27850] = 29'b0_110110011001_010_1_101100110010;
      patterns[27851] = 29'b0_110110011001_011_1_011001100101;
      patterns[27852] = 29'b0_110110011001_100_1_011011001100;
      patterns[27853] = 29'b0_110110011001_101_0_101101100110;
      patterns[27854] = 29'b0_110110011001_110_0_110110011001;
      patterns[27855] = 29'b0_110110011001_111_0_110110011001;
      patterns[27856] = 29'b0_110110011010_000_0_110110011010;
      patterns[27857] = 29'b0_110110011010_001_0_011010110110;
      patterns[27858] = 29'b0_110110011010_010_1_101100110100;
      patterns[27859] = 29'b0_110110011010_011_1_011001101001;
      patterns[27860] = 29'b0_110110011010_100_0_011011001101;
      patterns[27861] = 29'b0_110110011010_101_1_001101100110;
      patterns[27862] = 29'b0_110110011010_110_0_110110011010;
      patterns[27863] = 29'b0_110110011010_111_0_110110011010;
      patterns[27864] = 29'b0_110110011011_000_0_110110011011;
      patterns[27865] = 29'b0_110110011011_001_0_011011110110;
      patterns[27866] = 29'b0_110110011011_010_1_101100110110;
      patterns[27867] = 29'b0_110110011011_011_1_011001101101;
      patterns[27868] = 29'b0_110110011011_100_1_011011001101;
      patterns[27869] = 29'b0_110110011011_101_1_101101100110;
      patterns[27870] = 29'b0_110110011011_110_0_110110011011;
      patterns[27871] = 29'b0_110110011011_111_0_110110011011;
      patterns[27872] = 29'b0_110110011100_000_0_110110011100;
      patterns[27873] = 29'b0_110110011100_001_0_011100110110;
      patterns[27874] = 29'b0_110110011100_010_1_101100111000;
      patterns[27875] = 29'b0_110110011100_011_1_011001110001;
      patterns[27876] = 29'b0_110110011100_100_0_011011001110;
      patterns[27877] = 29'b0_110110011100_101_0_001101100111;
      patterns[27878] = 29'b0_110110011100_110_0_110110011100;
      patterns[27879] = 29'b0_110110011100_111_0_110110011100;
      patterns[27880] = 29'b0_110110011101_000_0_110110011101;
      patterns[27881] = 29'b0_110110011101_001_0_011101110110;
      patterns[27882] = 29'b0_110110011101_010_1_101100111010;
      patterns[27883] = 29'b0_110110011101_011_1_011001110101;
      patterns[27884] = 29'b0_110110011101_100_1_011011001110;
      patterns[27885] = 29'b0_110110011101_101_0_101101100111;
      patterns[27886] = 29'b0_110110011101_110_0_110110011101;
      patterns[27887] = 29'b0_110110011101_111_0_110110011101;
      patterns[27888] = 29'b0_110110011110_000_0_110110011110;
      patterns[27889] = 29'b0_110110011110_001_0_011110110110;
      patterns[27890] = 29'b0_110110011110_010_1_101100111100;
      patterns[27891] = 29'b0_110110011110_011_1_011001111001;
      patterns[27892] = 29'b0_110110011110_100_0_011011001111;
      patterns[27893] = 29'b0_110110011110_101_1_001101100111;
      patterns[27894] = 29'b0_110110011110_110_0_110110011110;
      patterns[27895] = 29'b0_110110011110_111_0_110110011110;
      patterns[27896] = 29'b0_110110011111_000_0_110110011111;
      patterns[27897] = 29'b0_110110011111_001_0_011111110110;
      patterns[27898] = 29'b0_110110011111_010_1_101100111110;
      patterns[27899] = 29'b0_110110011111_011_1_011001111101;
      patterns[27900] = 29'b0_110110011111_100_1_011011001111;
      patterns[27901] = 29'b0_110110011111_101_1_101101100111;
      patterns[27902] = 29'b0_110110011111_110_0_110110011111;
      patterns[27903] = 29'b0_110110011111_111_0_110110011111;
      patterns[27904] = 29'b0_110110100000_000_0_110110100000;
      patterns[27905] = 29'b0_110110100000_001_0_100000110110;
      patterns[27906] = 29'b0_110110100000_010_1_101101000000;
      patterns[27907] = 29'b0_110110100000_011_1_011010000001;
      patterns[27908] = 29'b0_110110100000_100_0_011011010000;
      patterns[27909] = 29'b0_110110100000_101_0_001101101000;
      patterns[27910] = 29'b0_110110100000_110_0_110110100000;
      patterns[27911] = 29'b0_110110100000_111_0_110110100000;
      patterns[27912] = 29'b0_110110100001_000_0_110110100001;
      patterns[27913] = 29'b0_110110100001_001_0_100001110110;
      patterns[27914] = 29'b0_110110100001_010_1_101101000010;
      patterns[27915] = 29'b0_110110100001_011_1_011010000101;
      patterns[27916] = 29'b0_110110100001_100_1_011011010000;
      patterns[27917] = 29'b0_110110100001_101_0_101101101000;
      patterns[27918] = 29'b0_110110100001_110_0_110110100001;
      patterns[27919] = 29'b0_110110100001_111_0_110110100001;
      patterns[27920] = 29'b0_110110100010_000_0_110110100010;
      patterns[27921] = 29'b0_110110100010_001_0_100010110110;
      patterns[27922] = 29'b0_110110100010_010_1_101101000100;
      patterns[27923] = 29'b0_110110100010_011_1_011010001001;
      patterns[27924] = 29'b0_110110100010_100_0_011011010001;
      patterns[27925] = 29'b0_110110100010_101_1_001101101000;
      patterns[27926] = 29'b0_110110100010_110_0_110110100010;
      patterns[27927] = 29'b0_110110100010_111_0_110110100010;
      patterns[27928] = 29'b0_110110100011_000_0_110110100011;
      patterns[27929] = 29'b0_110110100011_001_0_100011110110;
      patterns[27930] = 29'b0_110110100011_010_1_101101000110;
      patterns[27931] = 29'b0_110110100011_011_1_011010001101;
      patterns[27932] = 29'b0_110110100011_100_1_011011010001;
      patterns[27933] = 29'b0_110110100011_101_1_101101101000;
      patterns[27934] = 29'b0_110110100011_110_0_110110100011;
      patterns[27935] = 29'b0_110110100011_111_0_110110100011;
      patterns[27936] = 29'b0_110110100100_000_0_110110100100;
      patterns[27937] = 29'b0_110110100100_001_0_100100110110;
      patterns[27938] = 29'b0_110110100100_010_1_101101001000;
      patterns[27939] = 29'b0_110110100100_011_1_011010010001;
      patterns[27940] = 29'b0_110110100100_100_0_011011010010;
      patterns[27941] = 29'b0_110110100100_101_0_001101101001;
      patterns[27942] = 29'b0_110110100100_110_0_110110100100;
      patterns[27943] = 29'b0_110110100100_111_0_110110100100;
      patterns[27944] = 29'b0_110110100101_000_0_110110100101;
      patterns[27945] = 29'b0_110110100101_001_0_100101110110;
      patterns[27946] = 29'b0_110110100101_010_1_101101001010;
      patterns[27947] = 29'b0_110110100101_011_1_011010010101;
      patterns[27948] = 29'b0_110110100101_100_1_011011010010;
      patterns[27949] = 29'b0_110110100101_101_0_101101101001;
      patterns[27950] = 29'b0_110110100101_110_0_110110100101;
      patterns[27951] = 29'b0_110110100101_111_0_110110100101;
      patterns[27952] = 29'b0_110110100110_000_0_110110100110;
      patterns[27953] = 29'b0_110110100110_001_0_100110110110;
      patterns[27954] = 29'b0_110110100110_010_1_101101001100;
      patterns[27955] = 29'b0_110110100110_011_1_011010011001;
      patterns[27956] = 29'b0_110110100110_100_0_011011010011;
      patterns[27957] = 29'b0_110110100110_101_1_001101101001;
      patterns[27958] = 29'b0_110110100110_110_0_110110100110;
      patterns[27959] = 29'b0_110110100110_111_0_110110100110;
      patterns[27960] = 29'b0_110110100111_000_0_110110100111;
      patterns[27961] = 29'b0_110110100111_001_0_100111110110;
      patterns[27962] = 29'b0_110110100111_010_1_101101001110;
      patterns[27963] = 29'b0_110110100111_011_1_011010011101;
      patterns[27964] = 29'b0_110110100111_100_1_011011010011;
      patterns[27965] = 29'b0_110110100111_101_1_101101101001;
      patterns[27966] = 29'b0_110110100111_110_0_110110100111;
      patterns[27967] = 29'b0_110110100111_111_0_110110100111;
      patterns[27968] = 29'b0_110110101000_000_0_110110101000;
      patterns[27969] = 29'b0_110110101000_001_0_101000110110;
      patterns[27970] = 29'b0_110110101000_010_1_101101010000;
      patterns[27971] = 29'b0_110110101000_011_1_011010100001;
      patterns[27972] = 29'b0_110110101000_100_0_011011010100;
      patterns[27973] = 29'b0_110110101000_101_0_001101101010;
      patterns[27974] = 29'b0_110110101000_110_0_110110101000;
      patterns[27975] = 29'b0_110110101000_111_0_110110101000;
      patterns[27976] = 29'b0_110110101001_000_0_110110101001;
      patterns[27977] = 29'b0_110110101001_001_0_101001110110;
      patterns[27978] = 29'b0_110110101001_010_1_101101010010;
      patterns[27979] = 29'b0_110110101001_011_1_011010100101;
      patterns[27980] = 29'b0_110110101001_100_1_011011010100;
      patterns[27981] = 29'b0_110110101001_101_0_101101101010;
      patterns[27982] = 29'b0_110110101001_110_0_110110101001;
      patterns[27983] = 29'b0_110110101001_111_0_110110101001;
      patterns[27984] = 29'b0_110110101010_000_0_110110101010;
      patterns[27985] = 29'b0_110110101010_001_0_101010110110;
      patterns[27986] = 29'b0_110110101010_010_1_101101010100;
      patterns[27987] = 29'b0_110110101010_011_1_011010101001;
      patterns[27988] = 29'b0_110110101010_100_0_011011010101;
      patterns[27989] = 29'b0_110110101010_101_1_001101101010;
      patterns[27990] = 29'b0_110110101010_110_0_110110101010;
      patterns[27991] = 29'b0_110110101010_111_0_110110101010;
      patterns[27992] = 29'b0_110110101011_000_0_110110101011;
      patterns[27993] = 29'b0_110110101011_001_0_101011110110;
      patterns[27994] = 29'b0_110110101011_010_1_101101010110;
      patterns[27995] = 29'b0_110110101011_011_1_011010101101;
      patterns[27996] = 29'b0_110110101011_100_1_011011010101;
      patterns[27997] = 29'b0_110110101011_101_1_101101101010;
      patterns[27998] = 29'b0_110110101011_110_0_110110101011;
      patterns[27999] = 29'b0_110110101011_111_0_110110101011;
      patterns[28000] = 29'b0_110110101100_000_0_110110101100;
      patterns[28001] = 29'b0_110110101100_001_0_101100110110;
      patterns[28002] = 29'b0_110110101100_010_1_101101011000;
      patterns[28003] = 29'b0_110110101100_011_1_011010110001;
      patterns[28004] = 29'b0_110110101100_100_0_011011010110;
      patterns[28005] = 29'b0_110110101100_101_0_001101101011;
      patterns[28006] = 29'b0_110110101100_110_0_110110101100;
      patterns[28007] = 29'b0_110110101100_111_0_110110101100;
      patterns[28008] = 29'b0_110110101101_000_0_110110101101;
      patterns[28009] = 29'b0_110110101101_001_0_101101110110;
      patterns[28010] = 29'b0_110110101101_010_1_101101011010;
      patterns[28011] = 29'b0_110110101101_011_1_011010110101;
      patterns[28012] = 29'b0_110110101101_100_1_011011010110;
      patterns[28013] = 29'b0_110110101101_101_0_101101101011;
      patterns[28014] = 29'b0_110110101101_110_0_110110101101;
      patterns[28015] = 29'b0_110110101101_111_0_110110101101;
      patterns[28016] = 29'b0_110110101110_000_0_110110101110;
      patterns[28017] = 29'b0_110110101110_001_0_101110110110;
      patterns[28018] = 29'b0_110110101110_010_1_101101011100;
      patterns[28019] = 29'b0_110110101110_011_1_011010111001;
      patterns[28020] = 29'b0_110110101110_100_0_011011010111;
      patterns[28021] = 29'b0_110110101110_101_1_001101101011;
      patterns[28022] = 29'b0_110110101110_110_0_110110101110;
      patterns[28023] = 29'b0_110110101110_111_0_110110101110;
      patterns[28024] = 29'b0_110110101111_000_0_110110101111;
      patterns[28025] = 29'b0_110110101111_001_0_101111110110;
      patterns[28026] = 29'b0_110110101111_010_1_101101011110;
      patterns[28027] = 29'b0_110110101111_011_1_011010111101;
      patterns[28028] = 29'b0_110110101111_100_1_011011010111;
      patterns[28029] = 29'b0_110110101111_101_1_101101101011;
      patterns[28030] = 29'b0_110110101111_110_0_110110101111;
      patterns[28031] = 29'b0_110110101111_111_0_110110101111;
      patterns[28032] = 29'b0_110110110000_000_0_110110110000;
      patterns[28033] = 29'b0_110110110000_001_0_110000110110;
      patterns[28034] = 29'b0_110110110000_010_1_101101100000;
      patterns[28035] = 29'b0_110110110000_011_1_011011000001;
      patterns[28036] = 29'b0_110110110000_100_0_011011011000;
      patterns[28037] = 29'b0_110110110000_101_0_001101101100;
      patterns[28038] = 29'b0_110110110000_110_0_110110110000;
      patterns[28039] = 29'b0_110110110000_111_0_110110110000;
      patterns[28040] = 29'b0_110110110001_000_0_110110110001;
      patterns[28041] = 29'b0_110110110001_001_0_110001110110;
      patterns[28042] = 29'b0_110110110001_010_1_101101100010;
      patterns[28043] = 29'b0_110110110001_011_1_011011000101;
      patterns[28044] = 29'b0_110110110001_100_1_011011011000;
      patterns[28045] = 29'b0_110110110001_101_0_101101101100;
      patterns[28046] = 29'b0_110110110001_110_0_110110110001;
      patterns[28047] = 29'b0_110110110001_111_0_110110110001;
      patterns[28048] = 29'b0_110110110010_000_0_110110110010;
      patterns[28049] = 29'b0_110110110010_001_0_110010110110;
      patterns[28050] = 29'b0_110110110010_010_1_101101100100;
      patterns[28051] = 29'b0_110110110010_011_1_011011001001;
      patterns[28052] = 29'b0_110110110010_100_0_011011011001;
      patterns[28053] = 29'b0_110110110010_101_1_001101101100;
      patterns[28054] = 29'b0_110110110010_110_0_110110110010;
      patterns[28055] = 29'b0_110110110010_111_0_110110110010;
      patterns[28056] = 29'b0_110110110011_000_0_110110110011;
      patterns[28057] = 29'b0_110110110011_001_0_110011110110;
      patterns[28058] = 29'b0_110110110011_010_1_101101100110;
      patterns[28059] = 29'b0_110110110011_011_1_011011001101;
      patterns[28060] = 29'b0_110110110011_100_1_011011011001;
      patterns[28061] = 29'b0_110110110011_101_1_101101101100;
      patterns[28062] = 29'b0_110110110011_110_0_110110110011;
      patterns[28063] = 29'b0_110110110011_111_0_110110110011;
      patterns[28064] = 29'b0_110110110100_000_0_110110110100;
      patterns[28065] = 29'b0_110110110100_001_0_110100110110;
      patterns[28066] = 29'b0_110110110100_010_1_101101101000;
      patterns[28067] = 29'b0_110110110100_011_1_011011010001;
      patterns[28068] = 29'b0_110110110100_100_0_011011011010;
      patterns[28069] = 29'b0_110110110100_101_0_001101101101;
      patterns[28070] = 29'b0_110110110100_110_0_110110110100;
      patterns[28071] = 29'b0_110110110100_111_0_110110110100;
      patterns[28072] = 29'b0_110110110101_000_0_110110110101;
      patterns[28073] = 29'b0_110110110101_001_0_110101110110;
      patterns[28074] = 29'b0_110110110101_010_1_101101101010;
      patterns[28075] = 29'b0_110110110101_011_1_011011010101;
      patterns[28076] = 29'b0_110110110101_100_1_011011011010;
      patterns[28077] = 29'b0_110110110101_101_0_101101101101;
      patterns[28078] = 29'b0_110110110101_110_0_110110110101;
      patterns[28079] = 29'b0_110110110101_111_0_110110110101;
      patterns[28080] = 29'b0_110110110110_000_0_110110110110;
      patterns[28081] = 29'b0_110110110110_001_0_110110110110;
      patterns[28082] = 29'b0_110110110110_010_1_101101101100;
      patterns[28083] = 29'b0_110110110110_011_1_011011011001;
      patterns[28084] = 29'b0_110110110110_100_0_011011011011;
      patterns[28085] = 29'b0_110110110110_101_1_001101101101;
      patterns[28086] = 29'b0_110110110110_110_0_110110110110;
      patterns[28087] = 29'b0_110110110110_111_0_110110110110;
      patterns[28088] = 29'b0_110110110111_000_0_110110110111;
      patterns[28089] = 29'b0_110110110111_001_0_110111110110;
      patterns[28090] = 29'b0_110110110111_010_1_101101101110;
      patterns[28091] = 29'b0_110110110111_011_1_011011011101;
      patterns[28092] = 29'b0_110110110111_100_1_011011011011;
      patterns[28093] = 29'b0_110110110111_101_1_101101101101;
      patterns[28094] = 29'b0_110110110111_110_0_110110110111;
      patterns[28095] = 29'b0_110110110111_111_0_110110110111;
      patterns[28096] = 29'b0_110110111000_000_0_110110111000;
      patterns[28097] = 29'b0_110110111000_001_0_111000110110;
      patterns[28098] = 29'b0_110110111000_010_1_101101110000;
      patterns[28099] = 29'b0_110110111000_011_1_011011100001;
      patterns[28100] = 29'b0_110110111000_100_0_011011011100;
      patterns[28101] = 29'b0_110110111000_101_0_001101101110;
      patterns[28102] = 29'b0_110110111000_110_0_110110111000;
      patterns[28103] = 29'b0_110110111000_111_0_110110111000;
      patterns[28104] = 29'b0_110110111001_000_0_110110111001;
      patterns[28105] = 29'b0_110110111001_001_0_111001110110;
      patterns[28106] = 29'b0_110110111001_010_1_101101110010;
      patterns[28107] = 29'b0_110110111001_011_1_011011100101;
      patterns[28108] = 29'b0_110110111001_100_1_011011011100;
      patterns[28109] = 29'b0_110110111001_101_0_101101101110;
      patterns[28110] = 29'b0_110110111001_110_0_110110111001;
      patterns[28111] = 29'b0_110110111001_111_0_110110111001;
      patterns[28112] = 29'b0_110110111010_000_0_110110111010;
      patterns[28113] = 29'b0_110110111010_001_0_111010110110;
      patterns[28114] = 29'b0_110110111010_010_1_101101110100;
      patterns[28115] = 29'b0_110110111010_011_1_011011101001;
      patterns[28116] = 29'b0_110110111010_100_0_011011011101;
      patterns[28117] = 29'b0_110110111010_101_1_001101101110;
      patterns[28118] = 29'b0_110110111010_110_0_110110111010;
      patterns[28119] = 29'b0_110110111010_111_0_110110111010;
      patterns[28120] = 29'b0_110110111011_000_0_110110111011;
      patterns[28121] = 29'b0_110110111011_001_0_111011110110;
      patterns[28122] = 29'b0_110110111011_010_1_101101110110;
      patterns[28123] = 29'b0_110110111011_011_1_011011101101;
      patterns[28124] = 29'b0_110110111011_100_1_011011011101;
      patterns[28125] = 29'b0_110110111011_101_1_101101101110;
      patterns[28126] = 29'b0_110110111011_110_0_110110111011;
      patterns[28127] = 29'b0_110110111011_111_0_110110111011;
      patterns[28128] = 29'b0_110110111100_000_0_110110111100;
      patterns[28129] = 29'b0_110110111100_001_0_111100110110;
      patterns[28130] = 29'b0_110110111100_010_1_101101111000;
      patterns[28131] = 29'b0_110110111100_011_1_011011110001;
      patterns[28132] = 29'b0_110110111100_100_0_011011011110;
      patterns[28133] = 29'b0_110110111100_101_0_001101101111;
      patterns[28134] = 29'b0_110110111100_110_0_110110111100;
      patterns[28135] = 29'b0_110110111100_111_0_110110111100;
      patterns[28136] = 29'b0_110110111101_000_0_110110111101;
      patterns[28137] = 29'b0_110110111101_001_0_111101110110;
      patterns[28138] = 29'b0_110110111101_010_1_101101111010;
      patterns[28139] = 29'b0_110110111101_011_1_011011110101;
      patterns[28140] = 29'b0_110110111101_100_1_011011011110;
      patterns[28141] = 29'b0_110110111101_101_0_101101101111;
      patterns[28142] = 29'b0_110110111101_110_0_110110111101;
      patterns[28143] = 29'b0_110110111101_111_0_110110111101;
      patterns[28144] = 29'b0_110110111110_000_0_110110111110;
      patterns[28145] = 29'b0_110110111110_001_0_111110110110;
      patterns[28146] = 29'b0_110110111110_010_1_101101111100;
      patterns[28147] = 29'b0_110110111110_011_1_011011111001;
      patterns[28148] = 29'b0_110110111110_100_0_011011011111;
      patterns[28149] = 29'b0_110110111110_101_1_001101101111;
      patterns[28150] = 29'b0_110110111110_110_0_110110111110;
      patterns[28151] = 29'b0_110110111110_111_0_110110111110;
      patterns[28152] = 29'b0_110110111111_000_0_110110111111;
      patterns[28153] = 29'b0_110110111111_001_0_111111110110;
      patterns[28154] = 29'b0_110110111111_010_1_101101111110;
      patterns[28155] = 29'b0_110110111111_011_1_011011111101;
      patterns[28156] = 29'b0_110110111111_100_1_011011011111;
      patterns[28157] = 29'b0_110110111111_101_1_101101101111;
      patterns[28158] = 29'b0_110110111111_110_0_110110111111;
      patterns[28159] = 29'b0_110110111111_111_0_110110111111;
      patterns[28160] = 29'b0_110111000000_000_0_110111000000;
      patterns[28161] = 29'b0_110111000000_001_0_000000110111;
      patterns[28162] = 29'b0_110111000000_010_1_101110000000;
      patterns[28163] = 29'b0_110111000000_011_1_011100000001;
      patterns[28164] = 29'b0_110111000000_100_0_011011100000;
      patterns[28165] = 29'b0_110111000000_101_0_001101110000;
      patterns[28166] = 29'b0_110111000000_110_0_110111000000;
      patterns[28167] = 29'b0_110111000000_111_0_110111000000;
      patterns[28168] = 29'b0_110111000001_000_0_110111000001;
      patterns[28169] = 29'b0_110111000001_001_0_000001110111;
      patterns[28170] = 29'b0_110111000001_010_1_101110000010;
      patterns[28171] = 29'b0_110111000001_011_1_011100000101;
      patterns[28172] = 29'b0_110111000001_100_1_011011100000;
      patterns[28173] = 29'b0_110111000001_101_0_101101110000;
      patterns[28174] = 29'b0_110111000001_110_0_110111000001;
      patterns[28175] = 29'b0_110111000001_111_0_110111000001;
      patterns[28176] = 29'b0_110111000010_000_0_110111000010;
      patterns[28177] = 29'b0_110111000010_001_0_000010110111;
      patterns[28178] = 29'b0_110111000010_010_1_101110000100;
      patterns[28179] = 29'b0_110111000010_011_1_011100001001;
      patterns[28180] = 29'b0_110111000010_100_0_011011100001;
      patterns[28181] = 29'b0_110111000010_101_1_001101110000;
      patterns[28182] = 29'b0_110111000010_110_0_110111000010;
      patterns[28183] = 29'b0_110111000010_111_0_110111000010;
      patterns[28184] = 29'b0_110111000011_000_0_110111000011;
      patterns[28185] = 29'b0_110111000011_001_0_000011110111;
      patterns[28186] = 29'b0_110111000011_010_1_101110000110;
      patterns[28187] = 29'b0_110111000011_011_1_011100001101;
      patterns[28188] = 29'b0_110111000011_100_1_011011100001;
      patterns[28189] = 29'b0_110111000011_101_1_101101110000;
      patterns[28190] = 29'b0_110111000011_110_0_110111000011;
      patterns[28191] = 29'b0_110111000011_111_0_110111000011;
      patterns[28192] = 29'b0_110111000100_000_0_110111000100;
      patterns[28193] = 29'b0_110111000100_001_0_000100110111;
      patterns[28194] = 29'b0_110111000100_010_1_101110001000;
      patterns[28195] = 29'b0_110111000100_011_1_011100010001;
      patterns[28196] = 29'b0_110111000100_100_0_011011100010;
      patterns[28197] = 29'b0_110111000100_101_0_001101110001;
      patterns[28198] = 29'b0_110111000100_110_0_110111000100;
      patterns[28199] = 29'b0_110111000100_111_0_110111000100;
      patterns[28200] = 29'b0_110111000101_000_0_110111000101;
      patterns[28201] = 29'b0_110111000101_001_0_000101110111;
      patterns[28202] = 29'b0_110111000101_010_1_101110001010;
      patterns[28203] = 29'b0_110111000101_011_1_011100010101;
      patterns[28204] = 29'b0_110111000101_100_1_011011100010;
      patterns[28205] = 29'b0_110111000101_101_0_101101110001;
      patterns[28206] = 29'b0_110111000101_110_0_110111000101;
      patterns[28207] = 29'b0_110111000101_111_0_110111000101;
      patterns[28208] = 29'b0_110111000110_000_0_110111000110;
      patterns[28209] = 29'b0_110111000110_001_0_000110110111;
      patterns[28210] = 29'b0_110111000110_010_1_101110001100;
      patterns[28211] = 29'b0_110111000110_011_1_011100011001;
      patterns[28212] = 29'b0_110111000110_100_0_011011100011;
      patterns[28213] = 29'b0_110111000110_101_1_001101110001;
      patterns[28214] = 29'b0_110111000110_110_0_110111000110;
      patterns[28215] = 29'b0_110111000110_111_0_110111000110;
      patterns[28216] = 29'b0_110111000111_000_0_110111000111;
      patterns[28217] = 29'b0_110111000111_001_0_000111110111;
      patterns[28218] = 29'b0_110111000111_010_1_101110001110;
      patterns[28219] = 29'b0_110111000111_011_1_011100011101;
      patterns[28220] = 29'b0_110111000111_100_1_011011100011;
      patterns[28221] = 29'b0_110111000111_101_1_101101110001;
      patterns[28222] = 29'b0_110111000111_110_0_110111000111;
      patterns[28223] = 29'b0_110111000111_111_0_110111000111;
      patterns[28224] = 29'b0_110111001000_000_0_110111001000;
      patterns[28225] = 29'b0_110111001000_001_0_001000110111;
      patterns[28226] = 29'b0_110111001000_010_1_101110010000;
      patterns[28227] = 29'b0_110111001000_011_1_011100100001;
      patterns[28228] = 29'b0_110111001000_100_0_011011100100;
      patterns[28229] = 29'b0_110111001000_101_0_001101110010;
      patterns[28230] = 29'b0_110111001000_110_0_110111001000;
      patterns[28231] = 29'b0_110111001000_111_0_110111001000;
      patterns[28232] = 29'b0_110111001001_000_0_110111001001;
      patterns[28233] = 29'b0_110111001001_001_0_001001110111;
      patterns[28234] = 29'b0_110111001001_010_1_101110010010;
      patterns[28235] = 29'b0_110111001001_011_1_011100100101;
      patterns[28236] = 29'b0_110111001001_100_1_011011100100;
      patterns[28237] = 29'b0_110111001001_101_0_101101110010;
      patterns[28238] = 29'b0_110111001001_110_0_110111001001;
      patterns[28239] = 29'b0_110111001001_111_0_110111001001;
      patterns[28240] = 29'b0_110111001010_000_0_110111001010;
      patterns[28241] = 29'b0_110111001010_001_0_001010110111;
      patterns[28242] = 29'b0_110111001010_010_1_101110010100;
      patterns[28243] = 29'b0_110111001010_011_1_011100101001;
      patterns[28244] = 29'b0_110111001010_100_0_011011100101;
      patterns[28245] = 29'b0_110111001010_101_1_001101110010;
      patterns[28246] = 29'b0_110111001010_110_0_110111001010;
      patterns[28247] = 29'b0_110111001010_111_0_110111001010;
      patterns[28248] = 29'b0_110111001011_000_0_110111001011;
      patterns[28249] = 29'b0_110111001011_001_0_001011110111;
      patterns[28250] = 29'b0_110111001011_010_1_101110010110;
      patterns[28251] = 29'b0_110111001011_011_1_011100101101;
      patterns[28252] = 29'b0_110111001011_100_1_011011100101;
      patterns[28253] = 29'b0_110111001011_101_1_101101110010;
      patterns[28254] = 29'b0_110111001011_110_0_110111001011;
      patterns[28255] = 29'b0_110111001011_111_0_110111001011;
      patterns[28256] = 29'b0_110111001100_000_0_110111001100;
      patterns[28257] = 29'b0_110111001100_001_0_001100110111;
      patterns[28258] = 29'b0_110111001100_010_1_101110011000;
      patterns[28259] = 29'b0_110111001100_011_1_011100110001;
      patterns[28260] = 29'b0_110111001100_100_0_011011100110;
      patterns[28261] = 29'b0_110111001100_101_0_001101110011;
      patterns[28262] = 29'b0_110111001100_110_0_110111001100;
      patterns[28263] = 29'b0_110111001100_111_0_110111001100;
      patterns[28264] = 29'b0_110111001101_000_0_110111001101;
      patterns[28265] = 29'b0_110111001101_001_0_001101110111;
      patterns[28266] = 29'b0_110111001101_010_1_101110011010;
      patterns[28267] = 29'b0_110111001101_011_1_011100110101;
      patterns[28268] = 29'b0_110111001101_100_1_011011100110;
      patterns[28269] = 29'b0_110111001101_101_0_101101110011;
      patterns[28270] = 29'b0_110111001101_110_0_110111001101;
      patterns[28271] = 29'b0_110111001101_111_0_110111001101;
      patterns[28272] = 29'b0_110111001110_000_0_110111001110;
      patterns[28273] = 29'b0_110111001110_001_0_001110110111;
      patterns[28274] = 29'b0_110111001110_010_1_101110011100;
      patterns[28275] = 29'b0_110111001110_011_1_011100111001;
      patterns[28276] = 29'b0_110111001110_100_0_011011100111;
      patterns[28277] = 29'b0_110111001110_101_1_001101110011;
      patterns[28278] = 29'b0_110111001110_110_0_110111001110;
      patterns[28279] = 29'b0_110111001110_111_0_110111001110;
      patterns[28280] = 29'b0_110111001111_000_0_110111001111;
      patterns[28281] = 29'b0_110111001111_001_0_001111110111;
      patterns[28282] = 29'b0_110111001111_010_1_101110011110;
      patterns[28283] = 29'b0_110111001111_011_1_011100111101;
      patterns[28284] = 29'b0_110111001111_100_1_011011100111;
      patterns[28285] = 29'b0_110111001111_101_1_101101110011;
      patterns[28286] = 29'b0_110111001111_110_0_110111001111;
      patterns[28287] = 29'b0_110111001111_111_0_110111001111;
      patterns[28288] = 29'b0_110111010000_000_0_110111010000;
      patterns[28289] = 29'b0_110111010000_001_0_010000110111;
      patterns[28290] = 29'b0_110111010000_010_1_101110100000;
      patterns[28291] = 29'b0_110111010000_011_1_011101000001;
      patterns[28292] = 29'b0_110111010000_100_0_011011101000;
      patterns[28293] = 29'b0_110111010000_101_0_001101110100;
      patterns[28294] = 29'b0_110111010000_110_0_110111010000;
      patterns[28295] = 29'b0_110111010000_111_0_110111010000;
      patterns[28296] = 29'b0_110111010001_000_0_110111010001;
      patterns[28297] = 29'b0_110111010001_001_0_010001110111;
      patterns[28298] = 29'b0_110111010001_010_1_101110100010;
      patterns[28299] = 29'b0_110111010001_011_1_011101000101;
      patterns[28300] = 29'b0_110111010001_100_1_011011101000;
      patterns[28301] = 29'b0_110111010001_101_0_101101110100;
      patterns[28302] = 29'b0_110111010001_110_0_110111010001;
      patterns[28303] = 29'b0_110111010001_111_0_110111010001;
      patterns[28304] = 29'b0_110111010010_000_0_110111010010;
      patterns[28305] = 29'b0_110111010010_001_0_010010110111;
      patterns[28306] = 29'b0_110111010010_010_1_101110100100;
      patterns[28307] = 29'b0_110111010010_011_1_011101001001;
      patterns[28308] = 29'b0_110111010010_100_0_011011101001;
      patterns[28309] = 29'b0_110111010010_101_1_001101110100;
      patterns[28310] = 29'b0_110111010010_110_0_110111010010;
      patterns[28311] = 29'b0_110111010010_111_0_110111010010;
      patterns[28312] = 29'b0_110111010011_000_0_110111010011;
      patterns[28313] = 29'b0_110111010011_001_0_010011110111;
      patterns[28314] = 29'b0_110111010011_010_1_101110100110;
      patterns[28315] = 29'b0_110111010011_011_1_011101001101;
      patterns[28316] = 29'b0_110111010011_100_1_011011101001;
      patterns[28317] = 29'b0_110111010011_101_1_101101110100;
      patterns[28318] = 29'b0_110111010011_110_0_110111010011;
      patterns[28319] = 29'b0_110111010011_111_0_110111010011;
      patterns[28320] = 29'b0_110111010100_000_0_110111010100;
      patterns[28321] = 29'b0_110111010100_001_0_010100110111;
      patterns[28322] = 29'b0_110111010100_010_1_101110101000;
      patterns[28323] = 29'b0_110111010100_011_1_011101010001;
      patterns[28324] = 29'b0_110111010100_100_0_011011101010;
      patterns[28325] = 29'b0_110111010100_101_0_001101110101;
      patterns[28326] = 29'b0_110111010100_110_0_110111010100;
      patterns[28327] = 29'b0_110111010100_111_0_110111010100;
      patterns[28328] = 29'b0_110111010101_000_0_110111010101;
      patterns[28329] = 29'b0_110111010101_001_0_010101110111;
      patterns[28330] = 29'b0_110111010101_010_1_101110101010;
      patterns[28331] = 29'b0_110111010101_011_1_011101010101;
      patterns[28332] = 29'b0_110111010101_100_1_011011101010;
      patterns[28333] = 29'b0_110111010101_101_0_101101110101;
      patterns[28334] = 29'b0_110111010101_110_0_110111010101;
      patterns[28335] = 29'b0_110111010101_111_0_110111010101;
      patterns[28336] = 29'b0_110111010110_000_0_110111010110;
      patterns[28337] = 29'b0_110111010110_001_0_010110110111;
      patterns[28338] = 29'b0_110111010110_010_1_101110101100;
      patterns[28339] = 29'b0_110111010110_011_1_011101011001;
      patterns[28340] = 29'b0_110111010110_100_0_011011101011;
      patterns[28341] = 29'b0_110111010110_101_1_001101110101;
      patterns[28342] = 29'b0_110111010110_110_0_110111010110;
      patterns[28343] = 29'b0_110111010110_111_0_110111010110;
      patterns[28344] = 29'b0_110111010111_000_0_110111010111;
      patterns[28345] = 29'b0_110111010111_001_0_010111110111;
      patterns[28346] = 29'b0_110111010111_010_1_101110101110;
      patterns[28347] = 29'b0_110111010111_011_1_011101011101;
      patterns[28348] = 29'b0_110111010111_100_1_011011101011;
      patterns[28349] = 29'b0_110111010111_101_1_101101110101;
      patterns[28350] = 29'b0_110111010111_110_0_110111010111;
      patterns[28351] = 29'b0_110111010111_111_0_110111010111;
      patterns[28352] = 29'b0_110111011000_000_0_110111011000;
      patterns[28353] = 29'b0_110111011000_001_0_011000110111;
      patterns[28354] = 29'b0_110111011000_010_1_101110110000;
      patterns[28355] = 29'b0_110111011000_011_1_011101100001;
      patterns[28356] = 29'b0_110111011000_100_0_011011101100;
      patterns[28357] = 29'b0_110111011000_101_0_001101110110;
      patterns[28358] = 29'b0_110111011000_110_0_110111011000;
      patterns[28359] = 29'b0_110111011000_111_0_110111011000;
      patterns[28360] = 29'b0_110111011001_000_0_110111011001;
      patterns[28361] = 29'b0_110111011001_001_0_011001110111;
      patterns[28362] = 29'b0_110111011001_010_1_101110110010;
      patterns[28363] = 29'b0_110111011001_011_1_011101100101;
      patterns[28364] = 29'b0_110111011001_100_1_011011101100;
      patterns[28365] = 29'b0_110111011001_101_0_101101110110;
      patterns[28366] = 29'b0_110111011001_110_0_110111011001;
      patterns[28367] = 29'b0_110111011001_111_0_110111011001;
      patterns[28368] = 29'b0_110111011010_000_0_110111011010;
      patterns[28369] = 29'b0_110111011010_001_0_011010110111;
      patterns[28370] = 29'b0_110111011010_010_1_101110110100;
      patterns[28371] = 29'b0_110111011010_011_1_011101101001;
      patterns[28372] = 29'b0_110111011010_100_0_011011101101;
      patterns[28373] = 29'b0_110111011010_101_1_001101110110;
      patterns[28374] = 29'b0_110111011010_110_0_110111011010;
      patterns[28375] = 29'b0_110111011010_111_0_110111011010;
      patterns[28376] = 29'b0_110111011011_000_0_110111011011;
      patterns[28377] = 29'b0_110111011011_001_0_011011110111;
      patterns[28378] = 29'b0_110111011011_010_1_101110110110;
      patterns[28379] = 29'b0_110111011011_011_1_011101101101;
      patterns[28380] = 29'b0_110111011011_100_1_011011101101;
      patterns[28381] = 29'b0_110111011011_101_1_101101110110;
      patterns[28382] = 29'b0_110111011011_110_0_110111011011;
      patterns[28383] = 29'b0_110111011011_111_0_110111011011;
      patterns[28384] = 29'b0_110111011100_000_0_110111011100;
      patterns[28385] = 29'b0_110111011100_001_0_011100110111;
      patterns[28386] = 29'b0_110111011100_010_1_101110111000;
      patterns[28387] = 29'b0_110111011100_011_1_011101110001;
      patterns[28388] = 29'b0_110111011100_100_0_011011101110;
      patterns[28389] = 29'b0_110111011100_101_0_001101110111;
      patterns[28390] = 29'b0_110111011100_110_0_110111011100;
      patterns[28391] = 29'b0_110111011100_111_0_110111011100;
      patterns[28392] = 29'b0_110111011101_000_0_110111011101;
      patterns[28393] = 29'b0_110111011101_001_0_011101110111;
      patterns[28394] = 29'b0_110111011101_010_1_101110111010;
      patterns[28395] = 29'b0_110111011101_011_1_011101110101;
      patterns[28396] = 29'b0_110111011101_100_1_011011101110;
      patterns[28397] = 29'b0_110111011101_101_0_101101110111;
      patterns[28398] = 29'b0_110111011101_110_0_110111011101;
      patterns[28399] = 29'b0_110111011101_111_0_110111011101;
      patterns[28400] = 29'b0_110111011110_000_0_110111011110;
      patterns[28401] = 29'b0_110111011110_001_0_011110110111;
      patterns[28402] = 29'b0_110111011110_010_1_101110111100;
      patterns[28403] = 29'b0_110111011110_011_1_011101111001;
      patterns[28404] = 29'b0_110111011110_100_0_011011101111;
      patterns[28405] = 29'b0_110111011110_101_1_001101110111;
      patterns[28406] = 29'b0_110111011110_110_0_110111011110;
      patterns[28407] = 29'b0_110111011110_111_0_110111011110;
      patterns[28408] = 29'b0_110111011111_000_0_110111011111;
      patterns[28409] = 29'b0_110111011111_001_0_011111110111;
      patterns[28410] = 29'b0_110111011111_010_1_101110111110;
      patterns[28411] = 29'b0_110111011111_011_1_011101111101;
      patterns[28412] = 29'b0_110111011111_100_1_011011101111;
      patterns[28413] = 29'b0_110111011111_101_1_101101110111;
      patterns[28414] = 29'b0_110111011111_110_0_110111011111;
      patterns[28415] = 29'b0_110111011111_111_0_110111011111;
      patterns[28416] = 29'b0_110111100000_000_0_110111100000;
      patterns[28417] = 29'b0_110111100000_001_0_100000110111;
      patterns[28418] = 29'b0_110111100000_010_1_101111000000;
      patterns[28419] = 29'b0_110111100000_011_1_011110000001;
      patterns[28420] = 29'b0_110111100000_100_0_011011110000;
      patterns[28421] = 29'b0_110111100000_101_0_001101111000;
      patterns[28422] = 29'b0_110111100000_110_0_110111100000;
      patterns[28423] = 29'b0_110111100000_111_0_110111100000;
      patterns[28424] = 29'b0_110111100001_000_0_110111100001;
      patterns[28425] = 29'b0_110111100001_001_0_100001110111;
      patterns[28426] = 29'b0_110111100001_010_1_101111000010;
      patterns[28427] = 29'b0_110111100001_011_1_011110000101;
      patterns[28428] = 29'b0_110111100001_100_1_011011110000;
      patterns[28429] = 29'b0_110111100001_101_0_101101111000;
      patterns[28430] = 29'b0_110111100001_110_0_110111100001;
      patterns[28431] = 29'b0_110111100001_111_0_110111100001;
      patterns[28432] = 29'b0_110111100010_000_0_110111100010;
      patterns[28433] = 29'b0_110111100010_001_0_100010110111;
      patterns[28434] = 29'b0_110111100010_010_1_101111000100;
      patterns[28435] = 29'b0_110111100010_011_1_011110001001;
      patterns[28436] = 29'b0_110111100010_100_0_011011110001;
      patterns[28437] = 29'b0_110111100010_101_1_001101111000;
      patterns[28438] = 29'b0_110111100010_110_0_110111100010;
      patterns[28439] = 29'b0_110111100010_111_0_110111100010;
      patterns[28440] = 29'b0_110111100011_000_0_110111100011;
      patterns[28441] = 29'b0_110111100011_001_0_100011110111;
      patterns[28442] = 29'b0_110111100011_010_1_101111000110;
      patterns[28443] = 29'b0_110111100011_011_1_011110001101;
      patterns[28444] = 29'b0_110111100011_100_1_011011110001;
      patterns[28445] = 29'b0_110111100011_101_1_101101111000;
      patterns[28446] = 29'b0_110111100011_110_0_110111100011;
      patterns[28447] = 29'b0_110111100011_111_0_110111100011;
      patterns[28448] = 29'b0_110111100100_000_0_110111100100;
      patterns[28449] = 29'b0_110111100100_001_0_100100110111;
      patterns[28450] = 29'b0_110111100100_010_1_101111001000;
      patterns[28451] = 29'b0_110111100100_011_1_011110010001;
      patterns[28452] = 29'b0_110111100100_100_0_011011110010;
      patterns[28453] = 29'b0_110111100100_101_0_001101111001;
      patterns[28454] = 29'b0_110111100100_110_0_110111100100;
      patterns[28455] = 29'b0_110111100100_111_0_110111100100;
      patterns[28456] = 29'b0_110111100101_000_0_110111100101;
      patterns[28457] = 29'b0_110111100101_001_0_100101110111;
      patterns[28458] = 29'b0_110111100101_010_1_101111001010;
      patterns[28459] = 29'b0_110111100101_011_1_011110010101;
      patterns[28460] = 29'b0_110111100101_100_1_011011110010;
      patterns[28461] = 29'b0_110111100101_101_0_101101111001;
      patterns[28462] = 29'b0_110111100101_110_0_110111100101;
      patterns[28463] = 29'b0_110111100101_111_0_110111100101;
      patterns[28464] = 29'b0_110111100110_000_0_110111100110;
      patterns[28465] = 29'b0_110111100110_001_0_100110110111;
      patterns[28466] = 29'b0_110111100110_010_1_101111001100;
      patterns[28467] = 29'b0_110111100110_011_1_011110011001;
      patterns[28468] = 29'b0_110111100110_100_0_011011110011;
      patterns[28469] = 29'b0_110111100110_101_1_001101111001;
      patterns[28470] = 29'b0_110111100110_110_0_110111100110;
      patterns[28471] = 29'b0_110111100110_111_0_110111100110;
      patterns[28472] = 29'b0_110111100111_000_0_110111100111;
      patterns[28473] = 29'b0_110111100111_001_0_100111110111;
      patterns[28474] = 29'b0_110111100111_010_1_101111001110;
      patterns[28475] = 29'b0_110111100111_011_1_011110011101;
      patterns[28476] = 29'b0_110111100111_100_1_011011110011;
      patterns[28477] = 29'b0_110111100111_101_1_101101111001;
      patterns[28478] = 29'b0_110111100111_110_0_110111100111;
      patterns[28479] = 29'b0_110111100111_111_0_110111100111;
      patterns[28480] = 29'b0_110111101000_000_0_110111101000;
      patterns[28481] = 29'b0_110111101000_001_0_101000110111;
      patterns[28482] = 29'b0_110111101000_010_1_101111010000;
      patterns[28483] = 29'b0_110111101000_011_1_011110100001;
      patterns[28484] = 29'b0_110111101000_100_0_011011110100;
      patterns[28485] = 29'b0_110111101000_101_0_001101111010;
      patterns[28486] = 29'b0_110111101000_110_0_110111101000;
      patterns[28487] = 29'b0_110111101000_111_0_110111101000;
      patterns[28488] = 29'b0_110111101001_000_0_110111101001;
      patterns[28489] = 29'b0_110111101001_001_0_101001110111;
      patterns[28490] = 29'b0_110111101001_010_1_101111010010;
      patterns[28491] = 29'b0_110111101001_011_1_011110100101;
      patterns[28492] = 29'b0_110111101001_100_1_011011110100;
      patterns[28493] = 29'b0_110111101001_101_0_101101111010;
      patterns[28494] = 29'b0_110111101001_110_0_110111101001;
      patterns[28495] = 29'b0_110111101001_111_0_110111101001;
      patterns[28496] = 29'b0_110111101010_000_0_110111101010;
      patterns[28497] = 29'b0_110111101010_001_0_101010110111;
      patterns[28498] = 29'b0_110111101010_010_1_101111010100;
      patterns[28499] = 29'b0_110111101010_011_1_011110101001;
      patterns[28500] = 29'b0_110111101010_100_0_011011110101;
      patterns[28501] = 29'b0_110111101010_101_1_001101111010;
      patterns[28502] = 29'b0_110111101010_110_0_110111101010;
      patterns[28503] = 29'b0_110111101010_111_0_110111101010;
      patterns[28504] = 29'b0_110111101011_000_0_110111101011;
      patterns[28505] = 29'b0_110111101011_001_0_101011110111;
      patterns[28506] = 29'b0_110111101011_010_1_101111010110;
      patterns[28507] = 29'b0_110111101011_011_1_011110101101;
      patterns[28508] = 29'b0_110111101011_100_1_011011110101;
      patterns[28509] = 29'b0_110111101011_101_1_101101111010;
      patterns[28510] = 29'b0_110111101011_110_0_110111101011;
      patterns[28511] = 29'b0_110111101011_111_0_110111101011;
      patterns[28512] = 29'b0_110111101100_000_0_110111101100;
      patterns[28513] = 29'b0_110111101100_001_0_101100110111;
      patterns[28514] = 29'b0_110111101100_010_1_101111011000;
      patterns[28515] = 29'b0_110111101100_011_1_011110110001;
      patterns[28516] = 29'b0_110111101100_100_0_011011110110;
      patterns[28517] = 29'b0_110111101100_101_0_001101111011;
      patterns[28518] = 29'b0_110111101100_110_0_110111101100;
      patterns[28519] = 29'b0_110111101100_111_0_110111101100;
      patterns[28520] = 29'b0_110111101101_000_0_110111101101;
      patterns[28521] = 29'b0_110111101101_001_0_101101110111;
      patterns[28522] = 29'b0_110111101101_010_1_101111011010;
      patterns[28523] = 29'b0_110111101101_011_1_011110110101;
      patterns[28524] = 29'b0_110111101101_100_1_011011110110;
      patterns[28525] = 29'b0_110111101101_101_0_101101111011;
      patterns[28526] = 29'b0_110111101101_110_0_110111101101;
      patterns[28527] = 29'b0_110111101101_111_0_110111101101;
      patterns[28528] = 29'b0_110111101110_000_0_110111101110;
      patterns[28529] = 29'b0_110111101110_001_0_101110110111;
      patterns[28530] = 29'b0_110111101110_010_1_101111011100;
      patterns[28531] = 29'b0_110111101110_011_1_011110111001;
      patterns[28532] = 29'b0_110111101110_100_0_011011110111;
      patterns[28533] = 29'b0_110111101110_101_1_001101111011;
      patterns[28534] = 29'b0_110111101110_110_0_110111101110;
      patterns[28535] = 29'b0_110111101110_111_0_110111101110;
      patterns[28536] = 29'b0_110111101111_000_0_110111101111;
      patterns[28537] = 29'b0_110111101111_001_0_101111110111;
      patterns[28538] = 29'b0_110111101111_010_1_101111011110;
      patterns[28539] = 29'b0_110111101111_011_1_011110111101;
      patterns[28540] = 29'b0_110111101111_100_1_011011110111;
      patterns[28541] = 29'b0_110111101111_101_1_101101111011;
      patterns[28542] = 29'b0_110111101111_110_0_110111101111;
      patterns[28543] = 29'b0_110111101111_111_0_110111101111;
      patterns[28544] = 29'b0_110111110000_000_0_110111110000;
      patterns[28545] = 29'b0_110111110000_001_0_110000110111;
      patterns[28546] = 29'b0_110111110000_010_1_101111100000;
      patterns[28547] = 29'b0_110111110000_011_1_011111000001;
      patterns[28548] = 29'b0_110111110000_100_0_011011111000;
      patterns[28549] = 29'b0_110111110000_101_0_001101111100;
      patterns[28550] = 29'b0_110111110000_110_0_110111110000;
      patterns[28551] = 29'b0_110111110000_111_0_110111110000;
      patterns[28552] = 29'b0_110111110001_000_0_110111110001;
      patterns[28553] = 29'b0_110111110001_001_0_110001110111;
      patterns[28554] = 29'b0_110111110001_010_1_101111100010;
      patterns[28555] = 29'b0_110111110001_011_1_011111000101;
      patterns[28556] = 29'b0_110111110001_100_1_011011111000;
      patterns[28557] = 29'b0_110111110001_101_0_101101111100;
      patterns[28558] = 29'b0_110111110001_110_0_110111110001;
      patterns[28559] = 29'b0_110111110001_111_0_110111110001;
      patterns[28560] = 29'b0_110111110010_000_0_110111110010;
      patterns[28561] = 29'b0_110111110010_001_0_110010110111;
      patterns[28562] = 29'b0_110111110010_010_1_101111100100;
      patterns[28563] = 29'b0_110111110010_011_1_011111001001;
      patterns[28564] = 29'b0_110111110010_100_0_011011111001;
      patterns[28565] = 29'b0_110111110010_101_1_001101111100;
      patterns[28566] = 29'b0_110111110010_110_0_110111110010;
      patterns[28567] = 29'b0_110111110010_111_0_110111110010;
      patterns[28568] = 29'b0_110111110011_000_0_110111110011;
      patterns[28569] = 29'b0_110111110011_001_0_110011110111;
      patterns[28570] = 29'b0_110111110011_010_1_101111100110;
      patterns[28571] = 29'b0_110111110011_011_1_011111001101;
      patterns[28572] = 29'b0_110111110011_100_1_011011111001;
      patterns[28573] = 29'b0_110111110011_101_1_101101111100;
      patterns[28574] = 29'b0_110111110011_110_0_110111110011;
      patterns[28575] = 29'b0_110111110011_111_0_110111110011;
      patterns[28576] = 29'b0_110111110100_000_0_110111110100;
      patterns[28577] = 29'b0_110111110100_001_0_110100110111;
      patterns[28578] = 29'b0_110111110100_010_1_101111101000;
      patterns[28579] = 29'b0_110111110100_011_1_011111010001;
      patterns[28580] = 29'b0_110111110100_100_0_011011111010;
      patterns[28581] = 29'b0_110111110100_101_0_001101111101;
      patterns[28582] = 29'b0_110111110100_110_0_110111110100;
      patterns[28583] = 29'b0_110111110100_111_0_110111110100;
      patterns[28584] = 29'b0_110111110101_000_0_110111110101;
      patterns[28585] = 29'b0_110111110101_001_0_110101110111;
      patterns[28586] = 29'b0_110111110101_010_1_101111101010;
      patterns[28587] = 29'b0_110111110101_011_1_011111010101;
      patterns[28588] = 29'b0_110111110101_100_1_011011111010;
      patterns[28589] = 29'b0_110111110101_101_0_101101111101;
      patterns[28590] = 29'b0_110111110101_110_0_110111110101;
      patterns[28591] = 29'b0_110111110101_111_0_110111110101;
      patterns[28592] = 29'b0_110111110110_000_0_110111110110;
      patterns[28593] = 29'b0_110111110110_001_0_110110110111;
      patterns[28594] = 29'b0_110111110110_010_1_101111101100;
      patterns[28595] = 29'b0_110111110110_011_1_011111011001;
      patterns[28596] = 29'b0_110111110110_100_0_011011111011;
      patterns[28597] = 29'b0_110111110110_101_1_001101111101;
      patterns[28598] = 29'b0_110111110110_110_0_110111110110;
      patterns[28599] = 29'b0_110111110110_111_0_110111110110;
      patterns[28600] = 29'b0_110111110111_000_0_110111110111;
      patterns[28601] = 29'b0_110111110111_001_0_110111110111;
      patterns[28602] = 29'b0_110111110111_010_1_101111101110;
      patterns[28603] = 29'b0_110111110111_011_1_011111011101;
      patterns[28604] = 29'b0_110111110111_100_1_011011111011;
      patterns[28605] = 29'b0_110111110111_101_1_101101111101;
      patterns[28606] = 29'b0_110111110111_110_0_110111110111;
      patterns[28607] = 29'b0_110111110111_111_0_110111110111;
      patterns[28608] = 29'b0_110111111000_000_0_110111111000;
      patterns[28609] = 29'b0_110111111000_001_0_111000110111;
      patterns[28610] = 29'b0_110111111000_010_1_101111110000;
      patterns[28611] = 29'b0_110111111000_011_1_011111100001;
      patterns[28612] = 29'b0_110111111000_100_0_011011111100;
      patterns[28613] = 29'b0_110111111000_101_0_001101111110;
      patterns[28614] = 29'b0_110111111000_110_0_110111111000;
      patterns[28615] = 29'b0_110111111000_111_0_110111111000;
      patterns[28616] = 29'b0_110111111001_000_0_110111111001;
      patterns[28617] = 29'b0_110111111001_001_0_111001110111;
      patterns[28618] = 29'b0_110111111001_010_1_101111110010;
      patterns[28619] = 29'b0_110111111001_011_1_011111100101;
      patterns[28620] = 29'b0_110111111001_100_1_011011111100;
      patterns[28621] = 29'b0_110111111001_101_0_101101111110;
      patterns[28622] = 29'b0_110111111001_110_0_110111111001;
      patterns[28623] = 29'b0_110111111001_111_0_110111111001;
      patterns[28624] = 29'b0_110111111010_000_0_110111111010;
      patterns[28625] = 29'b0_110111111010_001_0_111010110111;
      patterns[28626] = 29'b0_110111111010_010_1_101111110100;
      patterns[28627] = 29'b0_110111111010_011_1_011111101001;
      patterns[28628] = 29'b0_110111111010_100_0_011011111101;
      patterns[28629] = 29'b0_110111111010_101_1_001101111110;
      patterns[28630] = 29'b0_110111111010_110_0_110111111010;
      patterns[28631] = 29'b0_110111111010_111_0_110111111010;
      patterns[28632] = 29'b0_110111111011_000_0_110111111011;
      patterns[28633] = 29'b0_110111111011_001_0_111011110111;
      patterns[28634] = 29'b0_110111111011_010_1_101111110110;
      patterns[28635] = 29'b0_110111111011_011_1_011111101101;
      patterns[28636] = 29'b0_110111111011_100_1_011011111101;
      patterns[28637] = 29'b0_110111111011_101_1_101101111110;
      patterns[28638] = 29'b0_110111111011_110_0_110111111011;
      patterns[28639] = 29'b0_110111111011_111_0_110111111011;
      patterns[28640] = 29'b0_110111111100_000_0_110111111100;
      patterns[28641] = 29'b0_110111111100_001_0_111100110111;
      patterns[28642] = 29'b0_110111111100_010_1_101111111000;
      patterns[28643] = 29'b0_110111111100_011_1_011111110001;
      patterns[28644] = 29'b0_110111111100_100_0_011011111110;
      patterns[28645] = 29'b0_110111111100_101_0_001101111111;
      patterns[28646] = 29'b0_110111111100_110_0_110111111100;
      patterns[28647] = 29'b0_110111111100_111_0_110111111100;
      patterns[28648] = 29'b0_110111111101_000_0_110111111101;
      patterns[28649] = 29'b0_110111111101_001_0_111101110111;
      patterns[28650] = 29'b0_110111111101_010_1_101111111010;
      patterns[28651] = 29'b0_110111111101_011_1_011111110101;
      patterns[28652] = 29'b0_110111111101_100_1_011011111110;
      patterns[28653] = 29'b0_110111111101_101_0_101101111111;
      patterns[28654] = 29'b0_110111111101_110_0_110111111101;
      patterns[28655] = 29'b0_110111111101_111_0_110111111101;
      patterns[28656] = 29'b0_110111111110_000_0_110111111110;
      patterns[28657] = 29'b0_110111111110_001_0_111110110111;
      patterns[28658] = 29'b0_110111111110_010_1_101111111100;
      patterns[28659] = 29'b0_110111111110_011_1_011111111001;
      patterns[28660] = 29'b0_110111111110_100_0_011011111111;
      patterns[28661] = 29'b0_110111111110_101_1_001101111111;
      patterns[28662] = 29'b0_110111111110_110_0_110111111110;
      patterns[28663] = 29'b0_110111111110_111_0_110111111110;
      patterns[28664] = 29'b0_110111111111_000_0_110111111111;
      patterns[28665] = 29'b0_110111111111_001_0_111111110111;
      patterns[28666] = 29'b0_110111111111_010_1_101111111110;
      patterns[28667] = 29'b0_110111111111_011_1_011111111101;
      patterns[28668] = 29'b0_110111111111_100_1_011011111111;
      patterns[28669] = 29'b0_110111111111_101_1_101101111111;
      patterns[28670] = 29'b0_110111111111_110_0_110111111111;
      patterns[28671] = 29'b0_110111111111_111_0_110111111111;
      patterns[28672] = 29'b0_111000000000_000_0_111000000000;
      patterns[28673] = 29'b0_111000000000_001_0_000000111000;
      patterns[28674] = 29'b0_111000000000_010_1_110000000000;
      patterns[28675] = 29'b0_111000000000_011_1_100000000001;
      patterns[28676] = 29'b0_111000000000_100_0_011100000000;
      patterns[28677] = 29'b0_111000000000_101_0_001110000000;
      patterns[28678] = 29'b0_111000000000_110_0_111000000000;
      patterns[28679] = 29'b0_111000000000_111_0_111000000000;
      patterns[28680] = 29'b0_111000000001_000_0_111000000001;
      patterns[28681] = 29'b0_111000000001_001_0_000001111000;
      patterns[28682] = 29'b0_111000000001_010_1_110000000010;
      patterns[28683] = 29'b0_111000000001_011_1_100000000101;
      patterns[28684] = 29'b0_111000000001_100_1_011100000000;
      patterns[28685] = 29'b0_111000000001_101_0_101110000000;
      patterns[28686] = 29'b0_111000000001_110_0_111000000001;
      patterns[28687] = 29'b0_111000000001_111_0_111000000001;
      patterns[28688] = 29'b0_111000000010_000_0_111000000010;
      patterns[28689] = 29'b0_111000000010_001_0_000010111000;
      patterns[28690] = 29'b0_111000000010_010_1_110000000100;
      patterns[28691] = 29'b0_111000000010_011_1_100000001001;
      patterns[28692] = 29'b0_111000000010_100_0_011100000001;
      patterns[28693] = 29'b0_111000000010_101_1_001110000000;
      patterns[28694] = 29'b0_111000000010_110_0_111000000010;
      patterns[28695] = 29'b0_111000000010_111_0_111000000010;
      patterns[28696] = 29'b0_111000000011_000_0_111000000011;
      patterns[28697] = 29'b0_111000000011_001_0_000011111000;
      patterns[28698] = 29'b0_111000000011_010_1_110000000110;
      patterns[28699] = 29'b0_111000000011_011_1_100000001101;
      patterns[28700] = 29'b0_111000000011_100_1_011100000001;
      patterns[28701] = 29'b0_111000000011_101_1_101110000000;
      patterns[28702] = 29'b0_111000000011_110_0_111000000011;
      patterns[28703] = 29'b0_111000000011_111_0_111000000011;
      patterns[28704] = 29'b0_111000000100_000_0_111000000100;
      patterns[28705] = 29'b0_111000000100_001_0_000100111000;
      patterns[28706] = 29'b0_111000000100_010_1_110000001000;
      patterns[28707] = 29'b0_111000000100_011_1_100000010001;
      patterns[28708] = 29'b0_111000000100_100_0_011100000010;
      patterns[28709] = 29'b0_111000000100_101_0_001110000001;
      patterns[28710] = 29'b0_111000000100_110_0_111000000100;
      patterns[28711] = 29'b0_111000000100_111_0_111000000100;
      patterns[28712] = 29'b0_111000000101_000_0_111000000101;
      patterns[28713] = 29'b0_111000000101_001_0_000101111000;
      patterns[28714] = 29'b0_111000000101_010_1_110000001010;
      patterns[28715] = 29'b0_111000000101_011_1_100000010101;
      patterns[28716] = 29'b0_111000000101_100_1_011100000010;
      patterns[28717] = 29'b0_111000000101_101_0_101110000001;
      patterns[28718] = 29'b0_111000000101_110_0_111000000101;
      patterns[28719] = 29'b0_111000000101_111_0_111000000101;
      patterns[28720] = 29'b0_111000000110_000_0_111000000110;
      patterns[28721] = 29'b0_111000000110_001_0_000110111000;
      patterns[28722] = 29'b0_111000000110_010_1_110000001100;
      patterns[28723] = 29'b0_111000000110_011_1_100000011001;
      patterns[28724] = 29'b0_111000000110_100_0_011100000011;
      patterns[28725] = 29'b0_111000000110_101_1_001110000001;
      patterns[28726] = 29'b0_111000000110_110_0_111000000110;
      patterns[28727] = 29'b0_111000000110_111_0_111000000110;
      patterns[28728] = 29'b0_111000000111_000_0_111000000111;
      patterns[28729] = 29'b0_111000000111_001_0_000111111000;
      patterns[28730] = 29'b0_111000000111_010_1_110000001110;
      patterns[28731] = 29'b0_111000000111_011_1_100000011101;
      patterns[28732] = 29'b0_111000000111_100_1_011100000011;
      patterns[28733] = 29'b0_111000000111_101_1_101110000001;
      patterns[28734] = 29'b0_111000000111_110_0_111000000111;
      patterns[28735] = 29'b0_111000000111_111_0_111000000111;
      patterns[28736] = 29'b0_111000001000_000_0_111000001000;
      patterns[28737] = 29'b0_111000001000_001_0_001000111000;
      patterns[28738] = 29'b0_111000001000_010_1_110000010000;
      patterns[28739] = 29'b0_111000001000_011_1_100000100001;
      patterns[28740] = 29'b0_111000001000_100_0_011100000100;
      patterns[28741] = 29'b0_111000001000_101_0_001110000010;
      patterns[28742] = 29'b0_111000001000_110_0_111000001000;
      patterns[28743] = 29'b0_111000001000_111_0_111000001000;
      patterns[28744] = 29'b0_111000001001_000_0_111000001001;
      patterns[28745] = 29'b0_111000001001_001_0_001001111000;
      patterns[28746] = 29'b0_111000001001_010_1_110000010010;
      patterns[28747] = 29'b0_111000001001_011_1_100000100101;
      patterns[28748] = 29'b0_111000001001_100_1_011100000100;
      patterns[28749] = 29'b0_111000001001_101_0_101110000010;
      patterns[28750] = 29'b0_111000001001_110_0_111000001001;
      patterns[28751] = 29'b0_111000001001_111_0_111000001001;
      patterns[28752] = 29'b0_111000001010_000_0_111000001010;
      patterns[28753] = 29'b0_111000001010_001_0_001010111000;
      patterns[28754] = 29'b0_111000001010_010_1_110000010100;
      patterns[28755] = 29'b0_111000001010_011_1_100000101001;
      patterns[28756] = 29'b0_111000001010_100_0_011100000101;
      patterns[28757] = 29'b0_111000001010_101_1_001110000010;
      patterns[28758] = 29'b0_111000001010_110_0_111000001010;
      patterns[28759] = 29'b0_111000001010_111_0_111000001010;
      patterns[28760] = 29'b0_111000001011_000_0_111000001011;
      patterns[28761] = 29'b0_111000001011_001_0_001011111000;
      patterns[28762] = 29'b0_111000001011_010_1_110000010110;
      patterns[28763] = 29'b0_111000001011_011_1_100000101101;
      patterns[28764] = 29'b0_111000001011_100_1_011100000101;
      patterns[28765] = 29'b0_111000001011_101_1_101110000010;
      patterns[28766] = 29'b0_111000001011_110_0_111000001011;
      patterns[28767] = 29'b0_111000001011_111_0_111000001011;
      patterns[28768] = 29'b0_111000001100_000_0_111000001100;
      patterns[28769] = 29'b0_111000001100_001_0_001100111000;
      patterns[28770] = 29'b0_111000001100_010_1_110000011000;
      patterns[28771] = 29'b0_111000001100_011_1_100000110001;
      patterns[28772] = 29'b0_111000001100_100_0_011100000110;
      patterns[28773] = 29'b0_111000001100_101_0_001110000011;
      patterns[28774] = 29'b0_111000001100_110_0_111000001100;
      patterns[28775] = 29'b0_111000001100_111_0_111000001100;
      patterns[28776] = 29'b0_111000001101_000_0_111000001101;
      patterns[28777] = 29'b0_111000001101_001_0_001101111000;
      patterns[28778] = 29'b0_111000001101_010_1_110000011010;
      patterns[28779] = 29'b0_111000001101_011_1_100000110101;
      patterns[28780] = 29'b0_111000001101_100_1_011100000110;
      patterns[28781] = 29'b0_111000001101_101_0_101110000011;
      patterns[28782] = 29'b0_111000001101_110_0_111000001101;
      patterns[28783] = 29'b0_111000001101_111_0_111000001101;
      patterns[28784] = 29'b0_111000001110_000_0_111000001110;
      patterns[28785] = 29'b0_111000001110_001_0_001110111000;
      patterns[28786] = 29'b0_111000001110_010_1_110000011100;
      patterns[28787] = 29'b0_111000001110_011_1_100000111001;
      patterns[28788] = 29'b0_111000001110_100_0_011100000111;
      patterns[28789] = 29'b0_111000001110_101_1_001110000011;
      patterns[28790] = 29'b0_111000001110_110_0_111000001110;
      patterns[28791] = 29'b0_111000001110_111_0_111000001110;
      patterns[28792] = 29'b0_111000001111_000_0_111000001111;
      patterns[28793] = 29'b0_111000001111_001_0_001111111000;
      patterns[28794] = 29'b0_111000001111_010_1_110000011110;
      patterns[28795] = 29'b0_111000001111_011_1_100000111101;
      patterns[28796] = 29'b0_111000001111_100_1_011100000111;
      patterns[28797] = 29'b0_111000001111_101_1_101110000011;
      patterns[28798] = 29'b0_111000001111_110_0_111000001111;
      patterns[28799] = 29'b0_111000001111_111_0_111000001111;
      patterns[28800] = 29'b0_111000010000_000_0_111000010000;
      patterns[28801] = 29'b0_111000010000_001_0_010000111000;
      patterns[28802] = 29'b0_111000010000_010_1_110000100000;
      patterns[28803] = 29'b0_111000010000_011_1_100001000001;
      patterns[28804] = 29'b0_111000010000_100_0_011100001000;
      patterns[28805] = 29'b0_111000010000_101_0_001110000100;
      patterns[28806] = 29'b0_111000010000_110_0_111000010000;
      patterns[28807] = 29'b0_111000010000_111_0_111000010000;
      patterns[28808] = 29'b0_111000010001_000_0_111000010001;
      patterns[28809] = 29'b0_111000010001_001_0_010001111000;
      patterns[28810] = 29'b0_111000010001_010_1_110000100010;
      patterns[28811] = 29'b0_111000010001_011_1_100001000101;
      patterns[28812] = 29'b0_111000010001_100_1_011100001000;
      patterns[28813] = 29'b0_111000010001_101_0_101110000100;
      patterns[28814] = 29'b0_111000010001_110_0_111000010001;
      patterns[28815] = 29'b0_111000010001_111_0_111000010001;
      patterns[28816] = 29'b0_111000010010_000_0_111000010010;
      patterns[28817] = 29'b0_111000010010_001_0_010010111000;
      patterns[28818] = 29'b0_111000010010_010_1_110000100100;
      patterns[28819] = 29'b0_111000010010_011_1_100001001001;
      patterns[28820] = 29'b0_111000010010_100_0_011100001001;
      patterns[28821] = 29'b0_111000010010_101_1_001110000100;
      patterns[28822] = 29'b0_111000010010_110_0_111000010010;
      patterns[28823] = 29'b0_111000010010_111_0_111000010010;
      patterns[28824] = 29'b0_111000010011_000_0_111000010011;
      patterns[28825] = 29'b0_111000010011_001_0_010011111000;
      patterns[28826] = 29'b0_111000010011_010_1_110000100110;
      patterns[28827] = 29'b0_111000010011_011_1_100001001101;
      patterns[28828] = 29'b0_111000010011_100_1_011100001001;
      patterns[28829] = 29'b0_111000010011_101_1_101110000100;
      patterns[28830] = 29'b0_111000010011_110_0_111000010011;
      patterns[28831] = 29'b0_111000010011_111_0_111000010011;
      patterns[28832] = 29'b0_111000010100_000_0_111000010100;
      patterns[28833] = 29'b0_111000010100_001_0_010100111000;
      patterns[28834] = 29'b0_111000010100_010_1_110000101000;
      patterns[28835] = 29'b0_111000010100_011_1_100001010001;
      patterns[28836] = 29'b0_111000010100_100_0_011100001010;
      patterns[28837] = 29'b0_111000010100_101_0_001110000101;
      patterns[28838] = 29'b0_111000010100_110_0_111000010100;
      patterns[28839] = 29'b0_111000010100_111_0_111000010100;
      patterns[28840] = 29'b0_111000010101_000_0_111000010101;
      patterns[28841] = 29'b0_111000010101_001_0_010101111000;
      patterns[28842] = 29'b0_111000010101_010_1_110000101010;
      patterns[28843] = 29'b0_111000010101_011_1_100001010101;
      patterns[28844] = 29'b0_111000010101_100_1_011100001010;
      patterns[28845] = 29'b0_111000010101_101_0_101110000101;
      patterns[28846] = 29'b0_111000010101_110_0_111000010101;
      patterns[28847] = 29'b0_111000010101_111_0_111000010101;
      patterns[28848] = 29'b0_111000010110_000_0_111000010110;
      patterns[28849] = 29'b0_111000010110_001_0_010110111000;
      patterns[28850] = 29'b0_111000010110_010_1_110000101100;
      patterns[28851] = 29'b0_111000010110_011_1_100001011001;
      patterns[28852] = 29'b0_111000010110_100_0_011100001011;
      patterns[28853] = 29'b0_111000010110_101_1_001110000101;
      patterns[28854] = 29'b0_111000010110_110_0_111000010110;
      patterns[28855] = 29'b0_111000010110_111_0_111000010110;
      patterns[28856] = 29'b0_111000010111_000_0_111000010111;
      patterns[28857] = 29'b0_111000010111_001_0_010111111000;
      patterns[28858] = 29'b0_111000010111_010_1_110000101110;
      patterns[28859] = 29'b0_111000010111_011_1_100001011101;
      patterns[28860] = 29'b0_111000010111_100_1_011100001011;
      patterns[28861] = 29'b0_111000010111_101_1_101110000101;
      patterns[28862] = 29'b0_111000010111_110_0_111000010111;
      patterns[28863] = 29'b0_111000010111_111_0_111000010111;
      patterns[28864] = 29'b0_111000011000_000_0_111000011000;
      patterns[28865] = 29'b0_111000011000_001_0_011000111000;
      patterns[28866] = 29'b0_111000011000_010_1_110000110000;
      patterns[28867] = 29'b0_111000011000_011_1_100001100001;
      patterns[28868] = 29'b0_111000011000_100_0_011100001100;
      patterns[28869] = 29'b0_111000011000_101_0_001110000110;
      patterns[28870] = 29'b0_111000011000_110_0_111000011000;
      patterns[28871] = 29'b0_111000011000_111_0_111000011000;
      patterns[28872] = 29'b0_111000011001_000_0_111000011001;
      patterns[28873] = 29'b0_111000011001_001_0_011001111000;
      patterns[28874] = 29'b0_111000011001_010_1_110000110010;
      patterns[28875] = 29'b0_111000011001_011_1_100001100101;
      patterns[28876] = 29'b0_111000011001_100_1_011100001100;
      patterns[28877] = 29'b0_111000011001_101_0_101110000110;
      patterns[28878] = 29'b0_111000011001_110_0_111000011001;
      patterns[28879] = 29'b0_111000011001_111_0_111000011001;
      patterns[28880] = 29'b0_111000011010_000_0_111000011010;
      patterns[28881] = 29'b0_111000011010_001_0_011010111000;
      patterns[28882] = 29'b0_111000011010_010_1_110000110100;
      patterns[28883] = 29'b0_111000011010_011_1_100001101001;
      patterns[28884] = 29'b0_111000011010_100_0_011100001101;
      patterns[28885] = 29'b0_111000011010_101_1_001110000110;
      patterns[28886] = 29'b0_111000011010_110_0_111000011010;
      patterns[28887] = 29'b0_111000011010_111_0_111000011010;
      patterns[28888] = 29'b0_111000011011_000_0_111000011011;
      patterns[28889] = 29'b0_111000011011_001_0_011011111000;
      patterns[28890] = 29'b0_111000011011_010_1_110000110110;
      patterns[28891] = 29'b0_111000011011_011_1_100001101101;
      patterns[28892] = 29'b0_111000011011_100_1_011100001101;
      patterns[28893] = 29'b0_111000011011_101_1_101110000110;
      patterns[28894] = 29'b0_111000011011_110_0_111000011011;
      patterns[28895] = 29'b0_111000011011_111_0_111000011011;
      patterns[28896] = 29'b0_111000011100_000_0_111000011100;
      patterns[28897] = 29'b0_111000011100_001_0_011100111000;
      patterns[28898] = 29'b0_111000011100_010_1_110000111000;
      patterns[28899] = 29'b0_111000011100_011_1_100001110001;
      patterns[28900] = 29'b0_111000011100_100_0_011100001110;
      patterns[28901] = 29'b0_111000011100_101_0_001110000111;
      patterns[28902] = 29'b0_111000011100_110_0_111000011100;
      patterns[28903] = 29'b0_111000011100_111_0_111000011100;
      patterns[28904] = 29'b0_111000011101_000_0_111000011101;
      patterns[28905] = 29'b0_111000011101_001_0_011101111000;
      patterns[28906] = 29'b0_111000011101_010_1_110000111010;
      patterns[28907] = 29'b0_111000011101_011_1_100001110101;
      patterns[28908] = 29'b0_111000011101_100_1_011100001110;
      patterns[28909] = 29'b0_111000011101_101_0_101110000111;
      patterns[28910] = 29'b0_111000011101_110_0_111000011101;
      patterns[28911] = 29'b0_111000011101_111_0_111000011101;
      patterns[28912] = 29'b0_111000011110_000_0_111000011110;
      patterns[28913] = 29'b0_111000011110_001_0_011110111000;
      patterns[28914] = 29'b0_111000011110_010_1_110000111100;
      patterns[28915] = 29'b0_111000011110_011_1_100001111001;
      patterns[28916] = 29'b0_111000011110_100_0_011100001111;
      patterns[28917] = 29'b0_111000011110_101_1_001110000111;
      patterns[28918] = 29'b0_111000011110_110_0_111000011110;
      patterns[28919] = 29'b0_111000011110_111_0_111000011110;
      patterns[28920] = 29'b0_111000011111_000_0_111000011111;
      patterns[28921] = 29'b0_111000011111_001_0_011111111000;
      patterns[28922] = 29'b0_111000011111_010_1_110000111110;
      patterns[28923] = 29'b0_111000011111_011_1_100001111101;
      patterns[28924] = 29'b0_111000011111_100_1_011100001111;
      patterns[28925] = 29'b0_111000011111_101_1_101110000111;
      patterns[28926] = 29'b0_111000011111_110_0_111000011111;
      patterns[28927] = 29'b0_111000011111_111_0_111000011111;
      patterns[28928] = 29'b0_111000100000_000_0_111000100000;
      patterns[28929] = 29'b0_111000100000_001_0_100000111000;
      patterns[28930] = 29'b0_111000100000_010_1_110001000000;
      patterns[28931] = 29'b0_111000100000_011_1_100010000001;
      patterns[28932] = 29'b0_111000100000_100_0_011100010000;
      patterns[28933] = 29'b0_111000100000_101_0_001110001000;
      patterns[28934] = 29'b0_111000100000_110_0_111000100000;
      patterns[28935] = 29'b0_111000100000_111_0_111000100000;
      patterns[28936] = 29'b0_111000100001_000_0_111000100001;
      patterns[28937] = 29'b0_111000100001_001_0_100001111000;
      patterns[28938] = 29'b0_111000100001_010_1_110001000010;
      patterns[28939] = 29'b0_111000100001_011_1_100010000101;
      patterns[28940] = 29'b0_111000100001_100_1_011100010000;
      patterns[28941] = 29'b0_111000100001_101_0_101110001000;
      patterns[28942] = 29'b0_111000100001_110_0_111000100001;
      patterns[28943] = 29'b0_111000100001_111_0_111000100001;
      patterns[28944] = 29'b0_111000100010_000_0_111000100010;
      patterns[28945] = 29'b0_111000100010_001_0_100010111000;
      patterns[28946] = 29'b0_111000100010_010_1_110001000100;
      patterns[28947] = 29'b0_111000100010_011_1_100010001001;
      patterns[28948] = 29'b0_111000100010_100_0_011100010001;
      patterns[28949] = 29'b0_111000100010_101_1_001110001000;
      patterns[28950] = 29'b0_111000100010_110_0_111000100010;
      patterns[28951] = 29'b0_111000100010_111_0_111000100010;
      patterns[28952] = 29'b0_111000100011_000_0_111000100011;
      patterns[28953] = 29'b0_111000100011_001_0_100011111000;
      patterns[28954] = 29'b0_111000100011_010_1_110001000110;
      patterns[28955] = 29'b0_111000100011_011_1_100010001101;
      patterns[28956] = 29'b0_111000100011_100_1_011100010001;
      patterns[28957] = 29'b0_111000100011_101_1_101110001000;
      patterns[28958] = 29'b0_111000100011_110_0_111000100011;
      patterns[28959] = 29'b0_111000100011_111_0_111000100011;
      patterns[28960] = 29'b0_111000100100_000_0_111000100100;
      patterns[28961] = 29'b0_111000100100_001_0_100100111000;
      patterns[28962] = 29'b0_111000100100_010_1_110001001000;
      patterns[28963] = 29'b0_111000100100_011_1_100010010001;
      patterns[28964] = 29'b0_111000100100_100_0_011100010010;
      patterns[28965] = 29'b0_111000100100_101_0_001110001001;
      patterns[28966] = 29'b0_111000100100_110_0_111000100100;
      patterns[28967] = 29'b0_111000100100_111_0_111000100100;
      patterns[28968] = 29'b0_111000100101_000_0_111000100101;
      patterns[28969] = 29'b0_111000100101_001_0_100101111000;
      patterns[28970] = 29'b0_111000100101_010_1_110001001010;
      patterns[28971] = 29'b0_111000100101_011_1_100010010101;
      patterns[28972] = 29'b0_111000100101_100_1_011100010010;
      patterns[28973] = 29'b0_111000100101_101_0_101110001001;
      patterns[28974] = 29'b0_111000100101_110_0_111000100101;
      patterns[28975] = 29'b0_111000100101_111_0_111000100101;
      patterns[28976] = 29'b0_111000100110_000_0_111000100110;
      patterns[28977] = 29'b0_111000100110_001_0_100110111000;
      patterns[28978] = 29'b0_111000100110_010_1_110001001100;
      patterns[28979] = 29'b0_111000100110_011_1_100010011001;
      patterns[28980] = 29'b0_111000100110_100_0_011100010011;
      patterns[28981] = 29'b0_111000100110_101_1_001110001001;
      patterns[28982] = 29'b0_111000100110_110_0_111000100110;
      patterns[28983] = 29'b0_111000100110_111_0_111000100110;
      patterns[28984] = 29'b0_111000100111_000_0_111000100111;
      patterns[28985] = 29'b0_111000100111_001_0_100111111000;
      patterns[28986] = 29'b0_111000100111_010_1_110001001110;
      patterns[28987] = 29'b0_111000100111_011_1_100010011101;
      patterns[28988] = 29'b0_111000100111_100_1_011100010011;
      patterns[28989] = 29'b0_111000100111_101_1_101110001001;
      patterns[28990] = 29'b0_111000100111_110_0_111000100111;
      patterns[28991] = 29'b0_111000100111_111_0_111000100111;
      patterns[28992] = 29'b0_111000101000_000_0_111000101000;
      patterns[28993] = 29'b0_111000101000_001_0_101000111000;
      patterns[28994] = 29'b0_111000101000_010_1_110001010000;
      patterns[28995] = 29'b0_111000101000_011_1_100010100001;
      patterns[28996] = 29'b0_111000101000_100_0_011100010100;
      patterns[28997] = 29'b0_111000101000_101_0_001110001010;
      patterns[28998] = 29'b0_111000101000_110_0_111000101000;
      patterns[28999] = 29'b0_111000101000_111_0_111000101000;
      patterns[29000] = 29'b0_111000101001_000_0_111000101001;
      patterns[29001] = 29'b0_111000101001_001_0_101001111000;
      patterns[29002] = 29'b0_111000101001_010_1_110001010010;
      patterns[29003] = 29'b0_111000101001_011_1_100010100101;
      patterns[29004] = 29'b0_111000101001_100_1_011100010100;
      patterns[29005] = 29'b0_111000101001_101_0_101110001010;
      patterns[29006] = 29'b0_111000101001_110_0_111000101001;
      patterns[29007] = 29'b0_111000101001_111_0_111000101001;
      patterns[29008] = 29'b0_111000101010_000_0_111000101010;
      patterns[29009] = 29'b0_111000101010_001_0_101010111000;
      patterns[29010] = 29'b0_111000101010_010_1_110001010100;
      patterns[29011] = 29'b0_111000101010_011_1_100010101001;
      patterns[29012] = 29'b0_111000101010_100_0_011100010101;
      patterns[29013] = 29'b0_111000101010_101_1_001110001010;
      patterns[29014] = 29'b0_111000101010_110_0_111000101010;
      patterns[29015] = 29'b0_111000101010_111_0_111000101010;
      patterns[29016] = 29'b0_111000101011_000_0_111000101011;
      patterns[29017] = 29'b0_111000101011_001_0_101011111000;
      patterns[29018] = 29'b0_111000101011_010_1_110001010110;
      patterns[29019] = 29'b0_111000101011_011_1_100010101101;
      patterns[29020] = 29'b0_111000101011_100_1_011100010101;
      patterns[29021] = 29'b0_111000101011_101_1_101110001010;
      patterns[29022] = 29'b0_111000101011_110_0_111000101011;
      patterns[29023] = 29'b0_111000101011_111_0_111000101011;
      patterns[29024] = 29'b0_111000101100_000_0_111000101100;
      patterns[29025] = 29'b0_111000101100_001_0_101100111000;
      patterns[29026] = 29'b0_111000101100_010_1_110001011000;
      patterns[29027] = 29'b0_111000101100_011_1_100010110001;
      patterns[29028] = 29'b0_111000101100_100_0_011100010110;
      patterns[29029] = 29'b0_111000101100_101_0_001110001011;
      patterns[29030] = 29'b0_111000101100_110_0_111000101100;
      patterns[29031] = 29'b0_111000101100_111_0_111000101100;
      patterns[29032] = 29'b0_111000101101_000_0_111000101101;
      patterns[29033] = 29'b0_111000101101_001_0_101101111000;
      patterns[29034] = 29'b0_111000101101_010_1_110001011010;
      patterns[29035] = 29'b0_111000101101_011_1_100010110101;
      patterns[29036] = 29'b0_111000101101_100_1_011100010110;
      patterns[29037] = 29'b0_111000101101_101_0_101110001011;
      patterns[29038] = 29'b0_111000101101_110_0_111000101101;
      patterns[29039] = 29'b0_111000101101_111_0_111000101101;
      patterns[29040] = 29'b0_111000101110_000_0_111000101110;
      patterns[29041] = 29'b0_111000101110_001_0_101110111000;
      patterns[29042] = 29'b0_111000101110_010_1_110001011100;
      patterns[29043] = 29'b0_111000101110_011_1_100010111001;
      patterns[29044] = 29'b0_111000101110_100_0_011100010111;
      patterns[29045] = 29'b0_111000101110_101_1_001110001011;
      patterns[29046] = 29'b0_111000101110_110_0_111000101110;
      patterns[29047] = 29'b0_111000101110_111_0_111000101110;
      patterns[29048] = 29'b0_111000101111_000_0_111000101111;
      patterns[29049] = 29'b0_111000101111_001_0_101111111000;
      patterns[29050] = 29'b0_111000101111_010_1_110001011110;
      patterns[29051] = 29'b0_111000101111_011_1_100010111101;
      patterns[29052] = 29'b0_111000101111_100_1_011100010111;
      patterns[29053] = 29'b0_111000101111_101_1_101110001011;
      patterns[29054] = 29'b0_111000101111_110_0_111000101111;
      patterns[29055] = 29'b0_111000101111_111_0_111000101111;
      patterns[29056] = 29'b0_111000110000_000_0_111000110000;
      patterns[29057] = 29'b0_111000110000_001_0_110000111000;
      patterns[29058] = 29'b0_111000110000_010_1_110001100000;
      patterns[29059] = 29'b0_111000110000_011_1_100011000001;
      patterns[29060] = 29'b0_111000110000_100_0_011100011000;
      patterns[29061] = 29'b0_111000110000_101_0_001110001100;
      patterns[29062] = 29'b0_111000110000_110_0_111000110000;
      patterns[29063] = 29'b0_111000110000_111_0_111000110000;
      patterns[29064] = 29'b0_111000110001_000_0_111000110001;
      patterns[29065] = 29'b0_111000110001_001_0_110001111000;
      patterns[29066] = 29'b0_111000110001_010_1_110001100010;
      patterns[29067] = 29'b0_111000110001_011_1_100011000101;
      patterns[29068] = 29'b0_111000110001_100_1_011100011000;
      patterns[29069] = 29'b0_111000110001_101_0_101110001100;
      patterns[29070] = 29'b0_111000110001_110_0_111000110001;
      patterns[29071] = 29'b0_111000110001_111_0_111000110001;
      patterns[29072] = 29'b0_111000110010_000_0_111000110010;
      patterns[29073] = 29'b0_111000110010_001_0_110010111000;
      patterns[29074] = 29'b0_111000110010_010_1_110001100100;
      patterns[29075] = 29'b0_111000110010_011_1_100011001001;
      patterns[29076] = 29'b0_111000110010_100_0_011100011001;
      patterns[29077] = 29'b0_111000110010_101_1_001110001100;
      patterns[29078] = 29'b0_111000110010_110_0_111000110010;
      patterns[29079] = 29'b0_111000110010_111_0_111000110010;
      patterns[29080] = 29'b0_111000110011_000_0_111000110011;
      patterns[29081] = 29'b0_111000110011_001_0_110011111000;
      patterns[29082] = 29'b0_111000110011_010_1_110001100110;
      patterns[29083] = 29'b0_111000110011_011_1_100011001101;
      patterns[29084] = 29'b0_111000110011_100_1_011100011001;
      patterns[29085] = 29'b0_111000110011_101_1_101110001100;
      patterns[29086] = 29'b0_111000110011_110_0_111000110011;
      patterns[29087] = 29'b0_111000110011_111_0_111000110011;
      patterns[29088] = 29'b0_111000110100_000_0_111000110100;
      patterns[29089] = 29'b0_111000110100_001_0_110100111000;
      patterns[29090] = 29'b0_111000110100_010_1_110001101000;
      patterns[29091] = 29'b0_111000110100_011_1_100011010001;
      patterns[29092] = 29'b0_111000110100_100_0_011100011010;
      patterns[29093] = 29'b0_111000110100_101_0_001110001101;
      patterns[29094] = 29'b0_111000110100_110_0_111000110100;
      patterns[29095] = 29'b0_111000110100_111_0_111000110100;
      patterns[29096] = 29'b0_111000110101_000_0_111000110101;
      patterns[29097] = 29'b0_111000110101_001_0_110101111000;
      patterns[29098] = 29'b0_111000110101_010_1_110001101010;
      patterns[29099] = 29'b0_111000110101_011_1_100011010101;
      patterns[29100] = 29'b0_111000110101_100_1_011100011010;
      patterns[29101] = 29'b0_111000110101_101_0_101110001101;
      patterns[29102] = 29'b0_111000110101_110_0_111000110101;
      patterns[29103] = 29'b0_111000110101_111_0_111000110101;
      patterns[29104] = 29'b0_111000110110_000_0_111000110110;
      patterns[29105] = 29'b0_111000110110_001_0_110110111000;
      patterns[29106] = 29'b0_111000110110_010_1_110001101100;
      patterns[29107] = 29'b0_111000110110_011_1_100011011001;
      patterns[29108] = 29'b0_111000110110_100_0_011100011011;
      patterns[29109] = 29'b0_111000110110_101_1_001110001101;
      patterns[29110] = 29'b0_111000110110_110_0_111000110110;
      patterns[29111] = 29'b0_111000110110_111_0_111000110110;
      patterns[29112] = 29'b0_111000110111_000_0_111000110111;
      patterns[29113] = 29'b0_111000110111_001_0_110111111000;
      patterns[29114] = 29'b0_111000110111_010_1_110001101110;
      patterns[29115] = 29'b0_111000110111_011_1_100011011101;
      patterns[29116] = 29'b0_111000110111_100_1_011100011011;
      patterns[29117] = 29'b0_111000110111_101_1_101110001101;
      patterns[29118] = 29'b0_111000110111_110_0_111000110111;
      patterns[29119] = 29'b0_111000110111_111_0_111000110111;
      patterns[29120] = 29'b0_111000111000_000_0_111000111000;
      patterns[29121] = 29'b0_111000111000_001_0_111000111000;
      patterns[29122] = 29'b0_111000111000_010_1_110001110000;
      patterns[29123] = 29'b0_111000111000_011_1_100011100001;
      patterns[29124] = 29'b0_111000111000_100_0_011100011100;
      patterns[29125] = 29'b0_111000111000_101_0_001110001110;
      patterns[29126] = 29'b0_111000111000_110_0_111000111000;
      patterns[29127] = 29'b0_111000111000_111_0_111000111000;
      patterns[29128] = 29'b0_111000111001_000_0_111000111001;
      patterns[29129] = 29'b0_111000111001_001_0_111001111000;
      patterns[29130] = 29'b0_111000111001_010_1_110001110010;
      patterns[29131] = 29'b0_111000111001_011_1_100011100101;
      patterns[29132] = 29'b0_111000111001_100_1_011100011100;
      patterns[29133] = 29'b0_111000111001_101_0_101110001110;
      patterns[29134] = 29'b0_111000111001_110_0_111000111001;
      patterns[29135] = 29'b0_111000111001_111_0_111000111001;
      patterns[29136] = 29'b0_111000111010_000_0_111000111010;
      patterns[29137] = 29'b0_111000111010_001_0_111010111000;
      patterns[29138] = 29'b0_111000111010_010_1_110001110100;
      patterns[29139] = 29'b0_111000111010_011_1_100011101001;
      patterns[29140] = 29'b0_111000111010_100_0_011100011101;
      patterns[29141] = 29'b0_111000111010_101_1_001110001110;
      patterns[29142] = 29'b0_111000111010_110_0_111000111010;
      patterns[29143] = 29'b0_111000111010_111_0_111000111010;
      patterns[29144] = 29'b0_111000111011_000_0_111000111011;
      patterns[29145] = 29'b0_111000111011_001_0_111011111000;
      patterns[29146] = 29'b0_111000111011_010_1_110001110110;
      patterns[29147] = 29'b0_111000111011_011_1_100011101101;
      patterns[29148] = 29'b0_111000111011_100_1_011100011101;
      patterns[29149] = 29'b0_111000111011_101_1_101110001110;
      patterns[29150] = 29'b0_111000111011_110_0_111000111011;
      patterns[29151] = 29'b0_111000111011_111_0_111000111011;
      patterns[29152] = 29'b0_111000111100_000_0_111000111100;
      patterns[29153] = 29'b0_111000111100_001_0_111100111000;
      patterns[29154] = 29'b0_111000111100_010_1_110001111000;
      patterns[29155] = 29'b0_111000111100_011_1_100011110001;
      patterns[29156] = 29'b0_111000111100_100_0_011100011110;
      patterns[29157] = 29'b0_111000111100_101_0_001110001111;
      patterns[29158] = 29'b0_111000111100_110_0_111000111100;
      patterns[29159] = 29'b0_111000111100_111_0_111000111100;
      patterns[29160] = 29'b0_111000111101_000_0_111000111101;
      patterns[29161] = 29'b0_111000111101_001_0_111101111000;
      patterns[29162] = 29'b0_111000111101_010_1_110001111010;
      patterns[29163] = 29'b0_111000111101_011_1_100011110101;
      patterns[29164] = 29'b0_111000111101_100_1_011100011110;
      patterns[29165] = 29'b0_111000111101_101_0_101110001111;
      patterns[29166] = 29'b0_111000111101_110_0_111000111101;
      patterns[29167] = 29'b0_111000111101_111_0_111000111101;
      patterns[29168] = 29'b0_111000111110_000_0_111000111110;
      patterns[29169] = 29'b0_111000111110_001_0_111110111000;
      patterns[29170] = 29'b0_111000111110_010_1_110001111100;
      patterns[29171] = 29'b0_111000111110_011_1_100011111001;
      patterns[29172] = 29'b0_111000111110_100_0_011100011111;
      patterns[29173] = 29'b0_111000111110_101_1_001110001111;
      patterns[29174] = 29'b0_111000111110_110_0_111000111110;
      patterns[29175] = 29'b0_111000111110_111_0_111000111110;
      patterns[29176] = 29'b0_111000111111_000_0_111000111111;
      patterns[29177] = 29'b0_111000111111_001_0_111111111000;
      patterns[29178] = 29'b0_111000111111_010_1_110001111110;
      patterns[29179] = 29'b0_111000111111_011_1_100011111101;
      patterns[29180] = 29'b0_111000111111_100_1_011100011111;
      patterns[29181] = 29'b0_111000111111_101_1_101110001111;
      patterns[29182] = 29'b0_111000111111_110_0_111000111111;
      patterns[29183] = 29'b0_111000111111_111_0_111000111111;
      patterns[29184] = 29'b0_111001000000_000_0_111001000000;
      patterns[29185] = 29'b0_111001000000_001_0_000000111001;
      patterns[29186] = 29'b0_111001000000_010_1_110010000000;
      patterns[29187] = 29'b0_111001000000_011_1_100100000001;
      patterns[29188] = 29'b0_111001000000_100_0_011100100000;
      patterns[29189] = 29'b0_111001000000_101_0_001110010000;
      patterns[29190] = 29'b0_111001000000_110_0_111001000000;
      patterns[29191] = 29'b0_111001000000_111_0_111001000000;
      patterns[29192] = 29'b0_111001000001_000_0_111001000001;
      patterns[29193] = 29'b0_111001000001_001_0_000001111001;
      patterns[29194] = 29'b0_111001000001_010_1_110010000010;
      patterns[29195] = 29'b0_111001000001_011_1_100100000101;
      patterns[29196] = 29'b0_111001000001_100_1_011100100000;
      patterns[29197] = 29'b0_111001000001_101_0_101110010000;
      patterns[29198] = 29'b0_111001000001_110_0_111001000001;
      patterns[29199] = 29'b0_111001000001_111_0_111001000001;
      patterns[29200] = 29'b0_111001000010_000_0_111001000010;
      patterns[29201] = 29'b0_111001000010_001_0_000010111001;
      patterns[29202] = 29'b0_111001000010_010_1_110010000100;
      patterns[29203] = 29'b0_111001000010_011_1_100100001001;
      patterns[29204] = 29'b0_111001000010_100_0_011100100001;
      patterns[29205] = 29'b0_111001000010_101_1_001110010000;
      patterns[29206] = 29'b0_111001000010_110_0_111001000010;
      patterns[29207] = 29'b0_111001000010_111_0_111001000010;
      patterns[29208] = 29'b0_111001000011_000_0_111001000011;
      patterns[29209] = 29'b0_111001000011_001_0_000011111001;
      patterns[29210] = 29'b0_111001000011_010_1_110010000110;
      patterns[29211] = 29'b0_111001000011_011_1_100100001101;
      patterns[29212] = 29'b0_111001000011_100_1_011100100001;
      patterns[29213] = 29'b0_111001000011_101_1_101110010000;
      patterns[29214] = 29'b0_111001000011_110_0_111001000011;
      patterns[29215] = 29'b0_111001000011_111_0_111001000011;
      patterns[29216] = 29'b0_111001000100_000_0_111001000100;
      patterns[29217] = 29'b0_111001000100_001_0_000100111001;
      patterns[29218] = 29'b0_111001000100_010_1_110010001000;
      patterns[29219] = 29'b0_111001000100_011_1_100100010001;
      patterns[29220] = 29'b0_111001000100_100_0_011100100010;
      patterns[29221] = 29'b0_111001000100_101_0_001110010001;
      patterns[29222] = 29'b0_111001000100_110_0_111001000100;
      patterns[29223] = 29'b0_111001000100_111_0_111001000100;
      patterns[29224] = 29'b0_111001000101_000_0_111001000101;
      patterns[29225] = 29'b0_111001000101_001_0_000101111001;
      patterns[29226] = 29'b0_111001000101_010_1_110010001010;
      patterns[29227] = 29'b0_111001000101_011_1_100100010101;
      patterns[29228] = 29'b0_111001000101_100_1_011100100010;
      patterns[29229] = 29'b0_111001000101_101_0_101110010001;
      patterns[29230] = 29'b0_111001000101_110_0_111001000101;
      patterns[29231] = 29'b0_111001000101_111_0_111001000101;
      patterns[29232] = 29'b0_111001000110_000_0_111001000110;
      patterns[29233] = 29'b0_111001000110_001_0_000110111001;
      patterns[29234] = 29'b0_111001000110_010_1_110010001100;
      patterns[29235] = 29'b0_111001000110_011_1_100100011001;
      patterns[29236] = 29'b0_111001000110_100_0_011100100011;
      patterns[29237] = 29'b0_111001000110_101_1_001110010001;
      patterns[29238] = 29'b0_111001000110_110_0_111001000110;
      patterns[29239] = 29'b0_111001000110_111_0_111001000110;
      patterns[29240] = 29'b0_111001000111_000_0_111001000111;
      patterns[29241] = 29'b0_111001000111_001_0_000111111001;
      patterns[29242] = 29'b0_111001000111_010_1_110010001110;
      patterns[29243] = 29'b0_111001000111_011_1_100100011101;
      patterns[29244] = 29'b0_111001000111_100_1_011100100011;
      patterns[29245] = 29'b0_111001000111_101_1_101110010001;
      patterns[29246] = 29'b0_111001000111_110_0_111001000111;
      patterns[29247] = 29'b0_111001000111_111_0_111001000111;
      patterns[29248] = 29'b0_111001001000_000_0_111001001000;
      patterns[29249] = 29'b0_111001001000_001_0_001000111001;
      patterns[29250] = 29'b0_111001001000_010_1_110010010000;
      patterns[29251] = 29'b0_111001001000_011_1_100100100001;
      patterns[29252] = 29'b0_111001001000_100_0_011100100100;
      patterns[29253] = 29'b0_111001001000_101_0_001110010010;
      patterns[29254] = 29'b0_111001001000_110_0_111001001000;
      patterns[29255] = 29'b0_111001001000_111_0_111001001000;
      patterns[29256] = 29'b0_111001001001_000_0_111001001001;
      patterns[29257] = 29'b0_111001001001_001_0_001001111001;
      patterns[29258] = 29'b0_111001001001_010_1_110010010010;
      patterns[29259] = 29'b0_111001001001_011_1_100100100101;
      patterns[29260] = 29'b0_111001001001_100_1_011100100100;
      patterns[29261] = 29'b0_111001001001_101_0_101110010010;
      patterns[29262] = 29'b0_111001001001_110_0_111001001001;
      patterns[29263] = 29'b0_111001001001_111_0_111001001001;
      patterns[29264] = 29'b0_111001001010_000_0_111001001010;
      patterns[29265] = 29'b0_111001001010_001_0_001010111001;
      patterns[29266] = 29'b0_111001001010_010_1_110010010100;
      patterns[29267] = 29'b0_111001001010_011_1_100100101001;
      patterns[29268] = 29'b0_111001001010_100_0_011100100101;
      patterns[29269] = 29'b0_111001001010_101_1_001110010010;
      patterns[29270] = 29'b0_111001001010_110_0_111001001010;
      patterns[29271] = 29'b0_111001001010_111_0_111001001010;
      patterns[29272] = 29'b0_111001001011_000_0_111001001011;
      patterns[29273] = 29'b0_111001001011_001_0_001011111001;
      patterns[29274] = 29'b0_111001001011_010_1_110010010110;
      patterns[29275] = 29'b0_111001001011_011_1_100100101101;
      patterns[29276] = 29'b0_111001001011_100_1_011100100101;
      patterns[29277] = 29'b0_111001001011_101_1_101110010010;
      patterns[29278] = 29'b0_111001001011_110_0_111001001011;
      patterns[29279] = 29'b0_111001001011_111_0_111001001011;
      patterns[29280] = 29'b0_111001001100_000_0_111001001100;
      patterns[29281] = 29'b0_111001001100_001_0_001100111001;
      patterns[29282] = 29'b0_111001001100_010_1_110010011000;
      patterns[29283] = 29'b0_111001001100_011_1_100100110001;
      patterns[29284] = 29'b0_111001001100_100_0_011100100110;
      patterns[29285] = 29'b0_111001001100_101_0_001110010011;
      patterns[29286] = 29'b0_111001001100_110_0_111001001100;
      patterns[29287] = 29'b0_111001001100_111_0_111001001100;
      patterns[29288] = 29'b0_111001001101_000_0_111001001101;
      patterns[29289] = 29'b0_111001001101_001_0_001101111001;
      patterns[29290] = 29'b0_111001001101_010_1_110010011010;
      patterns[29291] = 29'b0_111001001101_011_1_100100110101;
      patterns[29292] = 29'b0_111001001101_100_1_011100100110;
      patterns[29293] = 29'b0_111001001101_101_0_101110010011;
      patterns[29294] = 29'b0_111001001101_110_0_111001001101;
      patterns[29295] = 29'b0_111001001101_111_0_111001001101;
      patterns[29296] = 29'b0_111001001110_000_0_111001001110;
      patterns[29297] = 29'b0_111001001110_001_0_001110111001;
      patterns[29298] = 29'b0_111001001110_010_1_110010011100;
      patterns[29299] = 29'b0_111001001110_011_1_100100111001;
      patterns[29300] = 29'b0_111001001110_100_0_011100100111;
      patterns[29301] = 29'b0_111001001110_101_1_001110010011;
      patterns[29302] = 29'b0_111001001110_110_0_111001001110;
      patterns[29303] = 29'b0_111001001110_111_0_111001001110;
      patterns[29304] = 29'b0_111001001111_000_0_111001001111;
      patterns[29305] = 29'b0_111001001111_001_0_001111111001;
      patterns[29306] = 29'b0_111001001111_010_1_110010011110;
      patterns[29307] = 29'b0_111001001111_011_1_100100111101;
      patterns[29308] = 29'b0_111001001111_100_1_011100100111;
      patterns[29309] = 29'b0_111001001111_101_1_101110010011;
      patterns[29310] = 29'b0_111001001111_110_0_111001001111;
      patterns[29311] = 29'b0_111001001111_111_0_111001001111;
      patterns[29312] = 29'b0_111001010000_000_0_111001010000;
      patterns[29313] = 29'b0_111001010000_001_0_010000111001;
      patterns[29314] = 29'b0_111001010000_010_1_110010100000;
      patterns[29315] = 29'b0_111001010000_011_1_100101000001;
      patterns[29316] = 29'b0_111001010000_100_0_011100101000;
      patterns[29317] = 29'b0_111001010000_101_0_001110010100;
      patterns[29318] = 29'b0_111001010000_110_0_111001010000;
      patterns[29319] = 29'b0_111001010000_111_0_111001010000;
      patterns[29320] = 29'b0_111001010001_000_0_111001010001;
      patterns[29321] = 29'b0_111001010001_001_0_010001111001;
      patterns[29322] = 29'b0_111001010001_010_1_110010100010;
      patterns[29323] = 29'b0_111001010001_011_1_100101000101;
      patterns[29324] = 29'b0_111001010001_100_1_011100101000;
      patterns[29325] = 29'b0_111001010001_101_0_101110010100;
      patterns[29326] = 29'b0_111001010001_110_0_111001010001;
      patterns[29327] = 29'b0_111001010001_111_0_111001010001;
      patterns[29328] = 29'b0_111001010010_000_0_111001010010;
      patterns[29329] = 29'b0_111001010010_001_0_010010111001;
      patterns[29330] = 29'b0_111001010010_010_1_110010100100;
      patterns[29331] = 29'b0_111001010010_011_1_100101001001;
      patterns[29332] = 29'b0_111001010010_100_0_011100101001;
      patterns[29333] = 29'b0_111001010010_101_1_001110010100;
      patterns[29334] = 29'b0_111001010010_110_0_111001010010;
      patterns[29335] = 29'b0_111001010010_111_0_111001010010;
      patterns[29336] = 29'b0_111001010011_000_0_111001010011;
      patterns[29337] = 29'b0_111001010011_001_0_010011111001;
      patterns[29338] = 29'b0_111001010011_010_1_110010100110;
      patterns[29339] = 29'b0_111001010011_011_1_100101001101;
      patterns[29340] = 29'b0_111001010011_100_1_011100101001;
      patterns[29341] = 29'b0_111001010011_101_1_101110010100;
      patterns[29342] = 29'b0_111001010011_110_0_111001010011;
      patterns[29343] = 29'b0_111001010011_111_0_111001010011;
      patterns[29344] = 29'b0_111001010100_000_0_111001010100;
      patterns[29345] = 29'b0_111001010100_001_0_010100111001;
      patterns[29346] = 29'b0_111001010100_010_1_110010101000;
      patterns[29347] = 29'b0_111001010100_011_1_100101010001;
      patterns[29348] = 29'b0_111001010100_100_0_011100101010;
      patterns[29349] = 29'b0_111001010100_101_0_001110010101;
      patterns[29350] = 29'b0_111001010100_110_0_111001010100;
      patterns[29351] = 29'b0_111001010100_111_0_111001010100;
      patterns[29352] = 29'b0_111001010101_000_0_111001010101;
      patterns[29353] = 29'b0_111001010101_001_0_010101111001;
      patterns[29354] = 29'b0_111001010101_010_1_110010101010;
      patterns[29355] = 29'b0_111001010101_011_1_100101010101;
      patterns[29356] = 29'b0_111001010101_100_1_011100101010;
      patterns[29357] = 29'b0_111001010101_101_0_101110010101;
      patterns[29358] = 29'b0_111001010101_110_0_111001010101;
      patterns[29359] = 29'b0_111001010101_111_0_111001010101;
      patterns[29360] = 29'b0_111001010110_000_0_111001010110;
      patterns[29361] = 29'b0_111001010110_001_0_010110111001;
      patterns[29362] = 29'b0_111001010110_010_1_110010101100;
      patterns[29363] = 29'b0_111001010110_011_1_100101011001;
      patterns[29364] = 29'b0_111001010110_100_0_011100101011;
      patterns[29365] = 29'b0_111001010110_101_1_001110010101;
      patterns[29366] = 29'b0_111001010110_110_0_111001010110;
      patterns[29367] = 29'b0_111001010110_111_0_111001010110;
      patterns[29368] = 29'b0_111001010111_000_0_111001010111;
      patterns[29369] = 29'b0_111001010111_001_0_010111111001;
      patterns[29370] = 29'b0_111001010111_010_1_110010101110;
      patterns[29371] = 29'b0_111001010111_011_1_100101011101;
      patterns[29372] = 29'b0_111001010111_100_1_011100101011;
      patterns[29373] = 29'b0_111001010111_101_1_101110010101;
      patterns[29374] = 29'b0_111001010111_110_0_111001010111;
      patterns[29375] = 29'b0_111001010111_111_0_111001010111;
      patterns[29376] = 29'b0_111001011000_000_0_111001011000;
      patterns[29377] = 29'b0_111001011000_001_0_011000111001;
      patterns[29378] = 29'b0_111001011000_010_1_110010110000;
      patterns[29379] = 29'b0_111001011000_011_1_100101100001;
      patterns[29380] = 29'b0_111001011000_100_0_011100101100;
      patterns[29381] = 29'b0_111001011000_101_0_001110010110;
      patterns[29382] = 29'b0_111001011000_110_0_111001011000;
      patterns[29383] = 29'b0_111001011000_111_0_111001011000;
      patterns[29384] = 29'b0_111001011001_000_0_111001011001;
      patterns[29385] = 29'b0_111001011001_001_0_011001111001;
      patterns[29386] = 29'b0_111001011001_010_1_110010110010;
      patterns[29387] = 29'b0_111001011001_011_1_100101100101;
      patterns[29388] = 29'b0_111001011001_100_1_011100101100;
      patterns[29389] = 29'b0_111001011001_101_0_101110010110;
      patterns[29390] = 29'b0_111001011001_110_0_111001011001;
      patterns[29391] = 29'b0_111001011001_111_0_111001011001;
      patterns[29392] = 29'b0_111001011010_000_0_111001011010;
      patterns[29393] = 29'b0_111001011010_001_0_011010111001;
      patterns[29394] = 29'b0_111001011010_010_1_110010110100;
      patterns[29395] = 29'b0_111001011010_011_1_100101101001;
      patterns[29396] = 29'b0_111001011010_100_0_011100101101;
      patterns[29397] = 29'b0_111001011010_101_1_001110010110;
      patterns[29398] = 29'b0_111001011010_110_0_111001011010;
      patterns[29399] = 29'b0_111001011010_111_0_111001011010;
      patterns[29400] = 29'b0_111001011011_000_0_111001011011;
      patterns[29401] = 29'b0_111001011011_001_0_011011111001;
      patterns[29402] = 29'b0_111001011011_010_1_110010110110;
      patterns[29403] = 29'b0_111001011011_011_1_100101101101;
      patterns[29404] = 29'b0_111001011011_100_1_011100101101;
      patterns[29405] = 29'b0_111001011011_101_1_101110010110;
      patterns[29406] = 29'b0_111001011011_110_0_111001011011;
      patterns[29407] = 29'b0_111001011011_111_0_111001011011;
      patterns[29408] = 29'b0_111001011100_000_0_111001011100;
      patterns[29409] = 29'b0_111001011100_001_0_011100111001;
      patterns[29410] = 29'b0_111001011100_010_1_110010111000;
      patterns[29411] = 29'b0_111001011100_011_1_100101110001;
      patterns[29412] = 29'b0_111001011100_100_0_011100101110;
      patterns[29413] = 29'b0_111001011100_101_0_001110010111;
      patterns[29414] = 29'b0_111001011100_110_0_111001011100;
      patterns[29415] = 29'b0_111001011100_111_0_111001011100;
      patterns[29416] = 29'b0_111001011101_000_0_111001011101;
      patterns[29417] = 29'b0_111001011101_001_0_011101111001;
      patterns[29418] = 29'b0_111001011101_010_1_110010111010;
      patterns[29419] = 29'b0_111001011101_011_1_100101110101;
      patterns[29420] = 29'b0_111001011101_100_1_011100101110;
      patterns[29421] = 29'b0_111001011101_101_0_101110010111;
      patterns[29422] = 29'b0_111001011101_110_0_111001011101;
      patterns[29423] = 29'b0_111001011101_111_0_111001011101;
      patterns[29424] = 29'b0_111001011110_000_0_111001011110;
      patterns[29425] = 29'b0_111001011110_001_0_011110111001;
      patterns[29426] = 29'b0_111001011110_010_1_110010111100;
      patterns[29427] = 29'b0_111001011110_011_1_100101111001;
      patterns[29428] = 29'b0_111001011110_100_0_011100101111;
      patterns[29429] = 29'b0_111001011110_101_1_001110010111;
      patterns[29430] = 29'b0_111001011110_110_0_111001011110;
      patterns[29431] = 29'b0_111001011110_111_0_111001011110;
      patterns[29432] = 29'b0_111001011111_000_0_111001011111;
      patterns[29433] = 29'b0_111001011111_001_0_011111111001;
      patterns[29434] = 29'b0_111001011111_010_1_110010111110;
      patterns[29435] = 29'b0_111001011111_011_1_100101111101;
      patterns[29436] = 29'b0_111001011111_100_1_011100101111;
      patterns[29437] = 29'b0_111001011111_101_1_101110010111;
      patterns[29438] = 29'b0_111001011111_110_0_111001011111;
      patterns[29439] = 29'b0_111001011111_111_0_111001011111;
      patterns[29440] = 29'b0_111001100000_000_0_111001100000;
      patterns[29441] = 29'b0_111001100000_001_0_100000111001;
      patterns[29442] = 29'b0_111001100000_010_1_110011000000;
      patterns[29443] = 29'b0_111001100000_011_1_100110000001;
      patterns[29444] = 29'b0_111001100000_100_0_011100110000;
      patterns[29445] = 29'b0_111001100000_101_0_001110011000;
      patterns[29446] = 29'b0_111001100000_110_0_111001100000;
      patterns[29447] = 29'b0_111001100000_111_0_111001100000;
      patterns[29448] = 29'b0_111001100001_000_0_111001100001;
      patterns[29449] = 29'b0_111001100001_001_0_100001111001;
      patterns[29450] = 29'b0_111001100001_010_1_110011000010;
      patterns[29451] = 29'b0_111001100001_011_1_100110000101;
      patterns[29452] = 29'b0_111001100001_100_1_011100110000;
      patterns[29453] = 29'b0_111001100001_101_0_101110011000;
      patterns[29454] = 29'b0_111001100001_110_0_111001100001;
      patterns[29455] = 29'b0_111001100001_111_0_111001100001;
      patterns[29456] = 29'b0_111001100010_000_0_111001100010;
      patterns[29457] = 29'b0_111001100010_001_0_100010111001;
      patterns[29458] = 29'b0_111001100010_010_1_110011000100;
      patterns[29459] = 29'b0_111001100010_011_1_100110001001;
      patterns[29460] = 29'b0_111001100010_100_0_011100110001;
      patterns[29461] = 29'b0_111001100010_101_1_001110011000;
      patterns[29462] = 29'b0_111001100010_110_0_111001100010;
      patterns[29463] = 29'b0_111001100010_111_0_111001100010;
      patterns[29464] = 29'b0_111001100011_000_0_111001100011;
      patterns[29465] = 29'b0_111001100011_001_0_100011111001;
      patterns[29466] = 29'b0_111001100011_010_1_110011000110;
      patterns[29467] = 29'b0_111001100011_011_1_100110001101;
      patterns[29468] = 29'b0_111001100011_100_1_011100110001;
      patterns[29469] = 29'b0_111001100011_101_1_101110011000;
      patterns[29470] = 29'b0_111001100011_110_0_111001100011;
      patterns[29471] = 29'b0_111001100011_111_0_111001100011;
      patterns[29472] = 29'b0_111001100100_000_0_111001100100;
      patterns[29473] = 29'b0_111001100100_001_0_100100111001;
      patterns[29474] = 29'b0_111001100100_010_1_110011001000;
      patterns[29475] = 29'b0_111001100100_011_1_100110010001;
      patterns[29476] = 29'b0_111001100100_100_0_011100110010;
      patterns[29477] = 29'b0_111001100100_101_0_001110011001;
      patterns[29478] = 29'b0_111001100100_110_0_111001100100;
      patterns[29479] = 29'b0_111001100100_111_0_111001100100;
      patterns[29480] = 29'b0_111001100101_000_0_111001100101;
      patterns[29481] = 29'b0_111001100101_001_0_100101111001;
      patterns[29482] = 29'b0_111001100101_010_1_110011001010;
      patterns[29483] = 29'b0_111001100101_011_1_100110010101;
      patterns[29484] = 29'b0_111001100101_100_1_011100110010;
      patterns[29485] = 29'b0_111001100101_101_0_101110011001;
      patterns[29486] = 29'b0_111001100101_110_0_111001100101;
      patterns[29487] = 29'b0_111001100101_111_0_111001100101;
      patterns[29488] = 29'b0_111001100110_000_0_111001100110;
      patterns[29489] = 29'b0_111001100110_001_0_100110111001;
      patterns[29490] = 29'b0_111001100110_010_1_110011001100;
      patterns[29491] = 29'b0_111001100110_011_1_100110011001;
      patterns[29492] = 29'b0_111001100110_100_0_011100110011;
      patterns[29493] = 29'b0_111001100110_101_1_001110011001;
      patterns[29494] = 29'b0_111001100110_110_0_111001100110;
      patterns[29495] = 29'b0_111001100110_111_0_111001100110;
      patterns[29496] = 29'b0_111001100111_000_0_111001100111;
      patterns[29497] = 29'b0_111001100111_001_0_100111111001;
      patterns[29498] = 29'b0_111001100111_010_1_110011001110;
      patterns[29499] = 29'b0_111001100111_011_1_100110011101;
      patterns[29500] = 29'b0_111001100111_100_1_011100110011;
      patterns[29501] = 29'b0_111001100111_101_1_101110011001;
      patterns[29502] = 29'b0_111001100111_110_0_111001100111;
      patterns[29503] = 29'b0_111001100111_111_0_111001100111;
      patterns[29504] = 29'b0_111001101000_000_0_111001101000;
      patterns[29505] = 29'b0_111001101000_001_0_101000111001;
      patterns[29506] = 29'b0_111001101000_010_1_110011010000;
      patterns[29507] = 29'b0_111001101000_011_1_100110100001;
      patterns[29508] = 29'b0_111001101000_100_0_011100110100;
      patterns[29509] = 29'b0_111001101000_101_0_001110011010;
      patterns[29510] = 29'b0_111001101000_110_0_111001101000;
      patterns[29511] = 29'b0_111001101000_111_0_111001101000;
      patterns[29512] = 29'b0_111001101001_000_0_111001101001;
      patterns[29513] = 29'b0_111001101001_001_0_101001111001;
      patterns[29514] = 29'b0_111001101001_010_1_110011010010;
      patterns[29515] = 29'b0_111001101001_011_1_100110100101;
      patterns[29516] = 29'b0_111001101001_100_1_011100110100;
      patterns[29517] = 29'b0_111001101001_101_0_101110011010;
      patterns[29518] = 29'b0_111001101001_110_0_111001101001;
      patterns[29519] = 29'b0_111001101001_111_0_111001101001;
      patterns[29520] = 29'b0_111001101010_000_0_111001101010;
      patterns[29521] = 29'b0_111001101010_001_0_101010111001;
      patterns[29522] = 29'b0_111001101010_010_1_110011010100;
      patterns[29523] = 29'b0_111001101010_011_1_100110101001;
      patterns[29524] = 29'b0_111001101010_100_0_011100110101;
      patterns[29525] = 29'b0_111001101010_101_1_001110011010;
      patterns[29526] = 29'b0_111001101010_110_0_111001101010;
      patterns[29527] = 29'b0_111001101010_111_0_111001101010;
      patterns[29528] = 29'b0_111001101011_000_0_111001101011;
      patterns[29529] = 29'b0_111001101011_001_0_101011111001;
      patterns[29530] = 29'b0_111001101011_010_1_110011010110;
      patterns[29531] = 29'b0_111001101011_011_1_100110101101;
      patterns[29532] = 29'b0_111001101011_100_1_011100110101;
      patterns[29533] = 29'b0_111001101011_101_1_101110011010;
      patterns[29534] = 29'b0_111001101011_110_0_111001101011;
      patterns[29535] = 29'b0_111001101011_111_0_111001101011;
      patterns[29536] = 29'b0_111001101100_000_0_111001101100;
      patterns[29537] = 29'b0_111001101100_001_0_101100111001;
      patterns[29538] = 29'b0_111001101100_010_1_110011011000;
      patterns[29539] = 29'b0_111001101100_011_1_100110110001;
      patterns[29540] = 29'b0_111001101100_100_0_011100110110;
      patterns[29541] = 29'b0_111001101100_101_0_001110011011;
      patterns[29542] = 29'b0_111001101100_110_0_111001101100;
      patterns[29543] = 29'b0_111001101100_111_0_111001101100;
      patterns[29544] = 29'b0_111001101101_000_0_111001101101;
      patterns[29545] = 29'b0_111001101101_001_0_101101111001;
      patterns[29546] = 29'b0_111001101101_010_1_110011011010;
      patterns[29547] = 29'b0_111001101101_011_1_100110110101;
      patterns[29548] = 29'b0_111001101101_100_1_011100110110;
      patterns[29549] = 29'b0_111001101101_101_0_101110011011;
      patterns[29550] = 29'b0_111001101101_110_0_111001101101;
      patterns[29551] = 29'b0_111001101101_111_0_111001101101;
      patterns[29552] = 29'b0_111001101110_000_0_111001101110;
      patterns[29553] = 29'b0_111001101110_001_0_101110111001;
      patterns[29554] = 29'b0_111001101110_010_1_110011011100;
      patterns[29555] = 29'b0_111001101110_011_1_100110111001;
      patterns[29556] = 29'b0_111001101110_100_0_011100110111;
      patterns[29557] = 29'b0_111001101110_101_1_001110011011;
      patterns[29558] = 29'b0_111001101110_110_0_111001101110;
      patterns[29559] = 29'b0_111001101110_111_0_111001101110;
      patterns[29560] = 29'b0_111001101111_000_0_111001101111;
      patterns[29561] = 29'b0_111001101111_001_0_101111111001;
      patterns[29562] = 29'b0_111001101111_010_1_110011011110;
      patterns[29563] = 29'b0_111001101111_011_1_100110111101;
      patterns[29564] = 29'b0_111001101111_100_1_011100110111;
      patterns[29565] = 29'b0_111001101111_101_1_101110011011;
      patterns[29566] = 29'b0_111001101111_110_0_111001101111;
      patterns[29567] = 29'b0_111001101111_111_0_111001101111;
      patterns[29568] = 29'b0_111001110000_000_0_111001110000;
      patterns[29569] = 29'b0_111001110000_001_0_110000111001;
      patterns[29570] = 29'b0_111001110000_010_1_110011100000;
      patterns[29571] = 29'b0_111001110000_011_1_100111000001;
      patterns[29572] = 29'b0_111001110000_100_0_011100111000;
      patterns[29573] = 29'b0_111001110000_101_0_001110011100;
      patterns[29574] = 29'b0_111001110000_110_0_111001110000;
      patterns[29575] = 29'b0_111001110000_111_0_111001110000;
      patterns[29576] = 29'b0_111001110001_000_0_111001110001;
      patterns[29577] = 29'b0_111001110001_001_0_110001111001;
      patterns[29578] = 29'b0_111001110001_010_1_110011100010;
      patterns[29579] = 29'b0_111001110001_011_1_100111000101;
      patterns[29580] = 29'b0_111001110001_100_1_011100111000;
      patterns[29581] = 29'b0_111001110001_101_0_101110011100;
      patterns[29582] = 29'b0_111001110001_110_0_111001110001;
      patterns[29583] = 29'b0_111001110001_111_0_111001110001;
      patterns[29584] = 29'b0_111001110010_000_0_111001110010;
      patterns[29585] = 29'b0_111001110010_001_0_110010111001;
      patterns[29586] = 29'b0_111001110010_010_1_110011100100;
      patterns[29587] = 29'b0_111001110010_011_1_100111001001;
      patterns[29588] = 29'b0_111001110010_100_0_011100111001;
      patterns[29589] = 29'b0_111001110010_101_1_001110011100;
      patterns[29590] = 29'b0_111001110010_110_0_111001110010;
      patterns[29591] = 29'b0_111001110010_111_0_111001110010;
      patterns[29592] = 29'b0_111001110011_000_0_111001110011;
      patterns[29593] = 29'b0_111001110011_001_0_110011111001;
      patterns[29594] = 29'b0_111001110011_010_1_110011100110;
      patterns[29595] = 29'b0_111001110011_011_1_100111001101;
      patterns[29596] = 29'b0_111001110011_100_1_011100111001;
      patterns[29597] = 29'b0_111001110011_101_1_101110011100;
      patterns[29598] = 29'b0_111001110011_110_0_111001110011;
      patterns[29599] = 29'b0_111001110011_111_0_111001110011;
      patterns[29600] = 29'b0_111001110100_000_0_111001110100;
      patterns[29601] = 29'b0_111001110100_001_0_110100111001;
      patterns[29602] = 29'b0_111001110100_010_1_110011101000;
      patterns[29603] = 29'b0_111001110100_011_1_100111010001;
      patterns[29604] = 29'b0_111001110100_100_0_011100111010;
      patterns[29605] = 29'b0_111001110100_101_0_001110011101;
      patterns[29606] = 29'b0_111001110100_110_0_111001110100;
      patterns[29607] = 29'b0_111001110100_111_0_111001110100;
      patterns[29608] = 29'b0_111001110101_000_0_111001110101;
      patterns[29609] = 29'b0_111001110101_001_0_110101111001;
      patterns[29610] = 29'b0_111001110101_010_1_110011101010;
      patterns[29611] = 29'b0_111001110101_011_1_100111010101;
      patterns[29612] = 29'b0_111001110101_100_1_011100111010;
      patterns[29613] = 29'b0_111001110101_101_0_101110011101;
      patterns[29614] = 29'b0_111001110101_110_0_111001110101;
      patterns[29615] = 29'b0_111001110101_111_0_111001110101;
      patterns[29616] = 29'b0_111001110110_000_0_111001110110;
      patterns[29617] = 29'b0_111001110110_001_0_110110111001;
      patterns[29618] = 29'b0_111001110110_010_1_110011101100;
      patterns[29619] = 29'b0_111001110110_011_1_100111011001;
      patterns[29620] = 29'b0_111001110110_100_0_011100111011;
      patterns[29621] = 29'b0_111001110110_101_1_001110011101;
      patterns[29622] = 29'b0_111001110110_110_0_111001110110;
      patterns[29623] = 29'b0_111001110110_111_0_111001110110;
      patterns[29624] = 29'b0_111001110111_000_0_111001110111;
      patterns[29625] = 29'b0_111001110111_001_0_110111111001;
      patterns[29626] = 29'b0_111001110111_010_1_110011101110;
      patterns[29627] = 29'b0_111001110111_011_1_100111011101;
      patterns[29628] = 29'b0_111001110111_100_1_011100111011;
      patterns[29629] = 29'b0_111001110111_101_1_101110011101;
      patterns[29630] = 29'b0_111001110111_110_0_111001110111;
      patterns[29631] = 29'b0_111001110111_111_0_111001110111;
      patterns[29632] = 29'b0_111001111000_000_0_111001111000;
      patterns[29633] = 29'b0_111001111000_001_0_111000111001;
      patterns[29634] = 29'b0_111001111000_010_1_110011110000;
      patterns[29635] = 29'b0_111001111000_011_1_100111100001;
      patterns[29636] = 29'b0_111001111000_100_0_011100111100;
      patterns[29637] = 29'b0_111001111000_101_0_001110011110;
      patterns[29638] = 29'b0_111001111000_110_0_111001111000;
      patterns[29639] = 29'b0_111001111000_111_0_111001111000;
      patterns[29640] = 29'b0_111001111001_000_0_111001111001;
      patterns[29641] = 29'b0_111001111001_001_0_111001111001;
      patterns[29642] = 29'b0_111001111001_010_1_110011110010;
      patterns[29643] = 29'b0_111001111001_011_1_100111100101;
      patterns[29644] = 29'b0_111001111001_100_1_011100111100;
      patterns[29645] = 29'b0_111001111001_101_0_101110011110;
      patterns[29646] = 29'b0_111001111001_110_0_111001111001;
      patterns[29647] = 29'b0_111001111001_111_0_111001111001;
      patterns[29648] = 29'b0_111001111010_000_0_111001111010;
      patterns[29649] = 29'b0_111001111010_001_0_111010111001;
      patterns[29650] = 29'b0_111001111010_010_1_110011110100;
      patterns[29651] = 29'b0_111001111010_011_1_100111101001;
      patterns[29652] = 29'b0_111001111010_100_0_011100111101;
      patterns[29653] = 29'b0_111001111010_101_1_001110011110;
      patterns[29654] = 29'b0_111001111010_110_0_111001111010;
      patterns[29655] = 29'b0_111001111010_111_0_111001111010;
      patterns[29656] = 29'b0_111001111011_000_0_111001111011;
      patterns[29657] = 29'b0_111001111011_001_0_111011111001;
      patterns[29658] = 29'b0_111001111011_010_1_110011110110;
      patterns[29659] = 29'b0_111001111011_011_1_100111101101;
      patterns[29660] = 29'b0_111001111011_100_1_011100111101;
      patterns[29661] = 29'b0_111001111011_101_1_101110011110;
      patterns[29662] = 29'b0_111001111011_110_0_111001111011;
      patterns[29663] = 29'b0_111001111011_111_0_111001111011;
      patterns[29664] = 29'b0_111001111100_000_0_111001111100;
      patterns[29665] = 29'b0_111001111100_001_0_111100111001;
      patterns[29666] = 29'b0_111001111100_010_1_110011111000;
      patterns[29667] = 29'b0_111001111100_011_1_100111110001;
      patterns[29668] = 29'b0_111001111100_100_0_011100111110;
      patterns[29669] = 29'b0_111001111100_101_0_001110011111;
      patterns[29670] = 29'b0_111001111100_110_0_111001111100;
      patterns[29671] = 29'b0_111001111100_111_0_111001111100;
      patterns[29672] = 29'b0_111001111101_000_0_111001111101;
      patterns[29673] = 29'b0_111001111101_001_0_111101111001;
      patterns[29674] = 29'b0_111001111101_010_1_110011111010;
      patterns[29675] = 29'b0_111001111101_011_1_100111110101;
      patterns[29676] = 29'b0_111001111101_100_1_011100111110;
      patterns[29677] = 29'b0_111001111101_101_0_101110011111;
      patterns[29678] = 29'b0_111001111101_110_0_111001111101;
      patterns[29679] = 29'b0_111001111101_111_0_111001111101;
      patterns[29680] = 29'b0_111001111110_000_0_111001111110;
      patterns[29681] = 29'b0_111001111110_001_0_111110111001;
      patterns[29682] = 29'b0_111001111110_010_1_110011111100;
      patterns[29683] = 29'b0_111001111110_011_1_100111111001;
      patterns[29684] = 29'b0_111001111110_100_0_011100111111;
      patterns[29685] = 29'b0_111001111110_101_1_001110011111;
      patterns[29686] = 29'b0_111001111110_110_0_111001111110;
      patterns[29687] = 29'b0_111001111110_111_0_111001111110;
      patterns[29688] = 29'b0_111001111111_000_0_111001111111;
      patterns[29689] = 29'b0_111001111111_001_0_111111111001;
      patterns[29690] = 29'b0_111001111111_010_1_110011111110;
      patterns[29691] = 29'b0_111001111111_011_1_100111111101;
      patterns[29692] = 29'b0_111001111111_100_1_011100111111;
      patterns[29693] = 29'b0_111001111111_101_1_101110011111;
      patterns[29694] = 29'b0_111001111111_110_0_111001111111;
      patterns[29695] = 29'b0_111001111111_111_0_111001111111;
      patterns[29696] = 29'b0_111010000000_000_0_111010000000;
      patterns[29697] = 29'b0_111010000000_001_0_000000111010;
      patterns[29698] = 29'b0_111010000000_010_1_110100000000;
      patterns[29699] = 29'b0_111010000000_011_1_101000000001;
      patterns[29700] = 29'b0_111010000000_100_0_011101000000;
      patterns[29701] = 29'b0_111010000000_101_0_001110100000;
      patterns[29702] = 29'b0_111010000000_110_0_111010000000;
      patterns[29703] = 29'b0_111010000000_111_0_111010000000;
      patterns[29704] = 29'b0_111010000001_000_0_111010000001;
      patterns[29705] = 29'b0_111010000001_001_0_000001111010;
      patterns[29706] = 29'b0_111010000001_010_1_110100000010;
      patterns[29707] = 29'b0_111010000001_011_1_101000000101;
      patterns[29708] = 29'b0_111010000001_100_1_011101000000;
      patterns[29709] = 29'b0_111010000001_101_0_101110100000;
      patterns[29710] = 29'b0_111010000001_110_0_111010000001;
      patterns[29711] = 29'b0_111010000001_111_0_111010000001;
      patterns[29712] = 29'b0_111010000010_000_0_111010000010;
      patterns[29713] = 29'b0_111010000010_001_0_000010111010;
      patterns[29714] = 29'b0_111010000010_010_1_110100000100;
      patterns[29715] = 29'b0_111010000010_011_1_101000001001;
      patterns[29716] = 29'b0_111010000010_100_0_011101000001;
      patterns[29717] = 29'b0_111010000010_101_1_001110100000;
      patterns[29718] = 29'b0_111010000010_110_0_111010000010;
      patterns[29719] = 29'b0_111010000010_111_0_111010000010;
      patterns[29720] = 29'b0_111010000011_000_0_111010000011;
      patterns[29721] = 29'b0_111010000011_001_0_000011111010;
      patterns[29722] = 29'b0_111010000011_010_1_110100000110;
      patterns[29723] = 29'b0_111010000011_011_1_101000001101;
      patterns[29724] = 29'b0_111010000011_100_1_011101000001;
      patterns[29725] = 29'b0_111010000011_101_1_101110100000;
      patterns[29726] = 29'b0_111010000011_110_0_111010000011;
      patterns[29727] = 29'b0_111010000011_111_0_111010000011;
      patterns[29728] = 29'b0_111010000100_000_0_111010000100;
      patterns[29729] = 29'b0_111010000100_001_0_000100111010;
      patterns[29730] = 29'b0_111010000100_010_1_110100001000;
      patterns[29731] = 29'b0_111010000100_011_1_101000010001;
      patterns[29732] = 29'b0_111010000100_100_0_011101000010;
      patterns[29733] = 29'b0_111010000100_101_0_001110100001;
      patterns[29734] = 29'b0_111010000100_110_0_111010000100;
      patterns[29735] = 29'b0_111010000100_111_0_111010000100;
      patterns[29736] = 29'b0_111010000101_000_0_111010000101;
      patterns[29737] = 29'b0_111010000101_001_0_000101111010;
      patterns[29738] = 29'b0_111010000101_010_1_110100001010;
      patterns[29739] = 29'b0_111010000101_011_1_101000010101;
      patterns[29740] = 29'b0_111010000101_100_1_011101000010;
      patterns[29741] = 29'b0_111010000101_101_0_101110100001;
      patterns[29742] = 29'b0_111010000101_110_0_111010000101;
      patterns[29743] = 29'b0_111010000101_111_0_111010000101;
      patterns[29744] = 29'b0_111010000110_000_0_111010000110;
      patterns[29745] = 29'b0_111010000110_001_0_000110111010;
      patterns[29746] = 29'b0_111010000110_010_1_110100001100;
      patterns[29747] = 29'b0_111010000110_011_1_101000011001;
      patterns[29748] = 29'b0_111010000110_100_0_011101000011;
      patterns[29749] = 29'b0_111010000110_101_1_001110100001;
      patterns[29750] = 29'b0_111010000110_110_0_111010000110;
      patterns[29751] = 29'b0_111010000110_111_0_111010000110;
      patterns[29752] = 29'b0_111010000111_000_0_111010000111;
      patterns[29753] = 29'b0_111010000111_001_0_000111111010;
      patterns[29754] = 29'b0_111010000111_010_1_110100001110;
      patterns[29755] = 29'b0_111010000111_011_1_101000011101;
      patterns[29756] = 29'b0_111010000111_100_1_011101000011;
      patterns[29757] = 29'b0_111010000111_101_1_101110100001;
      patterns[29758] = 29'b0_111010000111_110_0_111010000111;
      patterns[29759] = 29'b0_111010000111_111_0_111010000111;
      patterns[29760] = 29'b0_111010001000_000_0_111010001000;
      patterns[29761] = 29'b0_111010001000_001_0_001000111010;
      patterns[29762] = 29'b0_111010001000_010_1_110100010000;
      patterns[29763] = 29'b0_111010001000_011_1_101000100001;
      patterns[29764] = 29'b0_111010001000_100_0_011101000100;
      patterns[29765] = 29'b0_111010001000_101_0_001110100010;
      patterns[29766] = 29'b0_111010001000_110_0_111010001000;
      patterns[29767] = 29'b0_111010001000_111_0_111010001000;
      patterns[29768] = 29'b0_111010001001_000_0_111010001001;
      patterns[29769] = 29'b0_111010001001_001_0_001001111010;
      patterns[29770] = 29'b0_111010001001_010_1_110100010010;
      patterns[29771] = 29'b0_111010001001_011_1_101000100101;
      patterns[29772] = 29'b0_111010001001_100_1_011101000100;
      patterns[29773] = 29'b0_111010001001_101_0_101110100010;
      patterns[29774] = 29'b0_111010001001_110_0_111010001001;
      patterns[29775] = 29'b0_111010001001_111_0_111010001001;
      patterns[29776] = 29'b0_111010001010_000_0_111010001010;
      patterns[29777] = 29'b0_111010001010_001_0_001010111010;
      patterns[29778] = 29'b0_111010001010_010_1_110100010100;
      patterns[29779] = 29'b0_111010001010_011_1_101000101001;
      patterns[29780] = 29'b0_111010001010_100_0_011101000101;
      patterns[29781] = 29'b0_111010001010_101_1_001110100010;
      patterns[29782] = 29'b0_111010001010_110_0_111010001010;
      patterns[29783] = 29'b0_111010001010_111_0_111010001010;
      patterns[29784] = 29'b0_111010001011_000_0_111010001011;
      patterns[29785] = 29'b0_111010001011_001_0_001011111010;
      patterns[29786] = 29'b0_111010001011_010_1_110100010110;
      patterns[29787] = 29'b0_111010001011_011_1_101000101101;
      patterns[29788] = 29'b0_111010001011_100_1_011101000101;
      patterns[29789] = 29'b0_111010001011_101_1_101110100010;
      patterns[29790] = 29'b0_111010001011_110_0_111010001011;
      patterns[29791] = 29'b0_111010001011_111_0_111010001011;
      patterns[29792] = 29'b0_111010001100_000_0_111010001100;
      patterns[29793] = 29'b0_111010001100_001_0_001100111010;
      patterns[29794] = 29'b0_111010001100_010_1_110100011000;
      patterns[29795] = 29'b0_111010001100_011_1_101000110001;
      patterns[29796] = 29'b0_111010001100_100_0_011101000110;
      patterns[29797] = 29'b0_111010001100_101_0_001110100011;
      patterns[29798] = 29'b0_111010001100_110_0_111010001100;
      patterns[29799] = 29'b0_111010001100_111_0_111010001100;
      patterns[29800] = 29'b0_111010001101_000_0_111010001101;
      patterns[29801] = 29'b0_111010001101_001_0_001101111010;
      patterns[29802] = 29'b0_111010001101_010_1_110100011010;
      patterns[29803] = 29'b0_111010001101_011_1_101000110101;
      patterns[29804] = 29'b0_111010001101_100_1_011101000110;
      patterns[29805] = 29'b0_111010001101_101_0_101110100011;
      patterns[29806] = 29'b0_111010001101_110_0_111010001101;
      patterns[29807] = 29'b0_111010001101_111_0_111010001101;
      patterns[29808] = 29'b0_111010001110_000_0_111010001110;
      patterns[29809] = 29'b0_111010001110_001_0_001110111010;
      patterns[29810] = 29'b0_111010001110_010_1_110100011100;
      patterns[29811] = 29'b0_111010001110_011_1_101000111001;
      patterns[29812] = 29'b0_111010001110_100_0_011101000111;
      patterns[29813] = 29'b0_111010001110_101_1_001110100011;
      patterns[29814] = 29'b0_111010001110_110_0_111010001110;
      patterns[29815] = 29'b0_111010001110_111_0_111010001110;
      patterns[29816] = 29'b0_111010001111_000_0_111010001111;
      patterns[29817] = 29'b0_111010001111_001_0_001111111010;
      patterns[29818] = 29'b0_111010001111_010_1_110100011110;
      patterns[29819] = 29'b0_111010001111_011_1_101000111101;
      patterns[29820] = 29'b0_111010001111_100_1_011101000111;
      patterns[29821] = 29'b0_111010001111_101_1_101110100011;
      patterns[29822] = 29'b0_111010001111_110_0_111010001111;
      patterns[29823] = 29'b0_111010001111_111_0_111010001111;
      patterns[29824] = 29'b0_111010010000_000_0_111010010000;
      patterns[29825] = 29'b0_111010010000_001_0_010000111010;
      patterns[29826] = 29'b0_111010010000_010_1_110100100000;
      patterns[29827] = 29'b0_111010010000_011_1_101001000001;
      patterns[29828] = 29'b0_111010010000_100_0_011101001000;
      patterns[29829] = 29'b0_111010010000_101_0_001110100100;
      patterns[29830] = 29'b0_111010010000_110_0_111010010000;
      patterns[29831] = 29'b0_111010010000_111_0_111010010000;
      patterns[29832] = 29'b0_111010010001_000_0_111010010001;
      patterns[29833] = 29'b0_111010010001_001_0_010001111010;
      patterns[29834] = 29'b0_111010010001_010_1_110100100010;
      patterns[29835] = 29'b0_111010010001_011_1_101001000101;
      patterns[29836] = 29'b0_111010010001_100_1_011101001000;
      patterns[29837] = 29'b0_111010010001_101_0_101110100100;
      patterns[29838] = 29'b0_111010010001_110_0_111010010001;
      patterns[29839] = 29'b0_111010010001_111_0_111010010001;
      patterns[29840] = 29'b0_111010010010_000_0_111010010010;
      patterns[29841] = 29'b0_111010010010_001_0_010010111010;
      patterns[29842] = 29'b0_111010010010_010_1_110100100100;
      patterns[29843] = 29'b0_111010010010_011_1_101001001001;
      patterns[29844] = 29'b0_111010010010_100_0_011101001001;
      patterns[29845] = 29'b0_111010010010_101_1_001110100100;
      patterns[29846] = 29'b0_111010010010_110_0_111010010010;
      patterns[29847] = 29'b0_111010010010_111_0_111010010010;
      patterns[29848] = 29'b0_111010010011_000_0_111010010011;
      patterns[29849] = 29'b0_111010010011_001_0_010011111010;
      patterns[29850] = 29'b0_111010010011_010_1_110100100110;
      patterns[29851] = 29'b0_111010010011_011_1_101001001101;
      patterns[29852] = 29'b0_111010010011_100_1_011101001001;
      patterns[29853] = 29'b0_111010010011_101_1_101110100100;
      patterns[29854] = 29'b0_111010010011_110_0_111010010011;
      patterns[29855] = 29'b0_111010010011_111_0_111010010011;
      patterns[29856] = 29'b0_111010010100_000_0_111010010100;
      patterns[29857] = 29'b0_111010010100_001_0_010100111010;
      patterns[29858] = 29'b0_111010010100_010_1_110100101000;
      patterns[29859] = 29'b0_111010010100_011_1_101001010001;
      patterns[29860] = 29'b0_111010010100_100_0_011101001010;
      patterns[29861] = 29'b0_111010010100_101_0_001110100101;
      patterns[29862] = 29'b0_111010010100_110_0_111010010100;
      patterns[29863] = 29'b0_111010010100_111_0_111010010100;
      patterns[29864] = 29'b0_111010010101_000_0_111010010101;
      patterns[29865] = 29'b0_111010010101_001_0_010101111010;
      patterns[29866] = 29'b0_111010010101_010_1_110100101010;
      patterns[29867] = 29'b0_111010010101_011_1_101001010101;
      patterns[29868] = 29'b0_111010010101_100_1_011101001010;
      patterns[29869] = 29'b0_111010010101_101_0_101110100101;
      patterns[29870] = 29'b0_111010010101_110_0_111010010101;
      patterns[29871] = 29'b0_111010010101_111_0_111010010101;
      patterns[29872] = 29'b0_111010010110_000_0_111010010110;
      patterns[29873] = 29'b0_111010010110_001_0_010110111010;
      patterns[29874] = 29'b0_111010010110_010_1_110100101100;
      patterns[29875] = 29'b0_111010010110_011_1_101001011001;
      patterns[29876] = 29'b0_111010010110_100_0_011101001011;
      patterns[29877] = 29'b0_111010010110_101_1_001110100101;
      patterns[29878] = 29'b0_111010010110_110_0_111010010110;
      patterns[29879] = 29'b0_111010010110_111_0_111010010110;
      patterns[29880] = 29'b0_111010010111_000_0_111010010111;
      patterns[29881] = 29'b0_111010010111_001_0_010111111010;
      patterns[29882] = 29'b0_111010010111_010_1_110100101110;
      patterns[29883] = 29'b0_111010010111_011_1_101001011101;
      patterns[29884] = 29'b0_111010010111_100_1_011101001011;
      patterns[29885] = 29'b0_111010010111_101_1_101110100101;
      patterns[29886] = 29'b0_111010010111_110_0_111010010111;
      patterns[29887] = 29'b0_111010010111_111_0_111010010111;
      patterns[29888] = 29'b0_111010011000_000_0_111010011000;
      patterns[29889] = 29'b0_111010011000_001_0_011000111010;
      patterns[29890] = 29'b0_111010011000_010_1_110100110000;
      patterns[29891] = 29'b0_111010011000_011_1_101001100001;
      patterns[29892] = 29'b0_111010011000_100_0_011101001100;
      patterns[29893] = 29'b0_111010011000_101_0_001110100110;
      patterns[29894] = 29'b0_111010011000_110_0_111010011000;
      patterns[29895] = 29'b0_111010011000_111_0_111010011000;
      patterns[29896] = 29'b0_111010011001_000_0_111010011001;
      patterns[29897] = 29'b0_111010011001_001_0_011001111010;
      patterns[29898] = 29'b0_111010011001_010_1_110100110010;
      patterns[29899] = 29'b0_111010011001_011_1_101001100101;
      patterns[29900] = 29'b0_111010011001_100_1_011101001100;
      patterns[29901] = 29'b0_111010011001_101_0_101110100110;
      patterns[29902] = 29'b0_111010011001_110_0_111010011001;
      patterns[29903] = 29'b0_111010011001_111_0_111010011001;
      patterns[29904] = 29'b0_111010011010_000_0_111010011010;
      patterns[29905] = 29'b0_111010011010_001_0_011010111010;
      patterns[29906] = 29'b0_111010011010_010_1_110100110100;
      patterns[29907] = 29'b0_111010011010_011_1_101001101001;
      patterns[29908] = 29'b0_111010011010_100_0_011101001101;
      patterns[29909] = 29'b0_111010011010_101_1_001110100110;
      patterns[29910] = 29'b0_111010011010_110_0_111010011010;
      patterns[29911] = 29'b0_111010011010_111_0_111010011010;
      patterns[29912] = 29'b0_111010011011_000_0_111010011011;
      patterns[29913] = 29'b0_111010011011_001_0_011011111010;
      patterns[29914] = 29'b0_111010011011_010_1_110100110110;
      patterns[29915] = 29'b0_111010011011_011_1_101001101101;
      patterns[29916] = 29'b0_111010011011_100_1_011101001101;
      patterns[29917] = 29'b0_111010011011_101_1_101110100110;
      patterns[29918] = 29'b0_111010011011_110_0_111010011011;
      patterns[29919] = 29'b0_111010011011_111_0_111010011011;
      patterns[29920] = 29'b0_111010011100_000_0_111010011100;
      patterns[29921] = 29'b0_111010011100_001_0_011100111010;
      patterns[29922] = 29'b0_111010011100_010_1_110100111000;
      patterns[29923] = 29'b0_111010011100_011_1_101001110001;
      patterns[29924] = 29'b0_111010011100_100_0_011101001110;
      patterns[29925] = 29'b0_111010011100_101_0_001110100111;
      patterns[29926] = 29'b0_111010011100_110_0_111010011100;
      patterns[29927] = 29'b0_111010011100_111_0_111010011100;
      patterns[29928] = 29'b0_111010011101_000_0_111010011101;
      patterns[29929] = 29'b0_111010011101_001_0_011101111010;
      patterns[29930] = 29'b0_111010011101_010_1_110100111010;
      patterns[29931] = 29'b0_111010011101_011_1_101001110101;
      patterns[29932] = 29'b0_111010011101_100_1_011101001110;
      patterns[29933] = 29'b0_111010011101_101_0_101110100111;
      patterns[29934] = 29'b0_111010011101_110_0_111010011101;
      patterns[29935] = 29'b0_111010011101_111_0_111010011101;
      patterns[29936] = 29'b0_111010011110_000_0_111010011110;
      patterns[29937] = 29'b0_111010011110_001_0_011110111010;
      patterns[29938] = 29'b0_111010011110_010_1_110100111100;
      patterns[29939] = 29'b0_111010011110_011_1_101001111001;
      patterns[29940] = 29'b0_111010011110_100_0_011101001111;
      patterns[29941] = 29'b0_111010011110_101_1_001110100111;
      patterns[29942] = 29'b0_111010011110_110_0_111010011110;
      patterns[29943] = 29'b0_111010011110_111_0_111010011110;
      patterns[29944] = 29'b0_111010011111_000_0_111010011111;
      patterns[29945] = 29'b0_111010011111_001_0_011111111010;
      patterns[29946] = 29'b0_111010011111_010_1_110100111110;
      patterns[29947] = 29'b0_111010011111_011_1_101001111101;
      patterns[29948] = 29'b0_111010011111_100_1_011101001111;
      patterns[29949] = 29'b0_111010011111_101_1_101110100111;
      patterns[29950] = 29'b0_111010011111_110_0_111010011111;
      patterns[29951] = 29'b0_111010011111_111_0_111010011111;
      patterns[29952] = 29'b0_111010100000_000_0_111010100000;
      patterns[29953] = 29'b0_111010100000_001_0_100000111010;
      patterns[29954] = 29'b0_111010100000_010_1_110101000000;
      patterns[29955] = 29'b0_111010100000_011_1_101010000001;
      patterns[29956] = 29'b0_111010100000_100_0_011101010000;
      patterns[29957] = 29'b0_111010100000_101_0_001110101000;
      patterns[29958] = 29'b0_111010100000_110_0_111010100000;
      patterns[29959] = 29'b0_111010100000_111_0_111010100000;
      patterns[29960] = 29'b0_111010100001_000_0_111010100001;
      patterns[29961] = 29'b0_111010100001_001_0_100001111010;
      patterns[29962] = 29'b0_111010100001_010_1_110101000010;
      patterns[29963] = 29'b0_111010100001_011_1_101010000101;
      patterns[29964] = 29'b0_111010100001_100_1_011101010000;
      patterns[29965] = 29'b0_111010100001_101_0_101110101000;
      patterns[29966] = 29'b0_111010100001_110_0_111010100001;
      patterns[29967] = 29'b0_111010100001_111_0_111010100001;
      patterns[29968] = 29'b0_111010100010_000_0_111010100010;
      patterns[29969] = 29'b0_111010100010_001_0_100010111010;
      patterns[29970] = 29'b0_111010100010_010_1_110101000100;
      patterns[29971] = 29'b0_111010100010_011_1_101010001001;
      patterns[29972] = 29'b0_111010100010_100_0_011101010001;
      patterns[29973] = 29'b0_111010100010_101_1_001110101000;
      patterns[29974] = 29'b0_111010100010_110_0_111010100010;
      patterns[29975] = 29'b0_111010100010_111_0_111010100010;
      patterns[29976] = 29'b0_111010100011_000_0_111010100011;
      patterns[29977] = 29'b0_111010100011_001_0_100011111010;
      patterns[29978] = 29'b0_111010100011_010_1_110101000110;
      patterns[29979] = 29'b0_111010100011_011_1_101010001101;
      patterns[29980] = 29'b0_111010100011_100_1_011101010001;
      patterns[29981] = 29'b0_111010100011_101_1_101110101000;
      patterns[29982] = 29'b0_111010100011_110_0_111010100011;
      patterns[29983] = 29'b0_111010100011_111_0_111010100011;
      patterns[29984] = 29'b0_111010100100_000_0_111010100100;
      patterns[29985] = 29'b0_111010100100_001_0_100100111010;
      patterns[29986] = 29'b0_111010100100_010_1_110101001000;
      patterns[29987] = 29'b0_111010100100_011_1_101010010001;
      patterns[29988] = 29'b0_111010100100_100_0_011101010010;
      patterns[29989] = 29'b0_111010100100_101_0_001110101001;
      patterns[29990] = 29'b0_111010100100_110_0_111010100100;
      patterns[29991] = 29'b0_111010100100_111_0_111010100100;
      patterns[29992] = 29'b0_111010100101_000_0_111010100101;
      patterns[29993] = 29'b0_111010100101_001_0_100101111010;
      patterns[29994] = 29'b0_111010100101_010_1_110101001010;
      patterns[29995] = 29'b0_111010100101_011_1_101010010101;
      patterns[29996] = 29'b0_111010100101_100_1_011101010010;
      patterns[29997] = 29'b0_111010100101_101_0_101110101001;
      patterns[29998] = 29'b0_111010100101_110_0_111010100101;
      patterns[29999] = 29'b0_111010100101_111_0_111010100101;
      patterns[30000] = 29'b0_111010100110_000_0_111010100110;
      patterns[30001] = 29'b0_111010100110_001_0_100110111010;
      patterns[30002] = 29'b0_111010100110_010_1_110101001100;
      patterns[30003] = 29'b0_111010100110_011_1_101010011001;
      patterns[30004] = 29'b0_111010100110_100_0_011101010011;
      patterns[30005] = 29'b0_111010100110_101_1_001110101001;
      patterns[30006] = 29'b0_111010100110_110_0_111010100110;
      patterns[30007] = 29'b0_111010100110_111_0_111010100110;
      patterns[30008] = 29'b0_111010100111_000_0_111010100111;
      patterns[30009] = 29'b0_111010100111_001_0_100111111010;
      patterns[30010] = 29'b0_111010100111_010_1_110101001110;
      patterns[30011] = 29'b0_111010100111_011_1_101010011101;
      patterns[30012] = 29'b0_111010100111_100_1_011101010011;
      patterns[30013] = 29'b0_111010100111_101_1_101110101001;
      patterns[30014] = 29'b0_111010100111_110_0_111010100111;
      patterns[30015] = 29'b0_111010100111_111_0_111010100111;
      patterns[30016] = 29'b0_111010101000_000_0_111010101000;
      patterns[30017] = 29'b0_111010101000_001_0_101000111010;
      patterns[30018] = 29'b0_111010101000_010_1_110101010000;
      patterns[30019] = 29'b0_111010101000_011_1_101010100001;
      patterns[30020] = 29'b0_111010101000_100_0_011101010100;
      patterns[30021] = 29'b0_111010101000_101_0_001110101010;
      patterns[30022] = 29'b0_111010101000_110_0_111010101000;
      patterns[30023] = 29'b0_111010101000_111_0_111010101000;
      patterns[30024] = 29'b0_111010101001_000_0_111010101001;
      patterns[30025] = 29'b0_111010101001_001_0_101001111010;
      patterns[30026] = 29'b0_111010101001_010_1_110101010010;
      patterns[30027] = 29'b0_111010101001_011_1_101010100101;
      patterns[30028] = 29'b0_111010101001_100_1_011101010100;
      patterns[30029] = 29'b0_111010101001_101_0_101110101010;
      patterns[30030] = 29'b0_111010101001_110_0_111010101001;
      patterns[30031] = 29'b0_111010101001_111_0_111010101001;
      patterns[30032] = 29'b0_111010101010_000_0_111010101010;
      patterns[30033] = 29'b0_111010101010_001_0_101010111010;
      patterns[30034] = 29'b0_111010101010_010_1_110101010100;
      patterns[30035] = 29'b0_111010101010_011_1_101010101001;
      patterns[30036] = 29'b0_111010101010_100_0_011101010101;
      patterns[30037] = 29'b0_111010101010_101_1_001110101010;
      patterns[30038] = 29'b0_111010101010_110_0_111010101010;
      patterns[30039] = 29'b0_111010101010_111_0_111010101010;
      patterns[30040] = 29'b0_111010101011_000_0_111010101011;
      patterns[30041] = 29'b0_111010101011_001_0_101011111010;
      patterns[30042] = 29'b0_111010101011_010_1_110101010110;
      patterns[30043] = 29'b0_111010101011_011_1_101010101101;
      patterns[30044] = 29'b0_111010101011_100_1_011101010101;
      patterns[30045] = 29'b0_111010101011_101_1_101110101010;
      patterns[30046] = 29'b0_111010101011_110_0_111010101011;
      patterns[30047] = 29'b0_111010101011_111_0_111010101011;
      patterns[30048] = 29'b0_111010101100_000_0_111010101100;
      patterns[30049] = 29'b0_111010101100_001_0_101100111010;
      patterns[30050] = 29'b0_111010101100_010_1_110101011000;
      patterns[30051] = 29'b0_111010101100_011_1_101010110001;
      patterns[30052] = 29'b0_111010101100_100_0_011101010110;
      patterns[30053] = 29'b0_111010101100_101_0_001110101011;
      patterns[30054] = 29'b0_111010101100_110_0_111010101100;
      patterns[30055] = 29'b0_111010101100_111_0_111010101100;
      patterns[30056] = 29'b0_111010101101_000_0_111010101101;
      patterns[30057] = 29'b0_111010101101_001_0_101101111010;
      patterns[30058] = 29'b0_111010101101_010_1_110101011010;
      patterns[30059] = 29'b0_111010101101_011_1_101010110101;
      patterns[30060] = 29'b0_111010101101_100_1_011101010110;
      patterns[30061] = 29'b0_111010101101_101_0_101110101011;
      patterns[30062] = 29'b0_111010101101_110_0_111010101101;
      patterns[30063] = 29'b0_111010101101_111_0_111010101101;
      patterns[30064] = 29'b0_111010101110_000_0_111010101110;
      patterns[30065] = 29'b0_111010101110_001_0_101110111010;
      patterns[30066] = 29'b0_111010101110_010_1_110101011100;
      patterns[30067] = 29'b0_111010101110_011_1_101010111001;
      patterns[30068] = 29'b0_111010101110_100_0_011101010111;
      patterns[30069] = 29'b0_111010101110_101_1_001110101011;
      patterns[30070] = 29'b0_111010101110_110_0_111010101110;
      patterns[30071] = 29'b0_111010101110_111_0_111010101110;
      patterns[30072] = 29'b0_111010101111_000_0_111010101111;
      patterns[30073] = 29'b0_111010101111_001_0_101111111010;
      patterns[30074] = 29'b0_111010101111_010_1_110101011110;
      patterns[30075] = 29'b0_111010101111_011_1_101010111101;
      patterns[30076] = 29'b0_111010101111_100_1_011101010111;
      patterns[30077] = 29'b0_111010101111_101_1_101110101011;
      patterns[30078] = 29'b0_111010101111_110_0_111010101111;
      patterns[30079] = 29'b0_111010101111_111_0_111010101111;
      patterns[30080] = 29'b0_111010110000_000_0_111010110000;
      patterns[30081] = 29'b0_111010110000_001_0_110000111010;
      patterns[30082] = 29'b0_111010110000_010_1_110101100000;
      patterns[30083] = 29'b0_111010110000_011_1_101011000001;
      patterns[30084] = 29'b0_111010110000_100_0_011101011000;
      patterns[30085] = 29'b0_111010110000_101_0_001110101100;
      patterns[30086] = 29'b0_111010110000_110_0_111010110000;
      patterns[30087] = 29'b0_111010110000_111_0_111010110000;
      patterns[30088] = 29'b0_111010110001_000_0_111010110001;
      patterns[30089] = 29'b0_111010110001_001_0_110001111010;
      patterns[30090] = 29'b0_111010110001_010_1_110101100010;
      patterns[30091] = 29'b0_111010110001_011_1_101011000101;
      patterns[30092] = 29'b0_111010110001_100_1_011101011000;
      patterns[30093] = 29'b0_111010110001_101_0_101110101100;
      patterns[30094] = 29'b0_111010110001_110_0_111010110001;
      patterns[30095] = 29'b0_111010110001_111_0_111010110001;
      patterns[30096] = 29'b0_111010110010_000_0_111010110010;
      patterns[30097] = 29'b0_111010110010_001_0_110010111010;
      patterns[30098] = 29'b0_111010110010_010_1_110101100100;
      patterns[30099] = 29'b0_111010110010_011_1_101011001001;
      patterns[30100] = 29'b0_111010110010_100_0_011101011001;
      patterns[30101] = 29'b0_111010110010_101_1_001110101100;
      patterns[30102] = 29'b0_111010110010_110_0_111010110010;
      patterns[30103] = 29'b0_111010110010_111_0_111010110010;
      patterns[30104] = 29'b0_111010110011_000_0_111010110011;
      patterns[30105] = 29'b0_111010110011_001_0_110011111010;
      patterns[30106] = 29'b0_111010110011_010_1_110101100110;
      patterns[30107] = 29'b0_111010110011_011_1_101011001101;
      patterns[30108] = 29'b0_111010110011_100_1_011101011001;
      patterns[30109] = 29'b0_111010110011_101_1_101110101100;
      patterns[30110] = 29'b0_111010110011_110_0_111010110011;
      patterns[30111] = 29'b0_111010110011_111_0_111010110011;
      patterns[30112] = 29'b0_111010110100_000_0_111010110100;
      patterns[30113] = 29'b0_111010110100_001_0_110100111010;
      patterns[30114] = 29'b0_111010110100_010_1_110101101000;
      patterns[30115] = 29'b0_111010110100_011_1_101011010001;
      patterns[30116] = 29'b0_111010110100_100_0_011101011010;
      patterns[30117] = 29'b0_111010110100_101_0_001110101101;
      patterns[30118] = 29'b0_111010110100_110_0_111010110100;
      patterns[30119] = 29'b0_111010110100_111_0_111010110100;
      patterns[30120] = 29'b0_111010110101_000_0_111010110101;
      patterns[30121] = 29'b0_111010110101_001_0_110101111010;
      patterns[30122] = 29'b0_111010110101_010_1_110101101010;
      patterns[30123] = 29'b0_111010110101_011_1_101011010101;
      patterns[30124] = 29'b0_111010110101_100_1_011101011010;
      patterns[30125] = 29'b0_111010110101_101_0_101110101101;
      patterns[30126] = 29'b0_111010110101_110_0_111010110101;
      patterns[30127] = 29'b0_111010110101_111_0_111010110101;
      patterns[30128] = 29'b0_111010110110_000_0_111010110110;
      patterns[30129] = 29'b0_111010110110_001_0_110110111010;
      patterns[30130] = 29'b0_111010110110_010_1_110101101100;
      patterns[30131] = 29'b0_111010110110_011_1_101011011001;
      patterns[30132] = 29'b0_111010110110_100_0_011101011011;
      patterns[30133] = 29'b0_111010110110_101_1_001110101101;
      patterns[30134] = 29'b0_111010110110_110_0_111010110110;
      patterns[30135] = 29'b0_111010110110_111_0_111010110110;
      patterns[30136] = 29'b0_111010110111_000_0_111010110111;
      patterns[30137] = 29'b0_111010110111_001_0_110111111010;
      patterns[30138] = 29'b0_111010110111_010_1_110101101110;
      patterns[30139] = 29'b0_111010110111_011_1_101011011101;
      patterns[30140] = 29'b0_111010110111_100_1_011101011011;
      patterns[30141] = 29'b0_111010110111_101_1_101110101101;
      patterns[30142] = 29'b0_111010110111_110_0_111010110111;
      patterns[30143] = 29'b0_111010110111_111_0_111010110111;
      patterns[30144] = 29'b0_111010111000_000_0_111010111000;
      patterns[30145] = 29'b0_111010111000_001_0_111000111010;
      patterns[30146] = 29'b0_111010111000_010_1_110101110000;
      patterns[30147] = 29'b0_111010111000_011_1_101011100001;
      patterns[30148] = 29'b0_111010111000_100_0_011101011100;
      patterns[30149] = 29'b0_111010111000_101_0_001110101110;
      patterns[30150] = 29'b0_111010111000_110_0_111010111000;
      patterns[30151] = 29'b0_111010111000_111_0_111010111000;
      patterns[30152] = 29'b0_111010111001_000_0_111010111001;
      patterns[30153] = 29'b0_111010111001_001_0_111001111010;
      patterns[30154] = 29'b0_111010111001_010_1_110101110010;
      patterns[30155] = 29'b0_111010111001_011_1_101011100101;
      patterns[30156] = 29'b0_111010111001_100_1_011101011100;
      patterns[30157] = 29'b0_111010111001_101_0_101110101110;
      patterns[30158] = 29'b0_111010111001_110_0_111010111001;
      patterns[30159] = 29'b0_111010111001_111_0_111010111001;
      patterns[30160] = 29'b0_111010111010_000_0_111010111010;
      patterns[30161] = 29'b0_111010111010_001_0_111010111010;
      patterns[30162] = 29'b0_111010111010_010_1_110101110100;
      patterns[30163] = 29'b0_111010111010_011_1_101011101001;
      patterns[30164] = 29'b0_111010111010_100_0_011101011101;
      patterns[30165] = 29'b0_111010111010_101_1_001110101110;
      patterns[30166] = 29'b0_111010111010_110_0_111010111010;
      patterns[30167] = 29'b0_111010111010_111_0_111010111010;
      patterns[30168] = 29'b0_111010111011_000_0_111010111011;
      patterns[30169] = 29'b0_111010111011_001_0_111011111010;
      patterns[30170] = 29'b0_111010111011_010_1_110101110110;
      patterns[30171] = 29'b0_111010111011_011_1_101011101101;
      patterns[30172] = 29'b0_111010111011_100_1_011101011101;
      patterns[30173] = 29'b0_111010111011_101_1_101110101110;
      patterns[30174] = 29'b0_111010111011_110_0_111010111011;
      patterns[30175] = 29'b0_111010111011_111_0_111010111011;
      patterns[30176] = 29'b0_111010111100_000_0_111010111100;
      patterns[30177] = 29'b0_111010111100_001_0_111100111010;
      patterns[30178] = 29'b0_111010111100_010_1_110101111000;
      patterns[30179] = 29'b0_111010111100_011_1_101011110001;
      patterns[30180] = 29'b0_111010111100_100_0_011101011110;
      patterns[30181] = 29'b0_111010111100_101_0_001110101111;
      patterns[30182] = 29'b0_111010111100_110_0_111010111100;
      patterns[30183] = 29'b0_111010111100_111_0_111010111100;
      patterns[30184] = 29'b0_111010111101_000_0_111010111101;
      patterns[30185] = 29'b0_111010111101_001_0_111101111010;
      patterns[30186] = 29'b0_111010111101_010_1_110101111010;
      patterns[30187] = 29'b0_111010111101_011_1_101011110101;
      patterns[30188] = 29'b0_111010111101_100_1_011101011110;
      patterns[30189] = 29'b0_111010111101_101_0_101110101111;
      patterns[30190] = 29'b0_111010111101_110_0_111010111101;
      patterns[30191] = 29'b0_111010111101_111_0_111010111101;
      patterns[30192] = 29'b0_111010111110_000_0_111010111110;
      patterns[30193] = 29'b0_111010111110_001_0_111110111010;
      patterns[30194] = 29'b0_111010111110_010_1_110101111100;
      patterns[30195] = 29'b0_111010111110_011_1_101011111001;
      patterns[30196] = 29'b0_111010111110_100_0_011101011111;
      patterns[30197] = 29'b0_111010111110_101_1_001110101111;
      patterns[30198] = 29'b0_111010111110_110_0_111010111110;
      patterns[30199] = 29'b0_111010111110_111_0_111010111110;
      patterns[30200] = 29'b0_111010111111_000_0_111010111111;
      patterns[30201] = 29'b0_111010111111_001_0_111111111010;
      patterns[30202] = 29'b0_111010111111_010_1_110101111110;
      patterns[30203] = 29'b0_111010111111_011_1_101011111101;
      patterns[30204] = 29'b0_111010111111_100_1_011101011111;
      patterns[30205] = 29'b0_111010111111_101_1_101110101111;
      patterns[30206] = 29'b0_111010111111_110_0_111010111111;
      patterns[30207] = 29'b0_111010111111_111_0_111010111111;
      patterns[30208] = 29'b0_111011000000_000_0_111011000000;
      patterns[30209] = 29'b0_111011000000_001_0_000000111011;
      patterns[30210] = 29'b0_111011000000_010_1_110110000000;
      patterns[30211] = 29'b0_111011000000_011_1_101100000001;
      patterns[30212] = 29'b0_111011000000_100_0_011101100000;
      patterns[30213] = 29'b0_111011000000_101_0_001110110000;
      patterns[30214] = 29'b0_111011000000_110_0_111011000000;
      patterns[30215] = 29'b0_111011000000_111_0_111011000000;
      patterns[30216] = 29'b0_111011000001_000_0_111011000001;
      patterns[30217] = 29'b0_111011000001_001_0_000001111011;
      patterns[30218] = 29'b0_111011000001_010_1_110110000010;
      patterns[30219] = 29'b0_111011000001_011_1_101100000101;
      patterns[30220] = 29'b0_111011000001_100_1_011101100000;
      patterns[30221] = 29'b0_111011000001_101_0_101110110000;
      patterns[30222] = 29'b0_111011000001_110_0_111011000001;
      patterns[30223] = 29'b0_111011000001_111_0_111011000001;
      patterns[30224] = 29'b0_111011000010_000_0_111011000010;
      patterns[30225] = 29'b0_111011000010_001_0_000010111011;
      patterns[30226] = 29'b0_111011000010_010_1_110110000100;
      patterns[30227] = 29'b0_111011000010_011_1_101100001001;
      patterns[30228] = 29'b0_111011000010_100_0_011101100001;
      patterns[30229] = 29'b0_111011000010_101_1_001110110000;
      patterns[30230] = 29'b0_111011000010_110_0_111011000010;
      patterns[30231] = 29'b0_111011000010_111_0_111011000010;
      patterns[30232] = 29'b0_111011000011_000_0_111011000011;
      patterns[30233] = 29'b0_111011000011_001_0_000011111011;
      patterns[30234] = 29'b0_111011000011_010_1_110110000110;
      patterns[30235] = 29'b0_111011000011_011_1_101100001101;
      patterns[30236] = 29'b0_111011000011_100_1_011101100001;
      patterns[30237] = 29'b0_111011000011_101_1_101110110000;
      patterns[30238] = 29'b0_111011000011_110_0_111011000011;
      patterns[30239] = 29'b0_111011000011_111_0_111011000011;
      patterns[30240] = 29'b0_111011000100_000_0_111011000100;
      patterns[30241] = 29'b0_111011000100_001_0_000100111011;
      patterns[30242] = 29'b0_111011000100_010_1_110110001000;
      patterns[30243] = 29'b0_111011000100_011_1_101100010001;
      patterns[30244] = 29'b0_111011000100_100_0_011101100010;
      patterns[30245] = 29'b0_111011000100_101_0_001110110001;
      patterns[30246] = 29'b0_111011000100_110_0_111011000100;
      patterns[30247] = 29'b0_111011000100_111_0_111011000100;
      patterns[30248] = 29'b0_111011000101_000_0_111011000101;
      patterns[30249] = 29'b0_111011000101_001_0_000101111011;
      patterns[30250] = 29'b0_111011000101_010_1_110110001010;
      patterns[30251] = 29'b0_111011000101_011_1_101100010101;
      patterns[30252] = 29'b0_111011000101_100_1_011101100010;
      patterns[30253] = 29'b0_111011000101_101_0_101110110001;
      patterns[30254] = 29'b0_111011000101_110_0_111011000101;
      patterns[30255] = 29'b0_111011000101_111_0_111011000101;
      patterns[30256] = 29'b0_111011000110_000_0_111011000110;
      patterns[30257] = 29'b0_111011000110_001_0_000110111011;
      patterns[30258] = 29'b0_111011000110_010_1_110110001100;
      patterns[30259] = 29'b0_111011000110_011_1_101100011001;
      patterns[30260] = 29'b0_111011000110_100_0_011101100011;
      patterns[30261] = 29'b0_111011000110_101_1_001110110001;
      patterns[30262] = 29'b0_111011000110_110_0_111011000110;
      patterns[30263] = 29'b0_111011000110_111_0_111011000110;
      patterns[30264] = 29'b0_111011000111_000_0_111011000111;
      patterns[30265] = 29'b0_111011000111_001_0_000111111011;
      patterns[30266] = 29'b0_111011000111_010_1_110110001110;
      patterns[30267] = 29'b0_111011000111_011_1_101100011101;
      patterns[30268] = 29'b0_111011000111_100_1_011101100011;
      patterns[30269] = 29'b0_111011000111_101_1_101110110001;
      patterns[30270] = 29'b0_111011000111_110_0_111011000111;
      patterns[30271] = 29'b0_111011000111_111_0_111011000111;
      patterns[30272] = 29'b0_111011001000_000_0_111011001000;
      patterns[30273] = 29'b0_111011001000_001_0_001000111011;
      patterns[30274] = 29'b0_111011001000_010_1_110110010000;
      patterns[30275] = 29'b0_111011001000_011_1_101100100001;
      patterns[30276] = 29'b0_111011001000_100_0_011101100100;
      patterns[30277] = 29'b0_111011001000_101_0_001110110010;
      patterns[30278] = 29'b0_111011001000_110_0_111011001000;
      patterns[30279] = 29'b0_111011001000_111_0_111011001000;
      patterns[30280] = 29'b0_111011001001_000_0_111011001001;
      patterns[30281] = 29'b0_111011001001_001_0_001001111011;
      patterns[30282] = 29'b0_111011001001_010_1_110110010010;
      patterns[30283] = 29'b0_111011001001_011_1_101100100101;
      patterns[30284] = 29'b0_111011001001_100_1_011101100100;
      patterns[30285] = 29'b0_111011001001_101_0_101110110010;
      patterns[30286] = 29'b0_111011001001_110_0_111011001001;
      patterns[30287] = 29'b0_111011001001_111_0_111011001001;
      patterns[30288] = 29'b0_111011001010_000_0_111011001010;
      patterns[30289] = 29'b0_111011001010_001_0_001010111011;
      patterns[30290] = 29'b0_111011001010_010_1_110110010100;
      patterns[30291] = 29'b0_111011001010_011_1_101100101001;
      patterns[30292] = 29'b0_111011001010_100_0_011101100101;
      patterns[30293] = 29'b0_111011001010_101_1_001110110010;
      patterns[30294] = 29'b0_111011001010_110_0_111011001010;
      patterns[30295] = 29'b0_111011001010_111_0_111011001010;
      patterns[30296] = 29'b0_111011001011_000_0_111011001011;
      patterns[30297] = 29'b0_111011001011_001_0_001011111011;
      patterns[30298] = 29'b0_111011001011_010_1_110110010110;
      patterns[30299] = 29'b0_111011001011_011_1_101100101101;
      patterns[30300] = 29'b0_111011001011_100_1_011101100101;
      patterns[30301] = 29'b0_111011001011_101_1_101110110010;
      patterns[30302] = 29'b0_111011001011_110_0_111011001011;
      patterns[30303] = 29'b0_111011001011_111_0_111011001011;
      patterns[30304] = 29'b0_111011001100_000_0_111011001100;
      patterns[30305] = 29'b0_111011001100_001_0_001100111011;
      patterns[30306] = 29'b0_111011001100_010_1_110110011000;
      patterns[30307] = 29'b0_111011001100_011_1_101100110001;
      patterns[30308] = 29'b0_111011001100_100_0_011101100110;
      patterns[30309] = 29'b0_111011001100_101_0_001110110011;
      patterns[30310] = 29'b0_111011001100_110_0_111011001100;
      patterns[30311] = 29'b0_111011001100_111_0_111011001100;
      patterns[30312] = 29'b0_111011001101_000_0_111011001101;
      patterns[30313] = 29'b0_111011001101_001_0_001101111011;
      patterns[30314] = 29'b0_111011001101_010_1_110110011010;
      patterns[30315] = 29'b0_111011001101_011_1_101100110101;
      patterns[30316] = 29'b0_111011001101_100_1_011101100110;
      patterns[30317] = 29'b0_111011001101_101_0_101110110011;
      patterns[30318] = 29'b0_111011001101_110_0_111011001101;
      patterns[30319] = 29'b0_111011001101_111_0_111011001101;
      patterns[30320] = 29'b0_111011001110_000_0_111011001110;
      patterns[30321] = 29'b0_111011001110_001_0_001110111011;
      patterns[30322] = 29'b0_111011001110_010_1_110110011100;
      patterns[30323] = 29'b0_111011001110_011_1_101100111001;
      patterns[30324] = 29'b0_111011001110_100_0_011101100111;
      patterns[30325] = 29'b0_111011001110_101_1_001110110011;
      patterns[30326] = 29'b0_111011001110_110_0_111011001110;
      patterns[30327] = 29'b0_111011001110_111_0_111011001110;
      patterns[30328] = 29'b0_111011001111_000_0_111011001111;
      patterns[30329] = 29'b0_111011001111_001_0_001111111011;
      patterns[30330] = 29'b0_111011001111_010_1_110110011110;
      patterns[30331] = 29'b0_111011001111_011_1_101100111101;
      patterns[30332] = 29'b0_111011001111_100_1_011101100111;
      patterns[30333] = 29'b0_111011001111_101_1_101110110011;
      patterns[30334] = 29'b0_111011001111_110_0_111011001111;
      patterns[30335] = 29'b0_111011001111_111_0_111011001111;
      patterns[30336] = 29'b0_111011010000_000_0_111011010000;
      patterns[30337] = 29'b0_111011010000_001_0_010000111011;
      patterns[30338] = 29'b0_111011010000_010_1_110110100000;
      patterns[30339] = 29'b0_111011010000_011_1_101101000001;
      patterns[30340] = 29'b0_111011010000_100_0_011101101000;
      patterns[30341] = 29'b0_111011010000_101_0_001110110100;
      patterns[30342] = 29'b0_111011010000_110_0_111011010000;
      patterns[30343] = 29'b0_111011010000_111_0_111011010000;
      patterns[30344] = 29'b0_111011010001_000_0_111011010001;
      patterns[30345] = 29'b0_111011010001_001_0_010001111011;
      patterns[30346] = 29'b0_111011010001_010_1_110110100010;
      patterns[30347] = 29'b0_111011010001_011_1_101101000101;
      patterns[30348] = 29'b0_111011010001_100_1_011101101000;
      patterns[30349] = 29'b0_111011010001_101_0_101110110100;
      patterns[30350] = 29'b0_111011010001_110_0_111011010001;
      patterns[30351] = 29'b0_111011010001_111_0_111011010001;
      patterns[30352] = 29'b0_111011010010_000_0_111011010010;
      patterns[30353] = 29'b0_111011010010_001_0_010010111011;
      patterns[30354] = 29'b0_111011010010_010_1_110110100100;
      patterns[30355] = 29'b0_111011010010_011_1_101101001001;
      patterns[30356] = 29'b0_111011010010_100_0_011101101001;
      patterns[30357] = 29'b0_111011010010_101_1_001110110100;
      patterns[30358] = 29'b0_111011010010_110_0_111011010010;
      patterns[30359] = 29'b0_111011010010_111_0_111011010010;
      patterns[30360] = 29'b0_111011010011_000_0_111011010011;
      patterns[30361] = 29'b0_111011010011_001_0_010011111011;
      patterns[30362] = 29'b0_111011010011_010_1_110110100110;
      patterns[30363] = 29'b0_111011010011_011_1_101101001101;
      patterns[30364] = 29'b0_111011010011_100_1_011101101001;
      patterns[30365] = 29'b0_111011010011_101_1_101110110100;
      patterns[30366] = 29'b0_111011010011_110_0_111011010011;
      patterns[30367] = 29'b0_111011010011_111_0_111011010011;
      patterns[30368] = 29'b0_111011010100_000_0_111011010100;
      patterns[30369] = 29'b0_111011010100_001_0_010100111011;
      patterns[30370] = 29'b0_111011010100_010_1_110110101000;
      patterns[30371] = 29'b0_111011010100_011_1_101101010001;
      patterns[30372] = 29'b0_111011010100_100_0_011101101010;
      patterns[30373] = 29'b0_111011010100_101_0_001110110101;
      patterns[30374] = 29'b0_111011010100_110_0_111011010100;
      patterns[30375] = 29'b0_111011010100_111_0_111011010100;
      patterns[30376] = 29'b0_111011010101_000_0_111011010101;
      patterns[30377] = 29'b0_111011010101_001_0_010101111011;
      patterns[30378] = 29'b0_111011010101_010_1_110110101010;
      patterns[30379] = 29'b0_111011010101_011_1_101101010101;
      patterns[30380] = 29'b0_111011010101_100_1_011101101010;
      patterns[30381] = 29'b0_111011010101_101_0_101110110101;
      patterns[30382] = 29'b0_111011010101_110_0_111011010101;
      patterns[30383] = 29'b0_111011010101_111_0_111011010101;
      patterns[30384] = 29'b0_111011010110_000_0_111011010110;
      patterns[30385] = 29'b0_111011010110_001_0_010110111011;
      patterns[30386] = 29'b0_111011010110_010_1_110110101100;
      patterns[30387] = 29'b0_111011010110_011_1_101101011001;
      patterns[30388] = 29'b0_111011010110_100_0_011101101011;
      patterns[30389] = 29'b0_111011010110_101_1_001110110101;
      patterns[30390] = 29'b0_111011010110_110_0_111011010110;
      patterns[30391] = 29'b0_111011010110_111_0_111011010110;
      patterns[30392] = 29'b0_111011010111_000_0_111011010111;
      patterns[30393] = 29'b0_111011010111_001_0_010111111011;
      patterns[30394] = 29'b0_111011010111_010_1_110110101110;
      patterns[30395] = 29'b0_111011010111_011_1_101101011101;
      patterns[30396] = 29'b0_111011010111_100_1_011101101011;
      patterns[30397] = 29'b0_111011010111_101_1_101110110101;
      patterns[30398] = 29'b0_111011010111_110_0_111011010111;
      patterns[30399] = 29'b0_111011010111_111_0_111011010111;
      patterns[30400] = 29'b0_111011011000_000_0_111011011000;
      patterns[30401] = 29'b0_111011011000_001_0_011000111011;
      patterns[30402] = 29'b0_111011011000_010_1_110110110000;
      patterns[30403] = 29'b0_111011011000_011_1_101101100001;
      patterns[30404] = 29'b0_111011011000_100_0_011101101100;
      patterns[30405] = 29'b0_111011011000_101_0_001110110110;
      patterns[30406] = 29'b0_111011011000_110_0_111011011000;
      patterns[30407] = 29'b0_111011011000_111_0_111011011000;
      patterns[30408] = 29'b0_111011011001_000_0_111011011001;
      patterns[30409] = 29'b0_111011011001_001_0_011001111011;
      patterns[30410] = 29'b0_111011011001_010_1_110110110010;
      patterns[30411] = 29'b0_111011011001_011_1_101101100101;
      patterns[30412] = 29'b0_111011011001_100_1_011101101100;
      patterns[30413] = 29'b0_111011011001_101_0_101110110110;
      patterns[30414] = 29'b0_111011011001_110_0_111011011001;
      patterns[30415] = 29'b0_111011011001_111_0_111011011001;
      patterns[30416] = 29'b0_111011011010_000_0_111011011010;
      patterns[30417] = 29'b0_111011011010_001_0_011010111011;
      patterns[30418] = 29'b0_111011011010_010_1_110110110100;
      patterns[30419] = 29'b0_111011011010_011_1_101101101001;
      patterns[30420] = 29'b0_111011011010_100_0_011101101101;
      patterns[30421] = 29'b0_111011011010_101_1_001110110110;
      patterns[30422] = 29'b0_111011011010_110_0_111011011010;
      patterns[30423] = 29'b0_111011011010_111_0_111011011010;
      patterns[30424] = 29'b0_111011011011_000_0_111011011011;
      patterns[30425] = 29'b0_111011011011_001_0_011011111011;
      patterns[30426] = 29'b0_111011011011_010_1_110110110110;
      patterns[30427] = 29'b0_111011011011_011_1_101101101101;
      patterns[30428] = 29'b0_111011011011_100_1_011101101101;
      patterns[30429] = 29'b0_111011011011_101_1_101110110110;
      patterns[30430] = 29'b0_111011011011_110_0_111011011011;
      patterns[30431] = 29'b0_111011011011_111_0_111011011011;
      patterns[30432] = 29'b0_111011011100_000_0_111011011100;
      patterns[30433] = 29'b0_111011011100_001_0_011100111011;
      patterns[30434] = 29'b0_111011011100_010_1_110110111000;
      patterns[30435] = 29'b0_111011011100_011_1_101101110001;
      patterns[30436] = 29'b0_111011011100_100_0_011101101110;
      patterns[30437] = 29'b0_111011011100_101_0_001110110111;
      patterns[30438] = 29'b0_111011011100_110_0_111011011100;
      patterns[30439] = 29'b0_111011011100_111_0_111011011100;
      patterns[30440] = 29'b0_111011011101_000_0_111011011101;
      patterns[30441] = 29'b0_111011011101_001_0_011101111011;
      patterns[30442] = 29'b0_111011011101_010_1_110110111010;
      patterns[30443] = 29'b0_111011011101_011_1_101101110101;
      patterns[30444] = 29'b0_111011011101_100_1_011101101110;
      patterns[30445] = 29'b0_111011011101_101_0_101110110111;
      patterns[30446] = 29'b0_111011011101_110_0_111011011101;
      patterns[30447] = 29'b0_111011011101_111_0_111011011101;
      patterns[30448] = 29'b0_111011011110_000_0_111011011110;
      patterns[30449] = 29'b0_111011011110_001_0_011110111011;
      patterns[30450] = 29'b0_111011011110_010_1_110110111100;
      patterns[30451] = 29'b0_111011011110_011_1_101101111001;
      patterns[30452] = 29'b0_111011011110_100_0_011101101111;
      patterns[30453] = 29'b0_111011011110_101_1_001110110111;
      patterns[30454] = 29'b0_111011011110_110_0_111011011110;
      patterns[30455] = 29'b0_111011011110_111_0_111011011110;
      patterns[30456] = 29'b0_111011011111_000_0_111011011111;
      patterns[30457] = 29'b0_111011011111_001_0_011111111011;
      patterns[30458] = 29'b0_111011011111_010_1_110110111110;
      patterns[30459] = 29'b0_111011011111_011_1_101101111101;
      patterns[30460] = 29'b0_111011011111_100_1_011101101111;
      patterns[30461] = 29'b0_111011011111_101_1_101110110111;
      patterns[30462] = 29'b0_111011011111_110_0_111011011111;
      patterns[30463] = 29'b0_111011011111_111_0_111011011111;
      patterns[30464] = 29'b0_111011100000_000_0_111011100000;
      patterns[30465] = 29'b0_111011100000_001_0_100000111011;
      patterns[30466] = 29'b0_111011100000_010_1_110111000000;
      patterns[30467] = 29'b0_111011100000_011_1_101110000001;
      patterns[30468] = 29'b0_111011100000_100_0_011101110000;
      patterns[30469] = 29'b0_111011100000_101_0_001110111000;
      patterns[30470] = 29'b0_111011100000_110_0_111011100000;
      patterns[30471] = 29'b0_111011100000_111_0_111011100000;
      patterns[30472] = 29'b0_111011100001_000_0_111011100001;
      patterns[30473] = 29'b0_111011100001_001_0_100001111011;
      patterns[30474] = 29'b0_111011100001_010_1_110111000010;
      patterns[30475] = 29'b0_111011100001_011_1_101110000101;
      patterns[30476] = 29'b0_111011100001_100_1_011101110000;
      patterns[30477] = 29'b0_111011100001_101_0_101110111000;
      patterns[30478] = 29'b0_111011100001_110_0_111011100001;
      patterns[30479] = 29'b0_111011100001_111_0_111011100001;
      patterns[30480] = 29'b0_111011100010_000_0_111011100010;
      patterns[30481] = 29'b0_111011100010_001_0_100010111011;
      patterns[30482] = 29'b0_111011100010_010_1_110111000100;
      patterns[30483] = 29'b0_111011100010_011_1_101110001001;
      patterns[30484] = 29'b0_111011100010_100_0_011101110001;
      patterns[30485] = 29'b0_111011100010_101_1_001110111000;
      patterns[30486] = 29'b0_111011100010_110_0_111011100010;
      patterns[30487] = 29'b0_111011100010_111_0_111011100010;
      patterns[30488] = 29'b0_111011100011_000_0_111011100011;
      patterns[30489] = 29'b0_111011100011_001_0_100011111011;
      patterns[30490] = 29'b0_111011100011_010_1_110111000110;
      patterns[30491] = 29'b0_111011100011_011_1_101110001101;
      patterns[30492] = 29'b0_111011100011_100_1_011101110001;
      patterns[30493] = 29'b0_111011100011_101_1_101110111000;
      patterns[30494] = 29'b0_111011100011_110_0_111011100011;
      patterns[30495] = 29'b0_111011100011_111_0_111011100011;
      patterns[30496] = 29'b0_111011100100_000_0_111011100100;
      patterns[30497] = 29'b0_111011100100_001_0_100100111011;
      patterns[30498] = 29'b0_111011100100_010_1_110111001000;
      patterns[30499] = 29'b0_111011100100_011_1_101110010001;
      patterns[30500] = 29'b0_111011100100_100_0_011101110010;
      patterns[30501] = 29'b0_111011100100_101_0_001110111001;
      patterns[30502] = 29'b0_111011100100_110_0_111011100100;
      patterns[30503] = 29'b0_111011100100_111_0_111011100100;
      patterns[30504] = 29'b0_111011100101_000_0_111011100101;
      patterns[30505] = 29'b0_111011100101_001_0_100101111011;
      patterns[30506] = 29'b0_111011100101_010_1_110111001010;
      patterns[30507] = 29'b0_111011100101_011_1_101110010101;
      patterns[30508] = 29'b0_111011100101_100_1_011101110010;
      patterns[30509] = 29'b0_111011100101_101_0_101110111001;
      patterns[30510] = 29'b0_111011100101_110_0_111011100101;
      patterns[30511] = 29'b0_111011100101_111_0_111011100101;
      patterns[30512] = 29'b0_111011100110_000_0_111011100110;
      patterns[30513] = 29'b0_111011100110_001_0_100110111011;
      patterns[30514] = 29'b0_111011100110_010_1_110111001100;
      patterns[30515] = 29'b0_111011100110_011_1_101110011001;
      patterns[30516] = 29'b0_111011100110_100_0_011101110011;
      patterns[30517] = 29'b0_111011100110_101_1_001110111001;
      patterns[30518] = 29'b0_111011100110_110_0_111011100110;
      patterns[30519] = 29'b0_111011100110_111_0_111011100110;
      patterns[30520] = 29'b0_111011100111_000_0_111011100111;
      patterns[30521] = 29'b0_111011100111_001_0_100111111011;
      patterns[30522] = 29'b0_111011100111_010_1_110111001110;
      patterns[30523] = 29'b0_111011100111_011_1_101110011101;
      patterns[30524] = 29'b0_111011100111_100_1_011101110011;
      patterns[30525] = 29'b0_111011100111_101_1_101110111001;
      patterns[30526] = 29'b0_111011100111_110_0_111011100111;
      patterns[30527] = 29'b0_111011100111_111_0_111011100111;
      patterns[30528] = 29'b0_111011101000_000_0_111011101000;
      patterns[30529] = 29'b0_111011101000_001_0_101000111011;
      patterns[30530] = 29'b0_111011101000_010_1_110111010000;
      patterns[30531] = 29'b0_111011101000_011_1_101110100001;
      patterns[30532] = 29'b0_111011101000_100_0_011101110100;
      patterns[30533] = 29'b0_111011101000_101_0_001110111010;
      patterns[30534] = 29'b0_111011101000_110_0_111011101000;
      patterns[30535] = 29'b0_111011101000_111_0_111011101000;
      patterns[30536] = 29'b0_111011101001_000_0_111011101001;
      patterns[30537] = 29'b0_111011101001_001_0_101001111011;
      patterns[30538] = 29'b0_111011101001_010_1_110111010010;
      patterns[30539] = 29'b0_111011101001_011_1_101110100101;
      patterns[30540] = 29'b0_111011101001_100_1_011101110100;
      patterns[30541] = 29'b0_111011101001_101_0_101110111010;
      patterns[30542] = 29'b0_111011101001_110_0_111011101001;
      patterns[30543] = 29'b0_111011101001_111_0_111011101001;
      patterns[30544] = 29'b0_111011101010_000_0_111011101010;
      patterns[30545] = 29'b0_111011101010_001_0_101010111011;
      patterns[30546] = 29'b0_111011101010_010_1_110111010100;
      patterns[30547] = 29'b0_111011101010_011_1_101110101001;
      patterns[30548] = 29'b0_111011101010_100_0_011101110101;
      patterns[30549] = 29'b0_111011101010_101_1_001110111010;
      patterns[30550] = 29'b0_111011101010_110_0_111011101010;
      patterns[30551] = 29'b0_111011101010_111_0_111011101010;
      patterns[30552] = 29'b0_111011101011_000_0_111011101011;
      patterns[30553] = 29'b0_111011101011_001_0_101011111011;
      patterns[30554] = 29'b0_111011101011_010_1_110111010110;
      patterns[30555] = 29'b0_111011101011_011_1_101110101101;
      patterns[30556] = 29'b0_111011101011_100_1_011101110101;
      patterns[30557] = 29'b0_111011101011_101_1_101110111010;
      patterns[30558] = 29'b0_111011101011_110_0_111011101011;
      patterns[30559] = 29'b0_111011101011_111_0_111011101011;
      patterns[30560] = 29'b0_111011101100_000_0_111011101100;
      patterns[30561] = 29'b0_111011101100_001_0_101100111011;
      patterns[30562] = 29'b0_111011101100_010_1_110111011000;
      patterns[30563] = 29'b0_111011101100_011_1_101110110001;
      patterns[30564] = 29'b0_111011101100_100_0_011101110110;
      patterns[30565] = 29'b0_111011101100_101_0_001110111011;
      patterns[30566] = 29'b0_111011101100_110_0_111011101100;
      patterns[30567] = 29'b0_111011101100_111_0_111011101100;
      patterns[30568] = 29'b0_111011101101_000_0_111011101101;
      patterns[30569] = 29'b0_111011101101_001_0_101101111011;
      patterns[30570] = 29'b0_111011101101_010_1_110111011010;
      patterns[30571] = 29'b0_111011101101_011_1_101110110101;
      patterns[30572] = 29'b0_111011101101_100_1_011101110110;
      patterns[30573] = 29'b0_111011101101_101_0_101110111011;
      patterns[30574] = 29'b0_111011101101_110_0_111011101101;
      patterns[30575] = 29'b0_111011101101_111_0_111011101101;
      patterns[30576] = 29'b0_111011101110_000_0_111011101110;
      patterns[30577] = 29'b0_111011101110_001_0_101110111011;
      patterns[30578] = 29'b0_111011101110_010_1_110111011100;
      patterns[30579] = 29'b0_111011101110_011_1_101110111001;
      patterns[30580] = 29'b0_111011101110_100_0_011101110111;
      patterns[30581] = 29'b0_111011101110_101_1_001110111011;
      patterns[30582] = 29'b0_111011101110_110_0_111011101110;
      patterns[30583] = 29'b0_111011101110_111_0_111011101110;
      patterns[30584] = 29'b0_111011101111_000_0_111011101111;
      patterns[30585] = 29'b0_111011101111_001_0_101111111011;
      patterns[30586] = 29'b0_111011101111_010_1_110111011110;
      patterns[30587] = 29'b0_111011101111_011_1_101110111101;
      patterns[30588] = 29'b0_111011101111_100_1_011101110111;
      patterns[30589] = 29'b0_111011101111_101_1_101110111011;
      patterns[30590] = 29'b0_111011101111_110_0_111011101111;
      patterns[30591] = 29'b0_111011101111_111_0_111011101111;
      patterns[30592] = 29'b0_111011110000_000_0_111011110000;
      patterns[30593] = 29'b0_111011110000_001_0_110000111011;
      patterns[30594] = 29'b0_111011110000_010_1_110111100000;
      patterns[30595] = 29'b0_111011110000_011_1_101111000001;
      patterns[30596] = 29'b0_111011110000_100_0_011101111000;
      patterns[30597] = 29'b0_111011110000_101_0_001110111100;
      patterns[30598] = 29'b0_111011110000_110_0_111011110000;
      patterns[30599] = 29'b0_111011110000_111_0_111011110000;
      patterns[30600] = 29'b0_111011110001_000_0_111011110001;
      patterns[30601] = 29'b0_111011110001_001_0_110001111011;
      patterns[30602] = 29'b0_111011110001_010_1_110111100010;
      patterns[30603] = 29'b0_111011110001_011_1_101111000101;
      patterns[30604] = 29'b0_111011110001_100_1_011101111000;
      patterns[30605] = 29'b0_111011110001_101_0_101110111100;
      patterns[30606] = 29'b0_111011110001_110_0_111011110001;
      patterns[30607] = 29'b0_111011110001_111_0_111011110001;
      patterns[30608] = 29'b0_111011110010_000_0_111011110010;
      patterns[30609] = 29'b0_111011110010_001_0_110010111011;
      patterns[30610] = 29'b0_111011110010_010_1_110111100100;
      patterns[30611] = 29'b0_111011110010_011_1_101111001001;
      patterns[30612] = 29'b0_111011110010_100_0_011101111001;
      patterns[30613] = 29'b0_111011110010_101_1_001110111100;
      patterns[30614] = 29'b0_111011110010_110_0_111011110010;
      patterns[30615] = 29'b0_111011110010_111_0_111011110010;
      patterns[30616] = 29'b0_111011110011_000_0_111011110011;
      patterns[30617] = 29'b0_111011110011_001_0_110011111011;
      patterns[30618] = 29'b0_111011110011_010_1_110111100110;
      patterns[30619] = 29'b0_111011110011_011_1_101111001101;
      patterns[30620] = 29'b0_111011110011_100_1_011101111001;
      patterns[30621] = 29'b0_111011110011_101_1_101110111100;
      patterns[30622] = 29'b0_111011110011_110_0_111011110011;
      patterns[30623] = 29'b0_111011110011_111_0_111011110011;
      patterns[30624] = 29'b0_111011110100_000_0_111011110100;
      patterns[30625] = 29'b0_111011110100_001_0_110100111011;
      patterns[30626] = 29'b0_111011110100_010_1_110111101000;
      patterns[30627] = 29'b0_111011110100_011_1_101111010001;
      patterns[30628] = 29'b0_111011110100_100_0_011101111010;
      patterns[30629] = 29'b0_111011110100_101_0_001110111101;
      patterns[30630] = 29'b0_111011110100_110_0_111011110100;
      patterns[30631] = 29'b0_111011110100_111_0_111011110100;
      patterns[30632] = 29'b0_111011110101_000_0_111011110101;
      patterns[30633] = 29'b0_111011110101_001_0_110101111011;
      patterns[30634] = 29'b0_111011110101_010_1_110111101010;
      patterns[30635] = 29'b0_111011110101_011_1_101111010101;
      patterns[30636] = 29'b0_111011110101_100_1_011101111010;
      patterns[30637] = 29'b0_111011110101_101_0_101110111101;
      patterns[30638] = 29'b0_111011110101_110_0_111011110101;
      patterns[30639] = 29'b0_111011110101_111_0_111011110101;
      patterns[30640] = 29'b0_111011110110_000_0_111011110110;
      patterns[30641] = 29'b0_111011110110_001_0_110110111011;
      patterns[30642] = 29'b0_111011110110_010_1_110111101100;
      patterns[30643] = 29'b0_111011110110_011_1_101111011001;
      patterns[30644] = 29'b0_111011110110_100_0_011101111011;
      patterns[30645] = 29'b0_111011110110_101_1_001110111101;
      patterns[30646] = 29'b0_111011110110_110_0_111011110110;
      patterns[30647] = 29'b0_111011110110_111_0_111011110110;
      patterns[30648] = 29'b0_111011110111_000_0_111011110111;
      patterns[30649] = 29'b0_111011110111_001_0_110111111011;
      patterns[30650] = 29'b0_111011110111_010_1_110111101110;
      patterns[30651] = 29'b0_111011110111_011_1_101111011101;
      patterns[30652] = 29'b0_111011110111_100_1_011101111011;
      patterns[30653] = 29'b0_111011110111_101_1_101110111101;
      patterns[30654] = 29'b0_111011110111_110_0_111011110111;
      patterns[30655] = 29'b0_111011110111_111_0_111011110111;
      patterns[30656] = 29'b0_111011111000_000_0_111011111000;
      patterns[30657] = 29'b0_111011111000_001_0_111000111011;
      patterns[30658] = 29'b0_111011111000_010_1_110111110000;
      patterns[30659] = 29'b0_111011111000_011_1_101111100001;
      patterns[30660] = 29'b0_111011111000_100_0_011101111100;
      patterns[30661] = 29'b0_111011111000_101_0_001110111110;
      patterns[30662] = 29'b0_111011111000_110_0_111011111000;
      patterns[30663] = 29'b0_111011111000_111_0_111011111000;
      patterns[30664] = 29'b0_111011111001_000_0_111011111001;
      patterns[30665] = 29'b0_111011111001_001_0_111001111011;
      patterns[30666] = 29'b0_111011111001_010_1_110111110010;
      patterns[30667] = 29'b0_111011111001_011_1_101111100101;
      patterns[30668] = 29'b0_111011111001_100_1_011101111100;
      patterns[30669] = 29'b0_111011111001_101_0_101110111110;
      patterns[30670] = 29'b0_111011111001_110_0_111011111001;
      patterns[30671] = 29'b0_111011111001_111_0_111011111001;
      patterns[30672] = 29'b0_111011111010_000_0_111011111010;
      patterns[30673] = 29'b0_111011111010_001_0_111010111011;
      patterns[30674] = 29'b0_111011111010_010_1_110111110100;
      patterns[30675] = 29'b0_111011111010_011_1_101111101001;
      patterns[30676] = 29'b0_111011111010_100_0_011101111101;
      patterns[30677] = 29'b0_111011111010_101_1_001110111110;
      patterns[30678] = 29'b0_111011111010_110_0_111011111010;
      patterns[30679] = 29'b0_111011111010_111_0_111011111010;
      patterns[30680] = 29'b0_111011111011_000_0_111011111011;
      patterns[30681] = 29'b0_111011111011_001_0_111011111011;
      patterns[30682] = 29'b0_111011111011_010_1_110111110110;
      patterns[30683] = 29'b0_111011111011_011_1_101111101101;
      patterns[30684] = 29'b0_111011111011_100_1_011101111101;
      patterns[30685] = 29'b0_111011111011_101_1_101110111110;
      patterns[30686] = 29'b0_111011111011_110_0_111011111011;
      patterns[30687] = 29'b0_111011111011_111_0_111011111011;
      patterns[30688] = 29'b0_111011111100_000_0_111011111100;
      patterns[30689] = 29'b0_111011111100_001_0_111100111011;
      patterns[30690] = 29'b0_111011111100_010_1_110111111000;
      patterns[30691] = 29'b0_111011111100_011_1_101111110001;
      patterns[30692] = 29'b0_111011111100_100_0_011101111110;
      patterns[30693] = 29'b0_111011111100_101_0_001110111111;
      patterns[30694] = 29'b0_111011111100_110_0_111011111100;
      patterns[30695] = 29'b0_111011111100_111_0_111011111100;
      patterns[30696] = 29'b0_111011111101_000_0_111011111101;
      patterns[30697] = 29'b0_111011111101_001_0_111101111011;
      patterns[30698] = 29'b0_111011111101_010_1_110111111010;
      patterns[30699] = 29'b0_111011111101_011_1_101111110101;
      patterns[30700] = 29'b0_111011111101_100_1_011101111110;
      patterns[30701] = 29'b0_111011111101_101_0_101110111111;
      patterns[30702] = 29'b0_111011111101_110_0_111011111101;
      patterns[30703] = 29'b0_111011111101_111_0_111011111101;
      patterns[30704] = 29'b0_111011111110_000_0_111011111110;
      patterns[30705] = 29'b0_111011111110_001_0_111110111011;
      patterns[30706] = 29'b0_111011111110_010_1_110111111100;
      patterns[30707] = 29'b0_111011111110_011_1_101111111001;
      patterns[30708] = 29'b0_111011111110_100_0_011101111111;
      patterns[30709] = 29'b0_111011111110_101_1_001110111111;
      patterns[30710] = 29'b0_111011111110_110_0_111011111110;
      patterns[30711] = 29'b0_111011111110_111_0_111011111110;
      patterns[30712] = 29'b0_111011111111_000_0_111011111111;
      patterns[30713] = 29'b0_111011111111_001_0_111111111011;
      patterns[30714] = 29'b0_111011111111_010_1_110111111110;
      patterns[30715] = 29'b0_111011111111_011_1_101111111101;
      patterns[30716] = 29'b0_111011111111_100_1_011101111111;
      patterns[30717] = 29'b0_111011111111_101_1_101110111111;
      patterns[30718] = 29'b0_111011111111_110_0_111011111111;
      patterns[30719] = 29'b0_111011111111_111_0_111011111111;
      patterns[30720] = 29'b0_111100000000_000_0_111100000000;
      patterns[30721] = 29'b0_111100000000_001_0_000000111100;
      patterns[30722] = 29'b0_111100000000_010_1_111000000000;
      patterns[30723] = 29'b0_111100000000_011_1_110000000001;
      patterns[30724] = 29'b0_111100000000_100_0_011110000000;
      patterns[30725] = 29'b0_111100000000_101_0_001111000000;
      patterns[30726] = 29'b0_111100000000_110_0_111100000000;
      patterns[30727] = 29'b0_111100000000_111_0_111100000000;
      patterns[30728] = 29'b0_111100000001_000_0_111100000001;
      patterns[30729] = 29'b0_111100000001_001_0_000001111100;
      patterns[30730] = 29'b0_111100000001_010_1_111000000010;
      patterns[30731] = 29'b0_111100000001_011_1_110000000101;
      patterns[30732] = 29'b0_111100000001_100_1_011110000000;
      patterns[30733] = 29'b0_111100000001_101_0_101111000000;
      patterns[30734] = 29'b0_111100000001_110_0_111100000001;
      patterns[30735] = 29'b0_111100000001_111_0_111100000001;
      patterns[30736] = 29'b0_111100000010_000_0_111100000010;
      patterns[30737] = 29'b0_111100000010_001_0_000010111100;
      patterns[30738] = 29'b0_111100000010_010_1_111000000100;
      patterns[30739] = 29'b0_111100000010_011_1_110000001001;
      patterns[30740] = 29'b0_111100000010_100_0_011110000001;
      patterns[30741] = 29'b0_111100000010_101_1_001111000000;
      patterns[30742] = 29'b0_111100000010_110_0_111100000010;
      patterns[30743] = 29'b0_111100000010_111_0_111100000010;
      patterns[30744] = 29'b0_111100000011_000_0_111100000011;
      patterns[30745] = 29'b0_111100000011_001_0_000011111100;
      patterns[30746] = 29'b0_111100000011_010_1_111000000110;
      patterns[30747] = 29'b0_111100000011_011_1_110000001101;
      patterns[30748] = 29'b0_111100000011_100_1_011110000001;
      patterns[30749] = 29'b0_111100000011_101_1_101111000000;
      patterns[30750] = 29'b0_111100000011_110_0_111100000011;
      patterns[30751] = 29'b0_111100000011_111_0_111100000011;
      patterns[30752] = 29'b0_111100000100_000_0_111100000100;
      patterns[30753] = 29'b0_111100000100_001_0_000100111100;
      patterns[30754] = 29'b0_111100000100_010_1_111000001000;
      patterns[30755] = 29'b0_111100000100_011_1_110000010001;
      patterns[30756] = 29'b0_111100000100_100_0_011110000010;
      patterns[30757] = 29'b0_111100000100_101_0_001111000001;
      patterns[30758] = 29'b0_111100000100_110_0_111100000100;
      patterns[30759] = 29'b0_111100000100_111_0_111100000100;
      patterns[30760] = 29'b0_111100000101_000_0_111100000101;
      patterns[30761] = 29'b0_111100000101_001_0_000101111100;
      patterns[30762] = 29'b0_111100000101_010_1_111000001010;
      patterns[30763] = 29'b0_111100000101_011_1_110000010101;
      patterns[30764] = 29'b0_111100000101_100_1_011110000010;
      patterns[30765] = 29'b0_111100000101_101_0_101111000001;
      patterns[30766] = 29'b0_111100000101_110_0_111100000101;
      patterns[30767] = 29'b0_111100000101_111_0_111100000101;
      patterns[30768] = 29'b0_111100000110_000_0_111100000110;
      patterns[30769] = 29'b0_111100000110_001_0_000110111100;
      patterns[30770] = 29'b0_111100000110_010_1_111000001100;
      patterns[30771] = 29'b0_111100000110_011_1_110000011001;
      patterns[30772] = 29'b0_111100000110_100_0_011110000011;
      patterns[30773] = 29'b0_111100000110_101_1_001111000001;
      patterns[30774] = 29'b0_111100000110_110_0_111100000110;
      patterns[30775] = 29'b0_111100000110_111_0_111100000110;
      patterns[30776] = 29'b0_111100000111_000_0_111100000111;
      patterns[30777] = 29'b0_111100000111_001_0_000111111100;
      patterns[30778] = 29'b0_111100000111_010_1_111000001110;
      patterns[30779] = 29'b0_111100000111_011_1_110000011101;
      patterns[30780] = 29'b0_111100000111_100_1_011110000011;
      patterns[30781] = 29'b0_111100000111_101_1_101111000001;
      patterns[30782] = 29'b0_111100000111_110_0_111100000111;
      patterns[30783] = 29'b0_111100000111_111_0_111100000111;
      patterns[30784] = 29'b0_111100001000_000_0_111100001000;
      patterns[30785] = 29'b0_111100001000_001_0_001000111100;
      patterns[30786] = 29'b0_111100001000_010_1_111000010000;
      patterns[30787] = 29'b0_111100001000_011_1_110000100001;
      patterns[30788] = 29'b0_111100001000_100_0_011110000100;
      patterns[30789] = 29'b0_111100001000_101_0_001111000010;
      patterns[30790] = 29'b0_111100001000_110_0_111100001000;
      patterns[30791] = 29'b0_111100001000_111_0_111100001000;
      patterns[30792] = 29'b0_111100001001_000_0_111100001001;
      patterns[30793] = 29'b0_111100001001_001_0_001001111100;
      patterns[30794] = 29'b0_111100001001_010_1_111000010010;
      patterns[30795] = 29'b0_111100001001_011_1_110000100101;
      patterns[30796] = 29'b0_111100001001_100_1_011110000100;
      patterns[30797] = 29'b0_111100001001_101_0_101111000010;
      patterns[30798] = 29'b0_111100001001_110_0_111100001001;
      patterns[30799] = 29'b0_111100001001_111_0_111100001001;
      patterns[30800] = 29'b0_111100001010_000_0_111100001010;
      patterns[30801] = 29'b0_111100001010_001_0_001010111100;
      patterns[30802] = 29'b0_111100001010_010_1_111000010100;
      patterns[30803] = 29'b0_111100001010_011_1_110000101001;
      patterns[30804] = 29'b0_111100001010_100_0_011110000101;
      patterns[30805] = 29'b0_111100001010_101_1_001111000010;
      patterns[30806] = 29'b0_111100001010_110_0_111100001010;
      patterns[30807] = 29'b0_111100001010_111_0_111100001010;
      patterns[30808] = 29'b0_111100001011_000_0_111100001011;
      patterns[30809] = 29'b0_111100001011_001_0_001011111100;
      patterns[30810] = 29'b0_111100001011_010_1_111000010110;
      patterns[30811] = 29'b0_111100001011_011_1_110000101101;
      patterns[30812] = 29'b0_111100001011_100_1_011110000101;
      patterns[30813] = 29'b0_111100001011_101_1_101111000010;
      patterns[30814] = 29'b0_111100001011_110_0_111100001011;
      patterns[30815] = 29'b0_111100001011_111_0_111100001011;
      patterns[30816] = 29'b0_111100001100_000_0_111100001100;
      patterns[30817] = 29'b0_111100001100_001_0_001100111100;
      patterns[30818] = 29'b0_111100001100_010_1_111000011000;
      patterns[30819] = 29'b0_111100001100_011_1_110000110001;
      patterns[30820] = 29'b0_111100001100_100_0_011110000110;
      patterns[30821] = 29'b0_111100001100_101_0_001111000011;
      patterns[30822] = 29'b0_111100001100_110_0_111100001100;
      patterns[30823] = 29'b0_111100001100_111_0_111100001100;
      patterns[30824] = 29'b0_111100001101_000_0_111100001101;
      patterns[30825] = 29'b0_111100001101_001_0_001101111100;
      patterns[30826] = 29'b0_111100001101_010_1_111000011010;
      patterns[30827] = 29'b0_111100001101_011_1_110000110101;
      patterns[30828] = 29'b0_111100001101_100_1_011110000110;
      patterns[30829] = 29'b0_111100001101_101_0_101111000011;
      patterns[30830] = 29'b0_111100001101_110_0_111100001101;
      patterns[30831] = 29'b0_111100001101_111_0_111100001101;
      patterns[30832] = 29'b0_111100001110_000_0_111100001110;
      patterns[30833] = 29'b0_111100001110_001_0_001110111100;
      patterns[30834] = 29'b0_111100001110_010_1_111000011100;
      patterns[30835] = 29'b0_111100001110_011_1_110000111001;
      patterns[30836] = 29'b0_111100001110_100_0_011110000111;
      patterns[30837] = 29'b0_111100001110_101_1_001111000011;
      patterns[30838] = 29'b0_111100001110_110_0_111100001110;
      patterns[30839] = 29'b0_111100001110_111_0_111100001110;
      patterns[30840] = 29'b0_111100001111_000_0_111100001111;
      patterns[30841] = 29'b0_111100001111_001_0_001111111100;
      patterns[30842] = 29'b0_111100001111_010_1_111000011110;
      patterns[30843] = 29'b0_111100001111_011_1_110000111101;
      patterns[30844] = 29'b0_111100001111_100_1_011110000111;
      patterns[30845] = 29'b0_111100001111_101_1_101111000011;
      patterns[30846] = 29'b0_111100001111_110_0_111100001111;
      patterns[30847] = 29'b0_111100001111_111_0_111100001111;
      patterns[30848] = 29'b0_111100010000_000_0_111100010000;
      patterns[30849] = 29'b0_111100010000_001_0_010000111100;
      patterns[30850] = 29'b0_111100010000_010_1_111000100000;
      patterns[30851] = 29'b0_111100010000_011_1_110001000001;
      patterns[30852] = 29'b0_111100010000_100_0_011110001000;
      patterns[30853] = 29'b0_111100010000_101_0_001111000100;
      patterns[30854] = 29'b0_111100010000_110_0_111100010000;
      patterns[30855] = 29'b0_111100010000_111_0_111100010000;
      patterns[30856] = 29'b0_111100010001_000_0_111100010001;
      patterns[30857] = 29'b0_111100010001_001_0_010001111100;
      patterns[30858] = 29'b0_111100010001_010_1_111000100010;
      patterns[30859] = 29'b0_111100010001_011_1_110001000101;
      patterns[30860] = 29'b0_111100010001_100_1_011110001000;
      patterns[30861] = 29'b0_111100010001_101_0_101111000100;
      patterns[30862] = 29'b0_111100010001_110_0_111100010001;
      patterns[30863] = 29'b0_111100010001_111_0_111100010001;
      patterns[30864] = 29'b0_111100010010_000_0_111100010010;
      patterns[30865] = 29'b0_111100010010_001_0_010010111100;
      patterns[30866] = 29'b0_111100010010_010_1_111000100100;
      patterns[30867] = 29'b0_111100010010_011_1_110001001001;
      patterns[30868] = 29'b0_111100010010_100_0_011110001001;
      patterns[30869] = 29'b0_111100010010_101_1_001111000100;
      patterns[30870] = 29'b0_111100010010_110_0_111100010010;
      patterns[30871] = 29'b0_111100010010_111_0_111100010010;
      patterns[30872] = 29'b0_111100010011_000_0_111100010011;
      patterns[30873] = 29'b0_111100010011_001_0_010011111100;
      patterns[30874] = 29'b0_111100010011_010_1_111000100110;
      patterns[30875] = 29'b0_111100010011_011_1_110001001101;
      patterns[30876] = 29'b0_111100010011_100_1_011110001001;
      patterns[30877] = 29'b0_111100010011_101_1_101111000100;
      patterns[30878] = 29'b0_111100010011_110_0_111100010011;
      patterns[30879] = 29'b0_111100010011_111_0_111100010011;
      patterns[30880] = 29'b0_111100010100_000_0_111100010100;
      patterns[30881] = 29'b0_111100010100_001_0_010100111100;
      patterns[30882] = 29'b0_111100010100_010_1_111000101000;
      patterns[30883] = 29'b0_111100010100_011_1_110001010001;
      patterns[30884] = 29'b0_111100010100_100_0_011110001010;
      patterns[30885] = 29'b0_111100010100_101_0_001111000101;
      patterns[30886] = 29'b0_111100010100_110_0_111100010100;
      patterns[30887] = 29'b0_111100010100_111_0_111100010100;
      patterns[30888] = 29'b0_111100010101_000_0_111100010101;
      patterns[30889] = 29'b0_111100010101_001_0_010101111100;
      patterns[30890] = 29'b0_111100010101_010_1_111000101010;
      patterns[30891] = 29'b0_111100010101_011_1_110001010101;
      patterns[30892] = 29'b0_111100010101_100_1_011110001010;
      patterns[30893] = 29'b0_111100010101_101_0_101111000101;
      patterns[30894] = 29'b0_111100010101_110_0_111100010101;
      patterns[30895] = 29'b0_111100010101_111_0_111100010101;
      patterns[30896] = 29'b0_111100010110_000_0_111100010110;
      patterns[30897] = 29'b0_111100010110_001_0_010110111100;
      patterns[30898] = 29'b0_111100010110_010_1_111000101100;
      patterns[30899] = 29'b0_111100010110_011_1_110001011001;
      patterns[30900] = 29'b0_111100010110_100_0_011110001011;
      patterns[30901] = 29'b0_111100010110_101_1_001111000101;
      patterns[30902] = 29'b0_111100010110_110_0_111100010110;
      patterns[30903] = 29'b0_111100010110_111_0_111100010110;
      patterns[30904] = 29'b0_111100010111_000_0_111100010111;
      patterns[30905] = 29'b0_111100010111_001_0_010111111100;
      patterns[30906] = 29'b0_111100010111_010_1_111000101110;
      patterns[30907] = 29'b0_111100010111_011_1_110001011101;
      patterns[30908] = 29'b0_111100010111_100_1_011110001011;
      patterns[30909] = 29'b0_111100010111_101_1_101111000101;
      patterns[30910] = 29'b0_111100010111_110_0_111100010111;
      patterns[30911] = 29'b0_111100010111_111_0_111100010111;
      patterns[30912] = 29'b0_111100011000_000_0_111100011000;
      patterns[30913] = 29'b0_111100011000_001_0_011000111100;
      patterns[30914] = 29'b0_111100011000_010_1_111000110000;
      patterns[30915] = 29'b0_111100011000_011_1_110001100001;
      patterns[30916] = 29'b0_111100011000_100_0_011110001100;
      patterns[30917] = 29'b0_111100011000_101_0_001111000110;
      patterns[30918] = 29'b0_111100011000_110_0_111100011000;
      patterns[30919] = 29'b0_111100011000_111_0_111100011000;
      patterns[30920] = 29'b0_111100011001_000_0_111100011001;
      patterns[30921] = 29'b0_111100011001_001_0_011001111100;
      patterns[30922] = 29'b0_111100011001_010_1_111000110010;
      patterns[30923] = 29'b0_111100011001_011_1_110001100101;
      patterns[30924] = 29'b0_111100011001_100_1_011110001100;
      patterns[30925] = 29'b0_111100011001_101_0_101111000110;
      patterns[30926] = 29'b0_111100011001_110_0_111100011001;
      patterns[30927] = 29'b0_111100011001_111_0_111100011001;
      patterns[30928] = 29'b0_111100011010_000_0_111100011010;
      patterns[30929] = 29'b0_111100011010_001_0_011010111100;
      patterns[30930] = 29'b0_111100011010_010_1_111000110100;
      patterns[30931] = 29'b0_111100011010_011_1_110001101001;
      patterns[30932] = 29'b0_111100011010_100_0_011110001101;
      patterns[30933] = 29'b0_111100011010_101_1_001111000110;
      patterns[30934] = 29'b0_111100011010_110_0_111100011010;
      patterns[30935] = 29'b0_111100011010_111_0_111100011010;
      patterns[30936] = 29'b0_111100011011_000_0_111100011011;
      patterns[30937] = 29'b0_111100011011_001_0_011011111100;
      patterns[30938] = 29'b0_111100011011_010_1_111000110110;
      patterns[30939] = 29'b0_111100011011_011_1_110001101101;
      patterns[30940] = 29'b0_111100011011_100_1_011110001101;
      patterns[30941] = 29'b0_111100011011_101_1_101111000110;
      patterns[30942] = 29'b0_111100011011_110_0_111100011011;
      patterns[30943] = 29'b0_111100011011_111_0_111100011011;
      patterns[30944] = 29'b0_111100011100_000_0_111100011100;
      patterns[30945] = 29'b0_111100011100_001_0_011100111100;
      patterns[30946] = 29'b0_111100011100_010_1_111000111000;
      patterns[30947] = 29'b0_111100011100_011_1_110001110001;
      patterns[30948] = 29'b0_111100011100_100_0_011110001110;
      patterns[30949] = 29'b0_111100011100_101_0_001111000111;
      patterns[30950] = 29'b0_111100011100_110_0_111100011100;
      patterns[30951] = 29'b0_111100011100_111_0_111100011100;
      patterns[30952] = 29'b0_111100011101_000_0_111100011101;
      patterns[30953] = 29'b0_111100011101_001_0_011101111100;
      patterns[30954] = 29'b0_111100011101_010_1_111000111010;
      patterns[30955] = 29'b0_111100011101_011_1_110001110101;
      patterns[30956] = 29'b0_111100011101_100_1_011110001110;
      patterns[30957] = 29'b0_111100011101_101_0_101111000111;
      patterns[30958] = 29'b0_111100011101_110_0_111100011101;
      patterns[30959] = 29'b0_111100011101_111_0_111100011101;
      patterns[30960] = 29'b0_111100011110_000_0_111100011110;
      patterns[30961] = 29'b0_111100011110_001_0_011110111100;
      patterns[30962] = 29'b0_111100011110_010_1_111000111100;
      patterns[30963] = 29'b0_111100011110_011_1_110001111001;
      patterns[30964] = 29'b0_111100011110_100_0_011110001111;
      patterns[30965] = 29'b0_111100011110_101_1_001111000111;
      patterns[30966] = 29'b0_111100011110_110_0_111100011110;
      patterns[30967] = 29'b0_111100011110_111_0_111100011110;
      patterns[30968] = 29'b0_111100011111_000_0_111100011111;
      patterns[30969] = 29'b0_111100011111_001_0_011111111100;
      patterns[30970] = 29'b0_111100011111_010_1_111000111110;
      patterns[30971] = 29'b0_111100011111_011_1_110001111101;
      patterns[30972] = 29'b0_111100011111_100_1_011110001111;
      patterns[30973] = 29'b0_111100011111_101_1_101111000111;
      patterns[30974] = 29'b0_111100011111_110_0_111100011111;
      patterns[30975] = 29'b0_111100011111_111_0_111100011111;
      patterns[30976] = 29'b0_111100100000_000_0_111100100000;
      patterns[30977] = 29'b0_111100100000_001_0_100000111100;
      patterns[30978] = 29'b0_111100100000_010_1_111001000000;
      patterns[30979] = 29'b0_111100100000_011_1_110010000001;
      patterns[30980] = 29'b0_111100100000_100_0_011110010000;
      patterns[30981] = 29'b0_111100100000_101_0_001111001000;
      patterns[30982] = 29'b0_111100100000_110_0_111100100000;
      patterns[30983] = 29'b0_111100100000_111_0_111100100000;
      patterns[30984] = 29'b0_111100100001_000_0_111100100001;
      patterns[30985] = 29'b0_111100100001_001_0_100001111100;
      patterns[30986] = 29'b0_111100100001_010_1_111001000010;
      patterns[30987] = 29'b0_111100100001_011_1_110010000101;
      patterns[30988] = 29'b0_111100100001_100_1_011110010000;
      patterns[30989] = 29'b0_111100100001_101_0_101111001000;
      patterns[30990] = 29'b0_111100100001_110_0_111100100001;
      patterns[30991] = 29'b0_111100100001_111_0_111100100001;
      patterns[30992] = 29'b0_111100100010_000_0_111100100010;
      patterns[30993] = 29'b0_111100100010_001_0_100010111100;
      patterns[30994] = 29'b0_111100100010_010_1_111001000100;
      patterns[30995] = 29'b0_111100100010_011_1_110010001001;
      patterns[30996] = 29'b0_111100100010_100_0_011110010001;
      patterns[30997] = 29'b0_111100100010_101_1_001111001000;
      patterns[30998] = 29'b0_111100100010_110_0_111100100010;
      patterns[30999] = 29'b0_111100100010_111_0_111100100010;
      patterns[31000] = 29'b0_111100100011_000_0_111100100011;
      patterns[31001] = 29'b0_111100100011_001_0_100011111100;
      patterns[31002] = 29'b0_111100100011_010_1_111001000110;
      patterns[31003] = 29'b0_111100100011_011_1_110010001101;
      patterns[31004] = 29'b0_111100100011_100_1_011110010001;
      patterns[31005] = 29'b0_111100100011_101_1_101111001000;
      patterns[31006] = 29'b0_111100100011_110_0_111100100011;
      patterns[31007] = 29'b0_111100100011_111_0_111100100011;
      patterns[31008] = 29'b0_111100100100_000_0_111100100100;
      patterns[31009] = 29'b0_111100100100_001_0_100100111100;
      patterns[31010] = 29'b0_111100100100_010_1_111001001000;
      patterns[31011] = 29'b0_111100100100_011_1_110010010001;
      patterns[31012] = 29'b0_111100100100_100_0_011110010010;
      patterns[31013] = 29'b0_111100100100_101_0_001111001001;
      patterns[31014] = 29'b0_111100100100_110_0_111100100100;
      patterns[31015] = 29'b0_111100100100_111_0_111100100100;
      patterns[31016] = 29'b0_111100100101_000_0_111100100101;
      patterns[31017] = 29'b0_111100100101_001_0_100101111100;
      patterns[31018] = 29'b0_111100100101_010_1_111001001010;
      patterns[31019] = 29'b0_111100100101_011_1_110010010101;
      patterns[31020] = 29'b0_111100100101_100_1_011110010010;
      patterns[31021] = 29'b0_111100100101_101_0_101111001001;
      patterns[31022] = 29'b0_111100100101_110_0_111100100101;
      patterns[31023] = 29'b0_111100100101_111_0_111100100101;
      patterns[31024] = 29'b0_111100100110_000_0_111100100110;
      patterns[31025] = 29'b0_111100100110_001_0_100110111100;
      patterns[31026] = 29'b0_111100100110_010_1_111001001100;
      patterns[31027] = 29'b0_111100100110_011_1_110010011001;
      patterns[31028] = 29'b0_111100100110_100_0_011110010011;
      patterns[31029] = 29'b0_111100100110_101_1_001111001001;
      patterns[31030] = 29'b0_111100100110_110_0_111100100110;
      patterns[31031] = 29'b0_111100100110_111_0_111100100110;
      patterns[31032] = 29'b0_111100100111_000_0_111100100111;
      patterns[31033] = 29'b0_111100100111_001_0_100111111100;
      patterns[31034] = 29'b0_111100100111_010_1_111001001110;
      patterns[31035] = 29'b0_111100100111_011_1_110010011101;
      patterns[31036] = 29'b0_111100100111_100_1_011110010011;
      patterns[31037] = 29'b0_111100100111_101_1_101111001001;
      patterns[31038] = 29'b0_111100100111_110_0_111100100111;
      patterns[31039] = 29'b0_111100100111_111_0_111100100111;
      patterns[31040] = 29'b0_111100101000_000_0_111100101000;
      patterns[31041] = 29'b0_111100101000_001_0_101000111100;
      patterns[31042] = 29'b0_111100101000_010_1_111001010000;
      patterns[31043] = 29'b0_111100101000_011_1_110010100001;
      patterns[31044] = 29'b0_111100101000_100_0_011110010100;
      patterns[31045] = 29'b0_111100101000_101_0_001111001010;
      patterns[31046] = 29'b0_111100101000_110_0_111100101000;
      patterns[31047] = 29'b0_111100101000_111_0_111100101000;
      patterns[31048] = 29'b0_111100101001_000_0_111100101001;
      patterns[31049] = 29'b0_111100101001_001_0_101001111100;
      patterns[31050] = 29'b0_111100101001_010_1_111001010010;
      patterns[31051] = 29'b0_111100101001_011_1_110010100101;
      patterns[31052] = 29'b0_111100101001_100_1_011110010100;
      patterns[31053] = 29'b0_111100101001_101_0_101111001010;
      patterns[31054] = 29'b0_111100101001_110_0_111100101001;
      patterns[31055] = 29'b0_111100101001_111_0_111100101001;
      patterns[31056] = 29'b0_111100101010_000_0_111100101010;
      patterns[31057] = 29'b0_111100101010_001_0_101010111100;
      patterns[31058] = 29'b0_111100101010_010_1_111001010100;
      patterns[31059] = 29'b0_111100101010_011_1_110010101001;
      patterns[31060] = 29'b0_111100101010_100_0_011110010101;
      patterns[31061] = 29'b0_111100101010_101_1_001111001010;
      patterns[31062] = 29'b0_111100101010_110_0_111100101010;
      patterns[31063] = 29'b0_111100101010_111_0_111100101010;
      patterns[31064] = 29'b0_111100101011_000_0_111100101011;
      patterns[31065] = 29'b0_111100101011_001_0_101011111100;
      patterns[31066] = 29'b0_111100101011_010_1_111001010110;
      patterns[31067] = 29'b0_111100101011_011_1_110010101101;
      patterns[31068] = 29'b0_111100101011_100_1_011110010101;
      patterns[31069] = 29'b0_111100101011_101_1_101111001010;
      patterns[31070] = 29'b0_111100101011_110_0_111100101011;
      patterns[31071] = 29'b0_111100101011_111_0_111100101011;
      patterns[31072] = 29'b0_111100101100_000_0_111100101100;
      patterns[31073] = 29'b0_111100101100_001_0_101100111100;
      patterns[31074] = 29'b0_111100101100_010_1_111001011000;
      patterns[31075] = 29'b0_111100101100_011_1_110010110001;
      patterns[31076] = 29'b0_111100101100_100_0_011110010110;
      patterns[31077] = 29'b0_111100101100_101_0_001111001011;
      patterns[31078] = 29'b0_111100101100_110_0_111100101100;
      patterns[31079] = 29'b0_111100101100_111_0_111100101100;
      patterns[31080] = 29'b0_111100101101_000_0_111100101101;
      patterns[31081] = 29'b0_111100101101_001_0_101101111100;
      patterns[31082] = 29'b0_111100101101_010_1_111001011010;
      patterns[31083] = 29'b0_111100101101_011_1_110010110101;
      patterns[31084] = 29'b0_111100101101_100_1_011110010110;
      patterns[31085] = 29'b0_111100101101_101_0_101111001011;
      patterns[31086] = 29'b0_111100101101_110_0_111100101101;
      patterns[31087] = 29'b0_111100101101_111_0_111100101101;
      patterns[31088] = 29'b0_111100101110_000_0_111100101110;
      patterns[31089] = 29'b0_111100101110_001_0_101110111100;
      patterns[31090] = 29'b0_111100101110_010_1_111001011100;
      patterns[31091] = 29'b0_111100101110_011_1_110010111001;
      patterns[31092] = 29'b0_111100101110_100_0_011110010111;
      patterns[31093] = 29'b0_111100101110_101_1_001111001011;
      patterns[31094] = 29'b0_111100101110_110_0_111100101110;
      patterns[31095] = 29'b0_111100101110_111_0_111100101110;
      patterns[31096] = 29'b0_111100101111_000_0_111100101111;
      patterns[31097] = 29'b0_111100101111_001_0_101111111100;
      patterns[31098] = 29'b0_111100101111_010_1_111001011110;
      patterns[31099] = 29'b0_111100101111_011_1_110010111101;
      patterns[31100] = 29'b0_111100101111_100_1_011110010111;
      patterns[31101] = 29'b0_111100101111_101_1_101111001011;
      patterns[31102] = 29'b0_111100101111_110_0_111100101111;
      patterns[31103] = 29'b0_111100101111_111_0_111100101111;
      patterns[31104] = 29'b0_111100110000_000_0_111100110000;
      patterns[31105] = 29'b0_111100110000_001_0_110000111100;
      patterns[31106] = 29'b0_111100110000_010_1_111001100000;
      patterns[31107] = 29'b0_111100110000_011_1_110011000001;
      patterns[31108] = 29'b0_111100110000_100_0_011110011000;
      patterns[31109] = 29'b0_111100110000_101_0_001111001100;
      patterns[31110] = 29'b0_111100110000_110_0_111100110000;
      patterns[31111] = 29'b0_111100110000_111_0_111100110000;
      patterns[31112] = 29'b0_111100110001_000_0_111100110001;
      patterns[31113] = 29'b0_111100110001_001_0_110001111100;
      patterns[31114] = 29'b0_111100110001_010_1_111001100010;
      patterns[31115] = 29'b0_111100110001_011_1_110011000101;
      patterns[31116] = 29'b0_111100110001_100_1_011110011000;
      patterns[31117] = 29'b0_111100110001_101_0_101111001100;
      patterns[31118] = 29'b0_111100110001_110_0_111100110001;
      patterns[31119] = 29'b0_111100110001_111_0_111100110001;
      patterns[31120] = 29'b0_111100110010_000_0_111100110010;
      patterns[31121] = 29'b0_111100110010_001_0_110010111100;
      patterns[31122] = 29'b0_111100110010_010_1_111001100100;
      patterns[31123] = 29'b0_111100110010_011_1_110011001001;
      patterns[31124] = 29'b0_111100110010_100_0_011110011001;
      patterns[31125] = 29'b0_111100110010_101_1_001111001100;
      patterns[31126] = 29'b0_111100110010_110_0_111100110010;
      patterns[31127] = 29'b0_111100110010_111_0_111100110010;
      patterns[31128] = 29'b0_111100110011_000_0_111100110011;
      patterns[31129] = 29'b0_111100110011_001_0_110011111100;
      patterns[31130] = 29'b0_111100110011_010_1_111001100110;
      patterns[31131] = 29'b0_111100110011_011_1_110011001101;
      patterns[31132] = 29'b0_111100110011_100_1_011110011001;
      patterns[31133] = 29'b0_111100110011_101_1_101111001100;
      patterns[31134] = 29'b0_111100110011_110_0_111100110011;
      patterns[31135] = 29'b0_111100110011_111_0_111100110011;
      patterns[31136] = 29'b0_111100110100_000_0_111100110100;
      patterns[31137] = 29'b0_111100110100_001_0_110100111100;
      patterns[31138] = 29'b0_111100110100_010_1_111001101000;
      patterns[31139] = 29'b0_111100110100_011_1_110011010001;
      patterns[31140] = 29'b0_111100110100_100_0_011110011010;
      patterns[31141] = 29'b0_111100110100_101_0_001111001101;
      patterns[31142] = 29'b0_111100110100_110_0_111100110100;
      patterns[31143] = 29'b0_111100110100_111_0_111100110100;
      patterns[31144] = 29'b0_111100110101_000_0_111100110101;
      patterns[31145] = 29'b0_111100110101_001_0_110101111100;
      patterns[31146] = 29'b0_111100110101_010_1_111001101010;
      patterns[31147] = 29'b0_111100110101_011_1_110011010101;
      patterns[31148] = 29'b0_111100110101_100_1_011110011010;
      patterns[31149] = 29'b0_111100110101_101_0_101111001101;
      patterns[31150] = 29'b0_111100110101_110_0_111100110101;
      patterns[31151] = 29'b0_111100110101_111_0_111100110101;
      patterns[31152] = 29'b0_111100110110_000_0_111100110110;
      patterns[31153] = 29'b0_111100110110_001_0_110110111100;
      patterns[31154] = 29'b0_111100110110_010_1_111001101100;
      patterns[31155] = 29'b0_111100110110_011_1_110011011001;
      patterns[31156] = 29'b0_111100110110_100_0_011110011011;
      patterns[31157] = 29'b0_111100110110_101_1_001111001101;
      patterns[31158] = 29'b0_111100110110_110_0_111100110110;
      patterns[31159] = 29'b0_111100110110_111_0_111100110110;
      patterns[31160] = 29'b0_111100110111_000_0_111100110111;
      patterns[31161] = 29'b0_111100110111_001_0_110111111100;
      patterns[31162] = 29'b0_111100110111_010_1_111001101110;
      patterns[31163] = 29'b0_111100110111_011_1_110011011101;
      patterns[31164] = 29'b0_111100110111_100_1_011110011011;
      patterns[31165] = 29'b0_111100110111_101_1_101111001101;
      patterns[31166] = 29'b0_111100110111_110_0_111100110111;
      patterns[31167] = 29'b0_111100110111_111_0_111100110111;
      patterns[31168] = 29'b0_111100111000_000_0_111100111000;
      patterns[31169] = 29'b0_111100111000_001_0_111000111100;
      patterns[31170] = 29'b0_111100111000_010_1_111001110000;
      patterns[31171] = 29'b0_111100111000_011_1_110011100001;
      patterns[31172] = 29'b0_111100111000_100_0_011110011100;
      patterns[31173] = 29'b0_111100111000_101_0_001111001110;
      patterns[31174] = 29'b0_111100111000_110_0_111100111000;
      patterns[31175] = 29'b0_111100111000_111_0_111100111000;
      patterns[31176] = 29'b0_111100111001_000_0_111100111001;
      patterns[31177] = 29'b0_111100111001_001_0_111001111100;
      patterns[31178] = 29'b0_111100111001_010_1_111001110010;
      patterns[31179] = 29'b0_111100111001_011_1_110011100101;
      patterns[31180] = 29'b0_111100111001_100_1_011110011100;
      patterns[31181] = 29'b0_111100111001_101_0_101111001110;
      patterns[31182] = 29'b0_111100111001_110_0_111100111001;
      patterns[31183] = 29'b0_111100111001_111_0_111100111001;
      patterns[31184] = 29'b0_111100111010_000_0_111100111010;
      patterns[31185] = 29'b0_111100111010_001_0_111010111100;
      patterns[31186] = 29'b0_111100111010_010_1_111001110100;
      patterns[31187] = 29'b0_111100111010_011_1_110011101001;
      patterns[31188] = 29'b0_111100111010_100_0_011110011101;
      patterns[31189] = 29'b0_111100111010_101_1_001111001110;
      patterns[31190] = 29'b0_111100111010_110_0_111100111010;
      patterns[31191] = 29'b0_111100111010_111_0_111100111010;
      patterns[31192] = 29'b0_111100111011_000_0_111100111011;
      patterns[31193] = 29'b0_111100111011_001_0_111011111100;
      patterns[31194] = 29'b0_111100111011_010_1_111001110110;
      patterns[31195] = 29'b0_111100111011_011_1_110011101101;
      patterns[31196] = 29'b0_111100111011_100_1_011110011101;
      patterns[31197] = 29'b0_111100111011_101_1_101111001110;
      patterns[31198] = 29'b0_111100111011_110_0_111100111011;
      patterns[31199] = 29'b0_111100111011_111_0_111100111011;
      patterns[31200] = 29'b0_111100111100_000_0_111100111100;
      patterns[31201] = 29'b0_111100111100_001_0_111100111100;
      patterns[31202] = 29'b0_111100111100_010_1_111001111000;
      patterns[31203] = 29'b0_111100111100_011_1_110011110001;
      patterns[31204] = 29'b0_111100111100_100_0_011110011110;
      patterns[31205] = 29'b0_111100111100_101_0_001111001111;
      patterns[31206] = 29'b0_111100111100_110_0_111100111100;
      patterns[31207] = 29'b0_111100111100_111_0_111100111100;
      patterns[31208] = 29'b0_111100111101_000_0_111100111101;
      patterns[31209] = 29'b0_111100111101_001_0_111101111100;
      patterns[31210] = 29'b0_111100111101_010_1_111001111010;
      patterns[31211] = 29'b0_111100111101_011_1_110011110101;
      patterns[31212] = 29'b0_111100111101_100_1_011110011110;
      patterns[31213] = 29'b0_111100111101_101_0_101111001111;
      patterns[31214] = 29'b0_111100111101_110_0_111100111101;
      patterns[31215] = 29'b0_111100111101_111_0_111100111101;
      patterns[31216] = 29'b0_111100111110_000_0_111100111110;
      patterns[31217] = 29'b0_111100111110_001_0_111110111100;
      patterns[31218] = 29'b0_111100111110_010_1_111001111100;
      patterns[31219] = 29'b0_111100111110_011_1_110011111001;
      patterns[31220] = 29'b0_111100111110_100_0_011110011111;
      patterns[31221] = 29'b0_111100111110_101_1_001111001111;
      patterns[31222] = 29'b0_111100111110_110_0_111100111110;
      patterns[31223] = 29'b0_111100111110_111_0_111100111110;
      patterns[31224] = 29'b0_111100111111_000_0_111100111111;
      patterns[31225] = 29'b0_111100111111_001_0_111111111100;
      patterns[31226] = 29'b0_111100111111_010_1_111001111110;
      patterns[31227] = 29'b0_111100111111_011_1_110011111101;
      patterns[31228] = 29'b0_111100111111_100_1_011110011111;
      patterns[31229] = 29'b0_111100111111_101_1_101111001111;
      patterns[31230] = 29'b0_111100111111_110_0_111100111111;
      patterns[31231] = 29'b0_111100111111_111_0_111100111111;
      patterns[31232] = 29'b0_111101000000_000_0_111101000000;
      patterns[31233] = 29'b0_111101000000_001_0_000000111101;
      patterns[31234] = 29'b0_111101000000_010_1_111010000000;
      patterns[31235] = 29'b0_111101000000_011_1_110100000001;
      patterns[31236] = 29'b0_111101000000_100_0_011110100000;
      patterns[31237] = 29'b0_111101000000_101_0_001111010000;
      patterns[31238] = 29'b0_111101000000_110_0_111101000000;
      patterns[31239] = 29'b0_111101000000_111_0_111101000000;
      patterns[31240] = 29'b0_111101000001_000_0_111101000001;
      patterns[31241] = 29'b0_111101000001_001_0_000001111101;
      patterns[31242] = 29'b0_111101000001_010_1_111010000010;
      patterns[31243] = 29'b0_111101000001_011_1_110100000101;
      patterns[31244] = 29'b0_111101000001_100_1_011110100000;
      patterns[31245] = 29'b0_111101000001_101_0_101111010000;
      patterns[31246] = 29'b0_111101000001_110_0_111101000001;
      patterns[31247] = 29'b0_111101000001_111_0_111101000001;
      patterns[31248] = 29'b0_111101000010_000_0_111101000010;
      patterns[31249] = 29'b0_111101000010_001_0_000010111101;
      patterns[31250] = 29'b0_111101000010_010_1_111010000100;
      patterns[31251] = 29'b0_111101000010_011_1_110100001001;
      patterns[31252] = 29'b0_111101000010_100_0_011110100001;
      patterns[31253] = 29'b0_111101000010_101_1_001111010000;
      patterns[31254] = 29'b0_111101000010_110_0_111101000010;
      patterns[31255] = 29'b0_111101000010_111_0_111101000010;
      patterns[31256] = 29'b0_111101000011_000_0_111101000011;
      patterns[31257] = 29'b0_111101000011_001_0_000011111101;
      patterns[31258] = 29'b0_111101000011_010_1_111010000110;
      patterns[31259] = 29'b0_111101000011_011_1_110100001101;
      patterns[31260] = 29'b0_111101000011_100_1_011110100001;
      patterns[31261] = 29'b0_111101000011_101_1_101111010000;
      patterns[31262] = 29'b0_111101000011_110_0_111101000011;
      patterns[31263] = 29'b0_111101000011_111_0_111101000011;
      patterns[31264] = 29'b0_111101000100_000_0_111101000100;
      patterns[31265] = 29'b0_111101000100_001_0_000100111101;
      patterns[31266] = 29'b0_111101000100_010_1_111010001000;
      patterns[31267] = 29'b0_111101000100_011_1_110100010001;
      patterns[31268] = 29'b0_111101000100_100_0_011110100010;
      patterns[31269] = 29'b0_111101000100_101_0_001111010001;
      patterns[31270] = 29'b0_111101000100_110_0_111101000100;
      patterns[31271] = 29'b0_111101000100_111_0_111101000100;
      patterns[31272] = 29'b0_111101000101_000_0_111101000101;
      patterns[31273] = 29'b0_111101000101_001_0_000101111101;
      patterns[31274] = 29'b0_111101000101_010_1_111010001010;
      patterns[31275] = 29'b0_111101000101_011_1_110100010101;
      patterns[31276] = 29'b0_111101000101_100_1_011110100010;
      patterns[31277] = 29'b0_111101000101_101_0_101111010001;
      patterns[31278] = 29'b0_111101000101_110_0_111101000101;
      patterns[31279] = 29'b0_111101000101_111_0_111101000101;
      patterns[31280] = 29'b0_111101000110_000_0_111101000110;
      patterns[31281] = 29'b0_111101000110_001_0_000110111101;
      patterns[31282] = 29'b0_111101000110_010_1_111010001100;
      patterns[31283] = 29'b0_111101000110_011_1_110100011001;
      patterns[31284] = 29'b0_111101000110_100_0_011110100011;
      patterns[31285] = 29'b0_111101000110_101_1_001111010001;
      patterns[31286] = 29'b0_111101000110_110_0_111101000110;
      patterns[31287] = 29'b0_111101000110_111_0_111101000110;
      patterns[31288] = 29'b0_111101000111_000_0_111101000111;
      patterns[31289] = 29'b0_111101000111_001_0_000111111101;
      patterns[31290] = 29'b0_111101000111_010_1_111010001110;
      patterns[31291] = 29'b0_111101000111_011_1_110100011101;
      patterns[31292] = 29'b0_111101000111_100_1_011110100011;
      patterns[31293] = 29'b0_111101000111_101_1_101111010001;
      patterns[31294] = 29'b0_111101000111_110_0_111101000111;
      patterns[31295] = 29'b0_111101000111_111_0_111101000111;
      patterns[31296] = 29'b0_111101001000_000_0_111101001000;
      patterns[31297] = 29'b0_111101001000_001_0_001000111101;
      patterns[31298] = 29'b0_111101001000_010_1_111010010000;
      patterns[31299] = 29'b0_111101001000_011_1_110100100001;
      patterns[31300] = 29'b0_111101001000_100_0_011110100100;
      patterns[31301] = 29'b0_111101001000_101_0_001111010010;
      patterns[31302] = 29'b0_111101001000_110_0_111101001000;
      patterns[31303] = 29'b0_111101001000_111_0_111101001000;
      patterns[31304] = 29'b0_111101001001_000_0_111101001001;
      patterns[31305] = 29'b0_111101001001_001_0_001001111101;
      patterns[31306] = 29'b0_111101001001_010_1_111010010010;
      patterns[31307] = 29'b0_111101001001_011_1_110100100101;
      patterns[31308] = 29'b0_111101001001_100_1_011110100100;
      patterns[31309] = 29'b0_111101001001_101_0_101111010010;
      patterns[31310] = 29'b0_111101001001_110_0_111101001001;
      patterns[31311] = 29'b0_111101001001_111_0_111101001001;
      patterns[31312] = 29'b0_111101001010_000_0_111101001010;
      patterns[31313] = 29'b0_111101001010_001_0_001010111101;
      patterns[31314] = 29'b0_111101001010_010_1_111010010100;
      patterns[31315] = 29'b0_111101001010_011_1_110100101001;
      patterns[31316] = 29'b0_111101001010_100_0_011110100101;
      patterns[31317] = 29'b0_111101001010_101_1_001111010010;
      patterns[31318] = 29'b0_111101001010_110_0_111101001010;
      patterns[31319] = 29'b0_111101001010_111_0_111101001010;
      patterns[31320] = 29'b0_111101001011_000_0_111101001011;
      patterns[31321] = 29'b0_111101001011_001_0_001011111101;
      patterns[31322] = 29'b0_111101001011_010_1_111010010110;
      patterns[31323] = 29'b0_111101001011_011_1_110100101101;
      patterns[31324] = 29'b0_111101001011_100_1_011110100101;
      patterns[31325] = 29'b0_111101001011_101_1_101111010010;
      patterns[31326] = 29'b0_111101001011_110_0_111101001011;
      patterns[31327] = 29'b0_111101001011_111_0_111101001011;
      patterns[31328] = 29'b0_111101001100_000_0_111101001100;
      patterns[31329] = 29'b0_111101001100_001_0_001100111101;
      patterns[31330] = 29'b0_111101001100_010_1_111010011000;
      patterns[31331] = 29'b0_111101001100_011_1_110100110001;
      patterns[31332] = 29'b0_111101001100_100_0_011110100110;
      patterns[31333] = 29'b0_111101001100_101_0_001111010011;
      patterns[31334] = 29'b0_111101001100_110_0_111101001100;
      patterns[31335] = 29'b0_111101001100_111_0_111101001100;
      patterns[31336] = 29'b0_111101001101_000_0_111101001101;
      patterns[31337] = 29'b0_111101001101_001_0_001101111101;
      patterns[31338] = 29'b0_111101001101_010_1_111010011010;
      patterns[31339] = 29'b0_111101001101_011_1_110100110101;
      patterns[31340] = 29'b0_111101001101_100_1_011110100110;
      patterns[31341] = 29'b0_111101001101_101_0_101111010011;
      patterns[31342] = 29'b0_111101001101_110_0_111101001101;
      patterns[31343] = 29'b0_111101001101_111_0_111101001101;
      patterns[31344] = 29'b0_111101001110_000_0_111101001110;
      patterns[31345] = 29'b0_111101001110_001_0_001110111101;
      patterns[31346] = 29'b0_111101001110_010_1_111010011100;
      patterns[31347] = 29'b0_111101001110_011_1_110100111001;
      patterns[31348] = 29'b0_111101001110_100_0_011110100111;
      patterns[31349] = 29'b0_111101001110_101_1_001111010011;
      patterns[31350] = 29'b0_111101001110_110_0_111101001110;
      patterns[31351] = 29'b0_111101001110_111_0_111101001110;
      patterns[31352] = 29'b0_111101001111_000_0_111101001111;
      patterns[31353] = 29'b0_111101001111_001_0_001111111101;
      patterns[31354] = 29'b0_111101001111_010_1_111010011110;
      patterns[31355] = 29'b0_111101001111_011_1_110100111101;
      patterns[31356] = 29'b0_111101001111_100_1_011110100111;
      patterns[31357] = 29'b0_111101001111_101_1_101111010011;
      patterns[31358] = 29'b0_111101001111_110_0_111101001111;
      patterns[31359] = 29'b0_111101001111_111_0_111101001111;
      patterns[31360] = 29'b0_111101010000_000_0_111101010000;
      patterns[31361] = 29'b0_111101010000_001_0_010000111101;
      patterns[31362] = 29'b0_111101010000_010_1_111010100000;
      patterns[31363] = 29'b0_111101010000_011_1_110101000001;
      patterns[31364] = 29'b0_111101010000_100_0_011110101000;
      patterns[31365] = 29'b0_111101010000_101_0_001111010100;
      patterns[31366] = 29'b0_111101010000_110_0_111101010000;
      patterns[31367] = 29'b0_111101010000_111_0_111101010000;
      patterns[31368] = 29'b0_111101010001_000_0_111101010001;
      patterns[31369] = 29'b0_111101010001_001_0_010001111101;
      patterns[31370] = 29'b0_111101010001_010_1_111010100010;
      patterns[31371] = 29'b0_111101010001_011_1_110101000101;
      patterns[31372] = 29'b0_111101010001_100_1_011110101000;
      patterns[31373] = 29'b0_111101010001_101_0_101111010100;
      patterns[31374] = 29'b0_111101010001_110_0_111101010001;
      patterns[31375] = 29'b0_111101010001_111_0_111101010001;
      patterns[31376] = 29'b0_111101010010_000_0_111101010010;
      patterns[31377] = 29'b0_111101010010_001_0_010010111101;
      patterns[31378] = 29'b0_111101010010_010_1_111010100100;
      patterns[31379] = 29'b0_111101010010_011_1_110101001001;
      patterns[31380] = 29'b0_111101010010_100_0_011110101001;
      patterns[31381] = 29'b0_111101010010_101_1_001111010100;
      patterns[31382] = 29'b0_111101010010_110_0_111101010010;
      patterns[31383] = 29'b0_111101010010_111_0_111101010010;
      patterns[31384] = 29'b0_111101010011_000_0_111101010011;
      patterns[31385] = 29'b0_111101010011_001_0_010011111101;
      patterns[31386] = 29'b0_111101010011_010_1_111010100110;
      patterns[31387] = 29'b0_111101010011_011_1_110101001101;
      patterns[31388] = 29'b0_111101010011_100_1_011110101001;
      patterns[31389] = 29'b0_111101010011_101_1_101111010100;
      patterns[31390] = 29'b0_111101010011_110_0_111101010011;
      patterns[31391] = 29'b0_111101010011_111_0_111101010011;
      patterns[31392] = 29'b0_111101010100_000_0_111101010100;
      patterns[31393] = 29'b0_111101010100_001_0_010100111101;
      patterns[31394] = 29'b0_111101010100_010_1_111010101000;
      patterns[31395] = 29'b0_111101010100_011_1_110101010001;
      patterns[31396] = 29'b0_111101010100_100_0_011110101010;
      patterns[31397] = 29'b0_111101010100_101_0_001111010101;
      patterns[31398] = 29'b0_111101010100_110_0_111101010100;
      patterns[31399] = 29'b0_111101010100_111_0_111101010100;
      patterns[31400] = 29'b0_111101010101_000_0_111101010101;
      patterns[31401] = 29'b0_111101010101_001_0_010101111101;
      patterns[31402] = 29'b0_111101010101_010_1_111010101010;
      patterns[31403] = 29'b0_111101010101_011_1_110101010101;
      patterns[31404] = 29'b0_111101010101_100_1_011110101010;
      patterns[31405] = 29'b0_111101010101_101_0_101111010101;
      patterns[31406] = 29'b0_111101010101_110_0_111101010101;
      patterns[31407] = 29'b0_111101010101_111_0_111101010101;
      patterns[31408] = 29'b0_111101010110_000_0_111101010110;
      patterns[31409] = 29'b0_111101010110_001_0_010110111101;
      patterns[31410] = 29'b0_111101010110_010_1_111010101100;
      patterns[31411] = 29'b0_111101010110_011_1_110101011001;
      patterns[31412] = 29'b0_111101010110_100_0_011110101011;
      patterns[31413] = 29'b0_111101010110_101_1_001111010101;
      patterns[31414] = 29'b0_111101010110_110_0_111101010110;
      patterns[31415] = 29'b0_111101010110_111_0_111101010110;
      patterns[31416] = 29'b0_111101010111_000_0_111101010111;
      patterns[31417] = 29'b0_111101010111_001_0_010111111101;
      patterns[31418] = 29'b0_111101010111_010_1_111010101110;
      patterns[31419] = 29'b0_111101010111_011_1_110101011101;
      patterns[31420] = 29'b0_111101010111_100_1_011110101011;
      patterns[31421] = 29'b0_111101010111_101_1_101111010101;
      patterns[31422] = 29'b0_111101010111_110_0_111101010111;
      patterns[31423] = 29'b0_111101010111_111_0_111101010111;
      patterns[31424] = 29'b0_111101011000_000_0_111101011000;
      patterns[31425] = 29'b0_111101011000_001_0_011000111101;
      patterns[31426] = 29'b0_111101011000_010_1_111010110000;
      patterns[31427] = 29'b0_111101011000_011_1_110101100001;
      patterns[31428] = 29'b0_111101011000_100_0_011110101100;
      patterns[31429] = 29'b0_111101011000_101_0_001111010110;
      patterns[31430] = 29'b0_111101011000_110_0_111101011000;
      patterns[31431] = 29'b0_111101011000_111_0_111101011000;
      patterns[31432] = 29'b0_111101011001_000_0_111101011001;
      patterns[31433] = 29'b0_111101011001_001_0_011001111101;
      patterns[31434] = 29'b0_111101011001_010_1_111010110010;
      patterns[31435] = 29'b0_111101011001_011_1_110101100101;
      patterns[31436] = 29'b0_111101011001_100_1_011110101100;
      patterns[31437] = 29'b0_111101011001_101_0_101111010110;
      patterns[31438] = 29'b0_111101011001_110_0_111101011001;
      patterns[31439] = 29'b0_111101011001_111_0_111101011001;
      patterns[31440] = 29'b0_111101011010_000_0_111101011010;
      patterns[31441] = 29'b0_111101011010_001_0_011010111101;
      patterns[31442] = 29'b0_111101011010_010_1_111010110100;
      patterns[31443] = 29'b0_111101011010_011_1_110101101001;
      patterns[31444] = 29'b0_111101011010_100_0_011110101101;
      patterns[31445] = 29'b0_111101011010_101_1_001111010110;
      patterns[31446] = 29'b0_111101011010_110_0_111101011010;
      patterns[31447] = 29'b0_111101011010_111_0_111101011010;
      patterns[31448] = 29'b0_111101011011_000_0_111101011011;
      patterns[31449] = 29'b0_111101011011_001_0_011011111101;
      patterns[31450] = 29'b0_111101011011_010_1_111010110110;
      patterns[31451] = 29'b0_111101011011_011_1_110101101101;
      patterns[31452] = 29'b0_111101011011_100_1_011110101101;
      patterns[31453] = 29'b0_111101011011_101_1_101111010110;
      patterns[31454] = 29'b0_111101011011_110_0_111101011011;
      patterns[31455] = 29'b0_111101011011_111_0_111101011011;
      patterns[31456] = 29'b0_111101011100_000_0_111101011100;
      patterns[31457] = 29'b0_111101011100_001_0_011100111101;
      patterns[31458] = 29'b0_111101011100_010_1_111010111000;
      patterns[31459] = 29'b0_111101011100_011_1_110101110001;
      patterns[31460] = 29'b0_111101011100_100_0_011110101110;
      patterns[31461] = 29'b0_111101011100_101_0_001111010111;
      patterns[31462] = 29'b0_111101011100_110_0_111101011100;
      patterns[31463] = 29'b0_111101011100_111_0_111101011100;
      patterns[31464] = 29'b0_111101011101_000_0_111101011101;
      patterns[31465] = 29'b0_111101011101_001_0_011101111101;
      patterns[31466] = 29'b0_111101011101_010_1_111010111010;
      patterns[31467] = 29'b0_111101011101_011_1_110101110101;
      patterns[31468] = 29'b0_111101011101_100_1_011110101110;
      patterns[31469] = 29'b0_111101011101_101_0_101111010111;
      patterns[31470] = 29'b0_111101011101_110_0_111101011101;
      patterns[31471] = 29'b0_111101011101_111_0_111101011101;
      patterns[31472] = 29'b0_111101011110_000_0_111101011110;
      patterns[31473] = 29'b0_111101011110_001_0_011110111101;
      patterns[31474] = 29'b0_111101011110_010_1_111010111100;
      patterns[31475] = 29'b0_111101011110_011_1_110101111001;
      patterns[31476] = 29'b0_111101011110_100_0_011110101111;
      patterns[31477] = 29'b0_111101011110_101_1_001111010111;
      patterns[31478] = 29'b0_111101011110_110_0_111101011110;
      patterns[31479] = 29'b0_111101011110_111_0_111101011110;
      patterns[31480] = 29'b0_111101011111_000_0_111101011111;
      patterns[31481] = 29'b0_111101011111_001_0_011111111101;
      patterns[31482] = 29'b0_111101011111_010_1_111010111110;
      patterns[31483] = 29'b0_111101011111_011_1_110101111101;
      patterns[31484] = 29'b0_111101011111_100_1_011110101111;
      patterns[31485] = 29'b0_111101011111_101_1_101111010111;
      patterns[31486] = 29'b0_111101011111_110_0_111101011111;
      patterns[31487] = 29'b0_111101011111_111_0_111101011111;
      patterns[31488] = 29'b0_111101100000_000_0_111101100000;
      patterns[31489] = 29'b0_111101100000_001_0_100000111101;
      patterns[31490] = 29'b0_111101100000_010_1_111011000000;
      patterns[31491] = 29'b0_111101100000_011_1_110110000001;
      patterns[31492] = 29'b0_111101100000_100_0_011110110000;
      patterns[31493] = 29'b0_111101100000_101_0_001111011000;
      patterns[31494] = 29'b0_111101100000_110_0_111101100000;
      patterns[31495] = 29'b0_111101100000_111_0_111101100000;
      patterns[31496] = 29'b0_111101100001_000_0_111101100001;
      patterns[31497] = 29'b0_111101100001_001_0_100001111101;
      patterns[31498] = 29'b0_111101100001_010_1_111011000010;
      patterns[31499] = 29'b0_111101100001_011_1_110110000101;
      patterns[31500] = 29'b0_111101100001_100_1_011110110000;
      patterns[31501] = 29'b0_111101100001_101_0_101111011000;
      patterns[31502] = 29'b0_111101100001_110_0_111101100001;
      patterns[31503] = 29'b0_111101100001_111_0_111101100001;
      patterns[31504] = 29'b0_111101100010_000_0_111101100010;
      patterns[31505] = 29'b0_111101100010_001_0_100010111101;
      patterns[31506] = 29'b0_111101100010_010_1_111011000100;
      patterns[31507] = 29'b0_111101100010_011_1_110110001001;
      patterns[31508] = 29'b0_111101100010_100_0_011110110001;
      patterns[31509] = 29'b0_111101100010_101_1_001111011000;
      patterns[31510] = 29'b0_111101100010_110_0_111101100010;
      patterns[31511] = 29'b0_111101100010_111_0_111101100010;
      patterns[31512] = 29'b0_111101100011_000_0_111101100011;
      patterns[31513] = 29'b0_111101100011_001_0_100011111101;
      patterns[31514] = 29'b0_111101100011_010_1_111011000110;
      patterns[31515] = 29'b0_111101100011_011_1_110110001101;
      patterns[31516] = 29'b0_111101100011_100_1_011110110001;
      patterns[31517] = 29'b0_111101100011_101_1_101111011000;
      patterns[31518] = 29'b0_111101100011_110_0_111101100011;
      patterns[31519] = 29'b0_111101100011_111_0_111101100011;
      patterns[31520] = 29'b0_111101100100_000_0_111101100100;
      patterns[31521] = 29'b0_111101100100_001_0_100100111101;
      patterns[31522] = 29'b0_111101100100_010_1_111011001000;
      patterns[31523] = 29'b0_111101100100_011_1_110110010001;
      patterns[31524] = 29'b0_111101100100_100_0_011110110010;
      patterns[31525] = 29'b0_111101100100_101_0_001111011001;
      patterns[31526] = 29'b0_111101100100_110_0_111101100100;
      patterns[31527] = 29'b0_111101100100_111_0_111101100100;
      patterns[31528] = 29'b0_111101100101_000_0_111101100101;
      patterns[31529] = 29'b0_111101100101_001_0_100101111101;
      patterns[31530] = 29'b0_111101100101_010_1_111011001010;
      patterns[31531] = 29'b0_111101100101_011_1_110110010101;
      patterns[31532] = 29'b0_111101100101_100_1_011110110010;
      patterns[31533] = 29'b0_111101100101_101_0_101111011001;
      patterns[31534] = 29'b0_111101100101_110_0_111101100101;
      patterns[31535] = 29'b0_111101100101_111_0_111101100101;
      patterns[31536] = 29'b0_111101100110_000_0_111101100110;
      patterns[31537] = 29'b0_111101100110_001_0_100110111101;
      patterns[31538] = 29'b0_111101100110_010_1_111011001100;
      patterns[31539] = 29'b0_111101100110_011_1_110110011001;
      patterns[31540] = 29'b0_111101100110_100_0_011110110011;
      patterns[31541] = 29'b0_111101100110_101_1_001111011001;
      patterns[31542] = 29'b0_111101100110_110_0_111101100110;
      patterns[31543] = 29'b0_111101100110_111_0_111101100110;
      patterns[31544] = 29'b0_111101100111_000_0_111101100111;
      patterns[31545] = 29'b0_111101100111_001_0_100111111101;
      patterns[31546] = 29'b0_111101100111_010_1_111011001110;
      patterns[31547] = 29'b0_111101100111_011_1_110110011101;
      patterns[31548] = 29'b0_111101100111_100_1_011110110011;
      patterns[31549] = 29'b0_111101100111_101_1_101111011001;
      patterns[31550] = 29'b0_111101100111_110_0_111101100111;
      patterns[31551] = 29'b0_111101100111_111_0_111101100111;
      patterns[31552] = 29'b0_111101101000_000_0_111101101000;
      patterns[31553] = 29'b0_111101101000_001_0_101000111101;
      patterns[31554] = 29'b0_111101101000_010_1_111011010000;
      patterns[31555] = 29'b0_111101101000_011_1_110110100001;
      patterns[31556] = 29'b0_111101101000_100_0_011110110100;
      patterns[31557] = 29'b0_111101101000_101_0_001111011010;
      patterns[31558] = 29'b0_111101101000_110_0_111101101000;
      patterns[31559] = 29'b0_111101101000_111_0_111101101000;
      patterns[31560] = 29'b0_111101101001_000_0_111101101001;
      patterns[31561] = 29'b0_111101101001_001_0_101001111101;
      patterns[31562] = 29'b0_111101101001_010_1_111011010010;
      patterns[31563] = 29'b0_111101101001_011_1_110110100101;
      patterns[31564] = 29'b0_111101101001_100_1_011110110100;
      patterns[31565] = 29'b0_111101101001_101_0_101111011010;
      patterns[31566] = 29'b0_111101101001_110_0_111101101001;
      patterns[31567] = 29'b0_111101101001_111_0_111101101001;
      patterns[31568] = 29'b0_111101101010_000_0_111101101010;
      patterns[31569] = 29'b0_111101101010_001_0_101010111101;
      patterns[31570] = 29'b0_111101101010_010_1_111011010100;
      patterns[31571] = 29'b0_111101101010_011_1_110110101001;
      patterns[31572] = 29'b0_111101101010_100_0_011110110101;
      patterns[31573] = 29'b0_111101101010_101_1_001111011010;
      patterns[31574] = 29'b0_111101101010_110_0_111101101010;
      patterns[31575] = 29'b0_111101101010_111_0_111101101010;
      patterns[31576] = 29'b0_111101101011_000_0_111101101011;
      patterns[31577] = 29'b0_111101101011_001_0_101011111101;
      patterns[31578] = 29'b0_111101101011_010_1_111011010110;
      patterns[31579] = 29'b0_111101101011_011_1_110110101101;
      patterns[31580] = 29'b0_111101101011_100_1_011110110101;
      patterns[31581] = 29'b0_111101101011_101_1_101111011010;
      patterns[31582] = 29'b0_111101101011_110_0_111101101011;
      patterns[31583] = 29'b0_111101101011_111_0_111101101011;
      patterns[31584] = 29'b0_111101101100_000_0_111101101100;
      patterns[31585] = 29'b0_111101101100_001_0_101100111101;
      patterns[31586] = 29'b0_111101101100_010_1_111011011000;
      patterns[31587] = 29'b0_111101101100_011_1_110110110001;
      patterns[31588] = 29'b0_111101101100_100_0_011110110110;
      patterns[31589] = 29'b0_111101101100_101_0_001111011011;
      patterns[31590] = 29'b0_111101101100_110_0_111101101100;
      patterns[31591] = 29'b0_111101101100_111_0_111101101100;
      patterns[31592] = 29'b0_111101101101_000_0_111101101101;
      patterns[31593] = 29'b0_111101101101_001_0_101101111101;
      patterns[31594] = 29'b0_111101101101_010_1_111011011010;
      patterns[31595] = 29'b0_111101101101_011_1_110110110101;
      patterns[31596] = 29'b0_111101101101_100_1_011110110110;
      patterns[31597] = 29'b0_111101101101_101_0_101111011011;
      patterns[31598] = 29'b0_111101101101_110_0_111101101101;
      patterns[31599] = 29'b0_111101101101_111_0_111101101101;
      patterns[31600] = 29'b0_111101101110_000_0_111101101110;
      patterns[31601] = 29'b0_111101101110_001_0_101110111101;
      patterns[31602] = 29'b0_111101101110_010_1_111011011100;
      patterns[31603] = 29'b0_111101101110_011_1_110110111001;
      patterns[31604] = 29'b0_111101101110_100_0_011110110111;
      patterns[31605] = 29'b0_111101101110_101_1_001111011011;
      patterns[31606] = 29'b0_111101101110_110_0_111101101110;
      patterns[31607] = 29'b0_111101101110_111_0_111101101110;
      patterns[31608] = 29'b0_111101101111_000_0_111101101111;
      patterns[31609] = 29'b0_111101101111_001_0_101111111101;
      patterns[31610] = 29'b0_111101101111_010_1_111011011110;
      patterns[31611] = 29'b0_111101101111_011_1_110110111101;
      patterns[31612] = 29'b0_111101101111_100_1_011110110111;
      patterns[31613] = 29'b0_111101101111_101_1_101111011011;
      patterns[31614] = 29'b0_111101101111_110_0_111101101111;
      patterns[31615] = 29'b0_111101101111_111_0_111101101111;
      patterns[31616] = 29'b0_111101110000_000_0_111101110000;
      patterns[31617] = 29'b0_111101110000_001_0_110000111101;
      patterns[31618] = 29'b0_111101110000_010_1_111011100000;
      patterns[31619] = 29'b0_111101110000_011_1_110111000001;
      patterns[31620] = 29'b0_111101110000_100_0_011110111000;
      patterns[31621] = 29'b0_111101110000_101_0_001111011100;
      patterns[31622] = 29'b0_111101110000_110_0_111101110000;
      patterns[31623] = 29'b0_111101110000_111_0_111101110000;
      patterns[31624] = 29'b0_111101110001_000_0_111101110001;
      patterns[31625] = 29'b0_111101110001_001_0_110001111101;
      patterns[31626] = 29'b0_111101110001_010_1_111011100010;
      patterns[31627] = 29'b0_111101110001_011_1_110111000101;
      patterns[31628] = 29'b0_111101110001_100_1_011110111000;
      patterns[31629] = 29'b0_111101110001_101_0_101111011100;
      patterns[31630] = 29'b0_111101110001_110_0_111101110001;
      patterns[31631] = 29'b0_111101110001_111_0_111101110001;
      patterns[31632] = 29'b0_111101110010_000_0_111101110010;
      patterns[31633] = 29'b0_111101110010_001_0_110010111101;
      patterns[31634] = 29'b0_111101110010_010_1_111011100100;
      patterns[31635] = 29'b0_111101110010_011_1_110111001001;
      patterns[31636] = 29'b0_111101110010_100_0_011110111001;
      patterns[31637] = 29'b0_111101110010_101_1_001111011100;
      patterns[31638] = 29'b0_111101110010_110_0_111101110010;
      patterns[31639] = 29'b0_111101110010_111_0_111101110010;
      patterns[31640] = 29'b0_111101110011_000_0_111101110011;
      patterns[31641] = 29'b0_111101110011_001_0_110011111101;
      patterns[31642] = 29'b0_111101110011_010_1_111011100110;
      patterns[31643] = 29'b0_111101110011_011_1_110111001101;
      patterns[31644] = 29'b0_111101110011_100_1_011110111001;
      patterns[31645] = 29'b0_111101110011_101_1_101111011100;
      patterns[31646] = 29'b0_111101110011_110_0_111101110011;
      patterns[31647] = 29'b0_111101110011_111_0_111101110011;
      patterns[31648] = 29'b0_111101110100_000_0_111101110100;
      patterns[31649] = 29'b0_111101110100_001_0_110100111101;
      patterns[31650] = 29'b0_111101110100_010_1_111011101000;
      patterns[31651] = 29'b0_111101110100_011_1_110111010001;
      patterns[31652] = 29'b0_111101110100_100_0_011110111010;
      patterns[31653] = 29'b0_111101110100_101_0_001111011101;
      patterns[31654] = 29'b0_111101110100_110_0_111101110100;
      patterns[31655] = 29'b0_111101110100_111_0_111101110100;
      patterns[31656] = 29'b0_111101110101_000_0_111101110101;
      patterns[31657] = 29'b0_111101110101_001_0_110101111101;
      patterns[31658] = 29'b0_111101110101_010_1_111011101010;
      patterns[31659] = 29'b0_111101110101_011_1_110111010101;
      patterns[31660] = 29'b0_111101110101_100_1_011110111010;
      patterns[31661] = 29'b0_111101110101_101_0_101111011101;
      patterns[31662] = 29'b0_111101110101_110_0_111101110101;
      patterns[31663] = 29'b0_111101110101_111_0_111101110101;
      patterns[31664] = 29'b0_111101110110_000_0_111101110110;
      patterns[31665] = 29'b0_111101110110_001_0_110110111101;
      patterns[31666] = 29'b0_111101110110_010_1_111011101100;
      patterns[31667] = 29'b0_111101110110_011_1_110111011001;
      patterns[31668] = 29'b0_111101110110_100_0_011110111011;
      patterns[31669] = 29'b0_111101110110_101_1_001111011101;
      patterns[31670] = 29'b0_111101110110_110_0_111101110110;
      patterns[31671] = 29'b0_111101110110_111_0_111101110110;
      patterns[31672] = 29'b0_111101110111_000_0_111101110111;
      patterns[31673] = 29'b0_111101110111_001_0_110111111101;
      patterns[31674] = 29'b0_111101110111_010_1_111011101110;
      patterns[31675] = 29'b0_111101110111_011_1_110111011101;
      patterns[31676] = 29'b0_111101110111_100_1_011110111011;
      patterns[31677] = 29'b0_111101110111_101_1_101111011101;
      patterns[31678] = 29'b0_111101110111_110_0_111101110111;
      patterns[31679] = 29'b0_111101110111_111_0_111101110111;
      patterns[31680] = 29'b0_111101111000_000_0_111101111000;
      patterns[31681] = 29'b0_111101111000_001_0_111000111101;
      patterns[31682] = 29'b0_111101111000_010_1_111011110000;
      patterns[31683] = 29'b0_111101111000_011_1_110111100001;
      patterns[31684] = 29'b0_111101111000_100_0_011110111100;
      patterns[31685] = 29'b0_111101111000_101_0_001111011110;
      patterns[31686] = 29'b0_111101111000_110_0_111101111000;
      patterns[31687] = 29'b0_111101111000_111_0_111101111000;
      patterns[31688] = 29'b0_111101111001_000_0_111101111001;
      patterns[31689] = 29'b0_111101111001_001_0_111001111101;
      patterns[31690] = 29'b0_111101111001_010_1_111011110010;
      patterns[31691] = 29'b0_111101111001_011_1_110111100101;
      patterns[31692] = 29'b0_111101111001_100_1_011110111100;
      patterns[31693] = 29'b0_111101111001_101_0_101111011110;
      patterns[31694] = 29'b0_111101111001_110_0_111101111001;
      patterns[31695] = 29'b0_111101111001_111_0_111101111001;
      patterns[31696] = 29'b0_111101111010_000_0_111101111010;
      patterns[31697] = 29'b0_111101111010_001_0_111010111101;
      patterns[31698] = 29'b0_111101111010_010_1_111011110100;
      patterns[31699] = 29'b0_111101111010_011_1_110111101001;
      patterns[31700] = 29'b0_111101111010_100_0_011110111101;
      patterns[31701] = 29'b0_111101111010_101_1_001111011110;
      patterns[31702] = 29'b0_111101111010_110_0_111101111010;
      patterns[31703] = 29'b0_111101111010_111_0_111101111010;
      patterns[31704] = 29'b0_111101111011_000_0_111101111011;
      patterns[31705] = 29'b0_111101111011_001_0_111011111101;
      patterns[31706] = 29'b0_111101111011_010_1_111011110110;
      patterns[31707] = 29'b0_111101111011_011_1_110111101101;
      patterns[31708] = 29'b0_111101111011_100_1_011110111101;
      patterns[31709] = 29'b0_111101111011_101_1_101111011110;
      patterns[31710] = 29'b0_111101111011_110_0_111101111011;
      patterns[31711] = 29'b0_111101111011_111_0_111101111011;
      patterns[31712] = 29'b0_111101111100_000_0_111101111100;
      patterns[31713] = 29'b0_111101111100_001_0_111100111101;
      patterns[31714] = 29'b0_111101111100_010_1_111011111000;
      patterns[31715] = 29'b0_111101111100_011_1_110111110001;
      patterns[31716] = 29'b0_111101111100_100_0_011110111110;
      patterns[31717] = 29'b0_111101111100_101_0_001111011111;
      patterns[31718] = 29'b0_111101111100_110_0_111101111100;
      patterns[31719] = 29'b0_111101111100_111_0_111101111100;
      patterns[31720] = 29'b0_111101111101_000_0_111101111101;
      patterns[31721] = 29'b0_111101111101_001_0_111101111101;
      patterns[31722] = 29'b0_111101111101_010_1_111011111010;
      patterns[31723] = 29'b0_111101111101_011_1_110111110101;
      patterns[31724] = 29'b0_111101111101_100_1_011110111110;
      patterns[31725] = 29'b0_111101111101_101_0_101111011111;
      patterns[31726] = 29'b0_111101111101_110_0_111101111101;
      patterns[31727] = 29'b0_111101111101_111_0_111101111101;
      patterns[31728] = 29'b0_111101111110_000_0_111101111110;
      patterns[31729] = 29'b0_111101111110_001_0_111110111101;
      patterns[31730] = 29'b0_111101111110_010_1_111011111100;
      patterns[31731] = 29'b0_111101111110_011_1_110111111001;
      patterns[31732] = 29'b0_111101111110_100_0_011110111111;
      patterns[31733] = 29'b0_111101111110_101_1_001111011111;
      patterns[31734] = 29'b0_111101111110_110_0_111101111110;
      patterns[31735] = 29'b0_111101111110_111_0_111101111110;
      patterns[31736] = 29'b0_111101111111_000_0_111101111111;
      patterns[31737] = 29'b0_111101111111_001_0_111111111101;
      patterns[31738] = 29'b0_111101111111_010_1_111011111110;
      patterns[31739] = 29'b0_111101111111_011_1_110111111101;
      patterns[31740] = 29'b0_111101111111_100_1_011110111111;
      patterns[31741] = 29'b0_111101111111_101_1_101111011111;
      patterns[31742] = 29'b0_111101111111_110_0_111101111111;
      patterns[31743] = 29'b0_111101111111_111_0_111101111111;
      patterns[31744] = 29'b0_111110000000_000_0_111110000000;
      patterns[31745] = 29'b0_111110000000_001_0_000000111110;
      patterns[31746] = 29'b0_111110000000_010_1_111100000000;
      patterns[31747] = 29'b0_111110000000_011_1_111000000001;
      patterns[31748] = 29'b0_111110000000_100_0_011111000000;
      patterns[31749] = 29'b0_111110000000_101_0_001111100000;
      patterns[31750] = 29'b0_111110000000_110_0_111110000000;
      patterns[31751] = 29'b0_111110000000_111_0_111110000000;
      patterns[31752] = 29'b0_111110000001_000_0_111110000001;
      patterns[31753] = 29'b0_111110000001_001_0_000001111110;
      patterns[31754] = 29'b0_111110000001_010_1_111100000010;
      patterns[31755] = 29'b0_111110000001_011_1_111000000101;
      patterns[31756] = 29'b0_111110000001_100_1_011111000000;
      patterns[31757] = 29'b0_111110000001_101_0_101111100000;
      patterns[31758] = 29'b0_111110000001_110_0_111110000001;
      patterns[31759] = 29'b0_111110000001_111_0_111110000001;
      patterns[31760] = 29'b0_111110000010_000_0_111110000010;
      patterns[31761] = 29'b0_111110000010_001_0_000010111110;
      patterns[31762] = 29'b0_111110000010_010_1_111100000100;
      patterns[31763] = 29'b0_111110000010_011_1_111000001001;
      patterns[31764] = 29'b0_111110000010_100_0_011111000001;
      patterns[31765] = 29'b0_111110000010_101_1_001111100000;
      patterns[31766] = 29'b0_111110000010_110_0_111110000010;
      patterns[31767] = 29'b0_111110000010_111_0_111110000010;
      patterns[31768] = 29'b0_111110000011_000_0_111110000011;
      patterns[31769] = 29'b0_111110000011_001_0_000011111110;
      patterns[31770] = 29'b0_111110000011_010_1_111100000110;
      patterns[31771] = 29'b0_111110000011_011_1_111000001101;
      patterns[31772] = 29'b0_111110000011_100_1_011111000001;
      patterns[31773] = 29'b0_111110000011_101_1_101111100000;
      patterns[31774] = 29'b0_111110000011_110_0_111110000011;
      patterns[31775] = 29'b0_111110000011_111_0_111110000011;
      patterns[31776] = 29'b0_111110000100_000_0_111110000100;
      patterns[31777] = 29'b0_111110000100_001_0_000100111110;
      patterns[31778] = 29'b0_111110000100_010_1_111100001000;
      patterns[31779] = 29'b0_111110000100_011_1_111000010001;
      patterns[31780] = 29'b0_111110000100_100_0_011111000010;
      patterns[31781] = 29'b0_111110000100_101_0_001111100001;
      patterns[31782] = 29'b0_111110000100_110_0_111110000100;
      patterns[31783] = 29'b0_111110000100_111_0_111110000100;
      patterns[31784] = 29'b0_111110000101_000_0_111110000101;
      patterns[31785] = 29'b0_111110000101_001_0_000101111110;
      patterns[31786] = 29'b0_111110000101_010_1_111100001010;
      patterns[31787] = 29'b0_111110000101_011_1_111000010101;
      patterns[31788] = 29'b0_111110000101_100_1_011111000010;
      patterns[31789] = 29'b0_111110000101_101_0_101111100001;
      patterns[31790] = 29'b0_111110000101_110_0_111110000101;
      patterns[31791] = 29'b0_111110000101_111_0_111110000101;
      patterns[31792] = 29'b0_111110000110_000_0_111110000110;
      patterns[31793] = 29'b0_111110000110_001_0_000110111110;
      patterns[31794] = 29'b0_111110000110_010_1_111100001100;
      patterns[31795] = 29'b0_111110000110_011_1_111000011001;
      patterns[31796] = 29'b0_111110000110_100_0_011111000011;
      patterns[31797] = 29'b0_111110000110_101_1_001111100001;
      patterns[31798] = 29'b0_111110000110_110_0_111110000110;
      patterns[31799] = 29'b0_111110000110_111_0_111110000110;
      patterns[31800] = 29'b0_111110000111_000_0_111110000111;
      patterns[31801] = 29'b0_111110000111_001_0_000111111110;
      patterns[31802] = 29'b0_111110000111_010_1_111100001110;
      patterns[31803] = 29'b0_111110000111_011_1_111000011101;
      patterns[31804] = 29'b0_111110000111_100_1_011111000011;
      patterns[31805] = 29'b0_111110000111_101_1_101111100001;
      patterns[31806] = 29'b0_111110000111_110_0_111110000111;
      patterns[31807] = 29'b0_111110000111_111_0_111110000111;
      patterns[31808] = 29'b0_111110001000_000_0_111110001000;
      patterns[31809] = 29'b0_111110001000_001_0_001000111110;
      patterns[31810] = 29'b0_111110001000_010_1_111100010000;
      patterns[31811] = 29'b0_111110001000_011_1_111000100001;
      patterns[31812] = 29'b0_111110001000_100_0_011111000100;
      patterns[31813] = 29'b0_111110001000_101_0_001111100010;
      patterns[31814] = 29'b0_111110001000_110_0_111110001000;
      patterns[31815] = 29'b0_111110001000_111_0_111110001000;
      patterns[31816] = 29'b0_111110001001_000_0_111110001001;
      patterns[31817] = 29'b0_111110001001_001_0_001001111110;
      patterns[31818] = 29'b0_111110001001_010_1_111100010010;
      patterns[31819] = 29'b0_111110001001_011_1_111000100101;
      patterns[31820] = 29'b0_111110001001_100_1_011111000100;
      patterns[31821] = 29'b0_111110001001_101_0_101111100010;
      patterns[31822] = 29'b0_111110001001_110_0_111110001001;
      patterns[31823] = 29'b0_111110001001_111_0_111110001001;
      patterns[31824] = 29'b0_111110001010_000_0_111110001010;
      patterns[31825] = 29'b0_111110001010_001_0_001010111110;
      patterns[31826] = 29'b0_111110001010_010_1_111100010100;
      patterns[31827] = 29'b0_111110001010_011_1_111000101001;
      patterns[31828] = 29'b0_111110001010_100_0_011111000101;
      patterns[31829] = 29'b0_111110001010_101_1_001111100010;
      patterns[31830] = 29'b0_111110001010_110_0_111110001010;
      patterns[31831] = 29'b0_111110001010_111_0_111110001010;
      patterns[31832] = 29'b0_111110001011_000_0_111110001011;
      patterns[31833] = 29'b0_111110001011_001_0_001011111110;
      patterns[31834] = 29'b0_111110001011_010_1_111100010110;
      patterns[31835] = 29'b0_111110001011_011_1_111000101101;
      patterns[31836] = 29'b0_111110001011_100_1_011111000101;
      patterns[31837] = 29'b0_111110001011_101_1_101111100010;
      patterns[31838] = 29'b0_111110001011_110_0_111110001011;
      patterns[31839] = 29'b0_111110001011_111_0_111110001011;
      patterns[31840] = 29'b0_111110001100_000_0_111110001100;
      patterns[31841] = 29'b0_111110001100_001_0_001100111110;
      patterns[31842] = 29'b0_111110001100_010_1_111100011000;
      patterns[31843] = 29'b0_111110001100_011_1_111000110001;
      patterns[31844] = 29'b0_111110001100_100_0_011111000110;
      patterns[31845] = 29'b0_111110001100_101_0_001111100011;
      patterns[31846] = 29'b0_111110001100_110_0_111110001100;
      patterns[31847] = 29'b0_111110001100_111_0_111110001100;
      patterns[31848] = 29'b0_111110001101_000_0_111110001101;
      patterns[31849] = 29'b0_111110001101_001_0_001101111110;
      patterns[31850] = 29'b0_111110001101_010_1_111100011010;
      patterns[31851] = 29'b0_111110001101_011_1_111000110101;
      patterns[31852] = 29'b0_111110001101_100_1_011111000110;
      patterns[31853] = 29'b0_111110001101_101_0_101111100011;
      patterns[31854] = 29'b0_111110001101_110_0_111110001101;
      patterns[31855] = 29'b0_111110001101_111_0_111110001101;
      patterns[31856] = 29'b0_111110001110_000_0_111110001110;
      patterns[31857] = 29'b0_111110001110_001_0_001110111110;
      patterns[31858] = 29'b0_111110001110_010_1_111100011100;
      patterns[31859] = 29'b0_111110001110_011_1_111000111001;
      patterns[31860] = 29'b0_111110001110_100_0_011111000111;
      patterns[31861] = 29'b0_111110001110_101_1_001111100011;
      patterns[31862] = 29'b0_111110001110_110_0_111110001110;
      patterns[31863] = 29'b0_111110001110_111_0_111110001110;
      patterns[31864] = 29'b0_111110001111_000_0_111110001111;
      patterns[31865] = 29'b0_111110001111_001_0_001111111110;
      patterns[31866] = 29'b0_111110001111_010_1_111100011110;
      patterns[31867] = 29'b0_111110001111_011_1_111000111101;
      patterns[31868] = 29'b0_111110001111_100_1_011111000111;
      patterns[31869] = 29'b0_111110001111_101_1_101111100011;
      patterns[31870] = 29'b0_111110001111_110_0_111110001111;
      patterns[31871] = 29'b0_111110001111_111_0_111110001111;
      patterns[31872] = 29'b0_111110010000_000_0_111110010000;
      patterns[31873] = 29'b0_111110010000_001_0_010000111110;
      patterns[31874] = 29'b0_111110010000_010_1_111100100000;
      patterns[31875] = 29'b0_111110010000_011_1_111001000001;
      patterns[31876] = 29'b0_111110010000_100_0_011111001000;
      patterns[31877] = 29'b0_111110010000_101_0_001111100100;
      patterns[31878] = 29'b0_111110010000_110_0_111110010000;
      patterns[31879] = 29'b0_111110010000_111_0_111110010000;
      patterns[31880] = 29'b0_111110010001_000_0_111110010001;
      patterns[31881] = 29'b0_111110010001_001_0_010001111110;
      patterns[31882] = 29'b0_111110010001_010_1_111100100010;
      patterns[31883] = 29'b0_111110010001_011_1_111001000101;
      patterns[31884] = 29'b0_111110010001_100_1_011111001000;
      patterns[31885] = 29'b0_111110010001_101_0_101111100100;
      patterns[31886] = 29'b0_111110010001_110_0_111110010001;
      patterns[31887] = 29'b0_111110010001_111_0_111110010001;
      patterns[31888] = 29'b0_111110010010_000_0_111110010010;
      patterns[31889] = 29'b0_111110010010_001_0_010010111110;
      patterns[31890] = 29'b0_111110010010_010_1_111100100100;
      patterns[31891] = 29'b0_111110010010_011_1_111001001001;
      patterns[31892] = 29'b0_111110010010_100_0_011111001001;
      patterns[31893] = 29'b0_111110010010_101_1_001111100100;
      patterns[31894] = 29'b0_111110010010_110_0_111110010010;
      patterns[31895] = 29'b0_111110010010_111_0_111110010010;
      patterns[31896] = 29'b0_111110010011_000_0_111110010011;
      patterns[31897] = 29'b0_111110010011_001_0_010011111110;
      patterns[31898] = 29'b0_111110010011_010_1_111100100110;
      patterns[31899] = 29'b0_111110010011_011_1_111001001101;
      patterns[31900] = 29'b0_111110010011_100_1_011111001001;
      patterns[31901] = 29'b0_111110010011_101_1_101111100100;
      patterns[31902] = 29'b0_111110010011_110_0_111110010011;
      patterns[31903] = 29'b0_111110010011_111_0_111110010011;
      patterns[31904] = 29'b0_111110010100_000_0_111110010100;
      patterns[31905] = 29'b0_111110010100_001_0_010100111110;
      patterns[31906] = 29'b0_111110010100_010_1_111100101000;
      patterns[31907] = 29'b0_111110010100_011_1_111001010001;
      patterns[31908] = 29'b0_111110010100_100_0_011111001010;
      patterns[31909] = 29'b0_111110010100_101_0_001111100101;
      patterns[31910] = 29'b0_111110010100_110_0_111110010100;
      patterns[31911] = 29'b0_111110010100_111_0_111110010100;
      patterns[31912] = 29'b0_111110010101_000_0_111110010101;
      patterns[31913] = 29'b0_111110010101_001_0_010101111110;
      patterns[31914] = 29'b0_111110010101_010_1_111100101010;
      patterns[31915] = 29'b0_111110010101_011_1_111001010101;
      patterns[31916] = 29'b0_111110010101_100_1_011111001010;
      patterns[31917] = 29'b0_111110010101_101_0_101111100101;
      patterns[31918] = 29'b0_111110010101_110_0_111110010101;
      patterns[31919] = 29'b0_111110010101_111_0_111110010101;
      patterns[31920] = 29'b0_111110010110_000_0_111110010110;
      patterns[31921] = 29'b0_111110010110_001_0_010110111110;
      patterns[31922] = 29'b0_111110010110_010_1_111100101100;
      patterns[31923] = 29'b0_111110010110_011_1_111001011001;
      patterns[31924] = 29'b0_111110010110_100_0_011111001011;
      patterns[31925] = 29'b0_111110010110_101_1_001111100101;
      patterns[31926] = 29'b0_111110010110_110_0_111110010110;
      patterns[31927] = 29'b0_111110010110_111_0_111110010110;
      patterns[31928] = 29'b0_111110010111_000_0_111110010111;
      patterns[31929] = 29'b0_111110010111_001_0_010111111110;
      patterns[31930] = 29'b0_111110010111_010_1_111100101110;
      patterns[31931] = 29'b0_111110010111_011_1_111001011101;
      patterns[31932] = 29'b0_111110010111_100_1_011111001011;
      patterns[31933] = 29'b0_111110010111_101_1_101111100101;
      patterns[31934] = 29'b0_111110010111_110_0_111110010111;
      patterns[31935] = 29'b0_111110010111_111_0_111110010111;
      patterns[31936] = 29'b0_111110011000_000_0_111110011000;
      patterns[31937] = 29'b0_111110011000_001_0_011000111110;
      patterns[31938] = 29'b0_111110011000_010_1_111100110000;
      patterns[31939] = 29'b0_111110011000_011_1_111001100001;
      patterns[31940] = 29'b0_111110011000_100_0_011111001100;
      patterns[31941] = 29'b0_111110011000_101_0_001111100110;
      patterns[31942] = 29'b0_111110011000_110_0_111110011000;
      patterns[31943] = 29'b0_111110011000_111_0_111110011000;
      patterns[31944] = 29'b0_111110011001_000_0_111110011001;
      patterns[31945] = 29'b0_111110011001_001_0_011001111110;
      patterns[31946] = 29'b0_111110011001_010_1_111100110010;
      patterns[31947] = 29'b0_111110011001_011_1_111001100101;
      patterns[31948] = 29'b0_111110011001_100_1_011111001100;
      patterns[31949] = 29'b0_111110011001_101_0_101111100110;
      patterns[31950] = 29'b0_111110011001_110_0_111110011001;
      patterns[31951] = 29'b0_111110011001_111_0_111110011001;
      patterns[31952] = 29'b0_111110011010_000_0_111110011010;
      patterns[31953] = 29'b0_111110011010_001_0_011010111110;
      patterns[31954] = 29'b0_111110011010_010_1_111100110100;
      patterns[31955] = 29'b0_111110011010_011_1_111001101001;
      patterns[31956] = 29'b0_111110011010_100_0_011111001101;
      patterns[31957] = 29'b0_111110011010_101_1_001111100110;
      patterns[31958] = 29'b0_111110011010_110_0_111110011010;
      patterns[31959] = 29'b0_111110011010_111_0_111110011010;
      patterns[31960] = 29'b0_111110011011_000_0_111110011011;
      patterns[31961] = 29'b0_111110011011_001_0_011011111110;
      patterns[31962] = 29'b0_111110011011_010_1_111100110110;
      patterns[31963] = 29'b0_111110011011_011_1_111001101101;
      patterns[31964] = 29'b0_111110011011_100_1_011111001101;
      patterns[31965] = 29'b0_111110011011_101_1_101111100110;
      patterns[31966] = 29'b0_111110011011_110_0_111110011011;
      patterns[31967] = 29'b0_111110011011_111_0_111110011011;
      patterns[31968] = 29'b0_111110011100_000_0_111110011100;
      patterns[31969] = 29'b0_111110011100_001_0_011100111110;
      patterns[31970] = 29'b0_111110011100_010_1_111100111000;
      patterns[31971] = 29'b0_111110011100_011_1_111001110001;
      patterns[31972] = 29'b0_111110011100_100_0_011111001110;
      patterns[31973] = 29'b0_111110011100_101_0_001111100111;
      patterns[31974] = 29'b0_111110011100_110_0_111110011100;
      patterns[31975] = 29'b0_111110011100_111_0_111110011100;
      patterns[31976] = 29'b0_111110011101_000_0_111110011101;
      patterns[31977] = 29'b0_111110011101_001_0_011101111110;
      patterns[31978] = 29'b0_111110011101_010_1_111100111010;
      patterns[31979] = 29'b0_111110011101_011_1_111001110101;
      patterns[31980] = 29'b0_111110011101_100_1_011111001110;
      patterns[31981] = 29'b0_111110011101_101_0_101111100111;
      patterns[31982] = 29'b0_111110011101_110_0_111110011101;
      patterns[31983] = 29'b0_111110011101_111_0_111110011101;
      patterns[31984] = 29'b0_111110011110_000_0_111110011110;
      patterns[31985] = 29'b0_111110011110_001_0_011110111110;
      patterns[31986] = 29'b0_111110011110_010_1_111100111100;
      patterns[31987] = 29'b0_111110011110_011_1_111001111001;
      patterns[31988] = 29'b0_111110011110_100_0_011111001111;
      patterns[31989] = 29'b0_111110011110_101_1_001111100111;
      patterns[31990] = 29'b0_111110011110_110_0_111110011110;
      patterns[31991] = 29'b0_111110011110_111_0_111110011110;
      patterns[31992] = 29'b0_111110011111_000_0_111110011111;
      patterns[31993] = 29'b0_111110011111_001_0_011111111110;
      patterns[31994] = 29'b0_111110011111_010_1_111100111110;
      patterns[31995] = 29'b0_111110011111_011_1_111001111101;
      patterns[31996] = 29'b0_111110011111_100_1_011111001111;
      patterns[31997] = 29'b0_111110011111_101_1_101111100111;
      patterns[31998] = 29'b0_111110011111_110_0_111110011111;
      patterns[31999] = 29'b0_111110011111_111_0_111110011111;
      patterns[32000] = 29'b0_111110100000_000_0_111110100000;
      patterns[32001] = 29'b0_111110100000_001_0_100000111110;
      patterns[32002] = 29'b0_111110100000_010_1_111101000000;
      patterns[32003] = 29'b0_111110100000_011_1_111010000001;
      patterns[32004] = 29'b0_111110100000_100_0_011111010000;
      patterns[32005] = 29'b0_111110100000_101_0_001111101000;
      patterns[32006] = 29'b0_111110100000_110_0_111110100000;
      patterns[32007] = 29'b0_111110100000_111_0_111110100000;
      patterns[32008] = 29'b0_111110100001_000_0_111110100001;
      patterns[32009] = 29'b0_111110100001_001_0_100001111110;
      patterns[32010] = 29'b0_111110100001_010_1_111101000010;
      patterns[32011] = 29'b0_111110100001_011_1_111010000101;
      patterns[32012] = 29'b0_111110100001_100_1_011111010000;
      patterns[32013] = 29'b0_111110100001_101_0_101111101000;
      patterns[32014] = 29'b0_111110100001_110_0_111110100001;
      patterns[32015] = 29'b0_111110100001_111_0_111110100001;
      patterns[32016] = 29'b0_111110100010_000_0_111110100010;
      patterns[32017] = 29'b0_111110100010_001_0_100010111110;
      patterns[32018] = 29'b0_111110100010_010_1_111101000100;
      patterns[32019] = 29'b0_111110100010_011_1_111010001001;
      patterns[32020] = 29'b0_111110100010_100_0_011111010001;
      patterns[32021] = 29'b0_111110100010_101_1_001111101000;
      patterns[32022] = 29'b0_111110100010_110_0_111110100010;
      patterns[32023] = 29'b0_111110100010_111_0_111110100010;
      patterns[32024] = 29'b0_111110100011_000_0_111110100011;
      patterns[32025] = 29'b0_111110100011_001_0_100011111110;
      patterns[32026] = 29'b0_111110100011_010_1_111101000110;
      patterns[32027] = 29'b0_111110100011_011_1_111010001101;
      patterns[32028] = 29'b0_111110100011_100_1_011111010001;
      patterns[32029] = 29'b0_111110100011_101_1_101111101000;
      patterns[32030] = 29'b0_111110100011_110_0_111110100011;
      patterns[32031] = 29'b0_111110100011_111_0_111110100011;
      patterns[32032] = 29'b0_111110100100_000_0_111110100100;
      patterns[32033] = 29'b0_111110100100_001_0_100100111110;
      patterns[32034] = 29'b0_111110100100_010_1_111101001000;
      patterns[32035] = 29'b0_111110100100_011_1_111010010001;
      patterns[32036] = 29'b0_111110100100_100_0_011111010010;
      patterns[32037] = 29'b0_111110100100_101_0_001111101001;
      patterns[32038] = 29'b0_111110100100_110_0_111110100100;
      patterns[32039] = 29'b0_111110100100_111_0_111110100100;
      patterns[32040] = 29'b0_111110100101_000_0_111110100101;
      patterns[32041] = 29'b0_111110100101_001_0_100101111110;
      patterns[32042] = 29'b0_111110100101_010_1_111101001010;
      patterns[32043] = 29'b0_111110100101_011_1_111010010101;
      patterns[32044] = 29'b0_111110100101_100_1_011111010010;
      patterns[32045] = 29'b0_111110100101_101_0_101111101001;
      patterns[32046] = 29'b0_111110100101_110_0_111110100101;
      patterns[32047] = 29'b0_111110100101_111_0_111110100101;
      patterns[32048] = 29'b0_111110100110_000_0_111110100110;
      patterns[32049] = 29'b0_111110100110_001_0_100110111110;
      patterns[32050] = 29'b0_111110100110_010_1_111101001100;
      patterns[32051] = 29'b0_111110100110_011_1_111010011001;
      patterns[32052] = 29'b0_111110100110_100_0_011111010011;
      patterns[32053] = 29'b0_111110100110_101_1_001111101001;
      patterns[32054] = 29'b0_111110100110_110_0_111110100110;
      patterns[32055] = 29'b0_111110100110_111_0_111110100110;
      patterns[32056] = 29'b0_111110100111_000_0_111110100111;
      patterns[32057] = 29'b0_111110100111_001_0_100111111110;
      patterns[32058] = 29'b0_111110100111_010_1_111101001110;
      patterns[32059] = 29'b0_111110100111_011_1_111010011101;
      patterns[32060] = 29'b0_111110100111_100_1_011111010011;
      patterns[32061] = 29'b0_111110100111_101_1_101111101001;
      patterns[32062] = 29'b0_111110100111_110_0_111110100111;
      patterns[32063] = 29'b0_111110100111_111_0_111110100111;
      patterns[32064] = 29'b0_111110101000_000_0_111110101000;
      patterns[32065] = 29'b0_111110101000_001_0_101000111110;
      patterns[32066] = 29'b0_111110101000_010_1_111101010000;
      patterns[32067] = 29'b0_111110101000_011_1_111010100001;
      patterns[32068] = 29'b0_111110101000_100_0_011111010100;
      patterns[32069] = 29'b0_111110101000_101_0_001111101010;
      patterns[32070] = 29'b0_111110101000_110_0_111110101000;
      patterns[32071] = 29'b0_111110101000_111_0_111110101000;
      patterns[32072] = 29'b0_111110101001_000_0_111110101001;
      patterns[32073] = 29'b0_111110101001_001_0_101001111110;
      patterns[32074] = 29'b0_111110101001_010_1_111101010010;
      patterns[32075] = 29'b0_111110101001_011_1_111010100101;
      patterns[32076] = 29'b0_111110101001_100_1_011111010100;
      patterns[32077] = 29'b0_111110101001_101_0_101111101010;
      patterns[32078] = 29'b0_111110101001_110_0_111110101001;
      patterns[32079] = 29'b0_111110101001_111_0_111110101001;
      patterns[32080] = 29'b0_111110101010_000_0_111110101010;
      patterns[32081] = 29'b0_111110101010_001_0_101010111110;
      patterns[32082] = 29'b0_111110101010_010_1_111101010100;
      patterns[32083] = 29'b0_111110101010_011_1_111010101001;
      patterns[32084] = 29'b0_111110101010_100_0_011111010101;
      patterns[32085] = 29'b0_111110101010_101_1_001111101010;
      patterns[32086] = 29'b0_111110101010_110_0_111110101010;
      patterns[32087] = 29'b0_111110101010_111_0_111110101010;
      patterns[32088] = 29'b0_111110101011_000_0_111110101011;
      patterns[32089] = 29'b0_111110101011_001_0_101011111110;
      patterns[32090] = 29'b0_111110101011_010_1_111101010110;
      patterns[32091] = 29'b0_111110101011_011_1_111010101101;
      patterns[32092] = 29'b0_111110101011_100_1_011111010101;
      patterns[32093] = 29'b0_111110101011_101_1_101111101010;
      patterns[32094] = 29'b0_111110101011_110_0_111110101011;
      patterns[32095] = 29'b0_111110101011_111_0_111110101011;
      patterns[32096] = 29'b0_111110101100_000_0_111110101100;
      patterns[32097] = 29'b0_111110101100_001_0_101100111110;
      patterns[32098] = 29'b0_111110101100_010_1_111101011000;
      patterns[32099] = 29'b0_111110101100_011_1_111010110001;
      patterns[32100] = 29'b0_111110101100_100_0_011111010110;
      patterns[32101] = 29'b0_111110101100_101_0_001111101011;
      patterns[32102] = 29'b0_111110101100_110_0_111110101100;
      patterns[32103] = 29'b0_111110101100_111_0_111110101100;
      patterns[32104] = 29'b0_111110101101_000_0_111110101101;
      patterns[32105] = 29'b0_111110101101_001_0_101101111110;
      patterns[32106] = 29'b0_111110101101_010_1_111101011010;
      patterns[32107] = 29'b0_111110101101_011_1_111010110101;
      patterns[32108] = 29'b0_111110101101_100_1_011111010110;
      patterns[32109] = 29'b0_111110101101_101_0_101111101011;
      patterns[32110] = 29'b0_111110101101_110_0_111110101101;
      patterns[32111] = 29'b0_111110101101_111_0_111110101101;
      patterns[32112] = 29'b0_111110101110_000_0_111110101110;
      patterns[32113] = 29'b0_111110101110_001_0_101110111110;
      patterns[32114] = 29'b0_111110101110_010_1_111101011100;
      patterns[32115] = 29'b0_111110101110_011_1_111010111001;
      patterns[32116] = 29'b0_111110101110_100_0_011111010111;
      patterns[32117] = 29'b0_111110101110_101_1_001111101011;
      patterns[32118] = 29'b0_111110101110_110_0_111110101110;
      patterns[32119] = 29'b0_111110101110_111_0_111110101110;
      patterns[32120] = 29'b0_111110101111_000_0_111110101111;
      patterns[32121] = 29'b0_111110101111_001_0_101111111110;
      patterns[32122] = 29'b0_111110101111_010_1_111101011110;
      patterns[32123] = 29'b0_111110101111_011_1_111010111101;
      patterns[32124] = 29'b0_111110101111_100_1_011111010111;
      patterns[32125] = 29'b0_111110101111_101_1_101111101011;
      patterns[32126] = 29'b0_111110101111_110_0_111110101111;
      patterns[32127] = 29'b0_111110101111_111_0_111110101111;
      patterns[32128] = 29'b0_111110110000_000_0_111110110000;
      patterns[32129] = 29'b0_111110110000_001_0_110000111110;
      patterns[32130] = 29'b0_111110110000_010_1_111101100000;
      patterns[32131] = 29'b0_111110110000_011_1_111011000001;
      patterns[32132] = 29'b0_111110110000_100_0_011111011000;
      patterns[32133] = 29'b0_111110110000_101_0_001111101100;
      patterns[32134] = 29'b0_111110110000_110_0_111110110000;
      patterns[32135] = 29'b0_111110110000_111_0_111110110000;
      patterns[32136] = 29'b0_111110110001_000_0_111110110001;
      patterns[32137] = 29'b0_111110110001_001_0_110001111110;
      patterns[32138] = 29'b0_111110110001_010_1_111101100010;
      patterns[32139] = 29'b0_111110110001_011_1_111011000101;
      patterns[32140] = 29'b0_111110110001_100_1_011111011000;
      patterns[32141] = 29'b0_111110110001_101_0_101111101100;
      patterns[32142] = 29'b0_111110110001_110_0_111110110001;
      patterns[32143] = 29'b0_111110110001_111_0_111110110001;
      patterns[32144] = 29'b0_111110110010_000_0_111110110010;
      patterns[32145] = 29'b0_111110110010_001_0_110010111110;
      patterns[32146] = 29'b0_111110110010_010_1_111101100100;
      patterns[32147] = 29'b0_111110110010_011_1_111011001001;
      patterns[32148] = 29'b0_111110110010_100_0_011111011001;
      patterns[32149] = 29'b0_111110110010_101_1_001111101100;
      patterns[32150] = 29'b0_111110110010_110_0_111110110010;
      patterns[32151] = 29'b0_111110110010_111_0_111110110010;
      patterns[32152] = 29'b0_111110110011_000_0_111110110011;
      patterns[32153] = 29'b0_111110110011_001_0_110011111110;
      patterns[32154] = 29'b0_111110110011_010_1_111101100110;
      patterns[32155] = 29'b0_111110110011_011_1_111011001101;
      patterns[32156] = 29'b0_111110110011_100_1_011111011001;
      patterns[32157] = 29'b0_111110110011_101_1_101111101100;
      patterns[32158] = 29'b0_111110110011_110_0_111110110011;
      patterns[32159] = 29'b0_111110110011_111_0_111110110011;
      patterns[32160] = 29'b0_111110110100_000_0_111110110100;
      patterns[32161] = 29'b0_111110110100_001_0_110100111110;
      patterns[32162] = 29'b0_111110110100_010_1_111101101000;
      patterns[32163] = 29'b0_111110110100_011_1_111011010001;
      patterns[32164] = 29'b0_111110110100_100_0_011111011010;
      patterns[32165] = 29'b0_111110110100_101_0_001111101101;
      patterns[32166] = 29'b0_111110110100_110_0_111110110100;
      patterns[32167] = 29'b0_111110110100_111_0_111110110100;
      patterns[32168] = 29'b0_111110110101_000_0_111110110101;
      patterns[32169] = 29'b0_111110110101_001_0_110101111110;
      patterns[32170] = 29'b0_111110110101_010_1_111101101010;
      patterns[32171] = 29'b0_111110110101_011_1_111011010101;
      patterns[32172] = 29'b0_111110110101_100_1_011111011010;
      patterns[32173] = 29'b0_111110110101_101_0_101111101101;
      patterns[32174] = 29'b0_111110110101_110_0_111110110101;
      patterns[32175] = 29'b0_111110110101_111_0_111110110101;
      patterns[32176] = 29'b0_111110110110_000_0_111110110110;
      patterns[32177] = 29'b0_111110110110_001_0_110110111110;
      patterns[32178] = 29'b0_111110110110_010_1_111101101100;
      patterns[32179] = 29'b0_111110110110_011_1_111011011001;
      patterns[32180] = 29'b0_111110110110_100_0_011111011011;
      patterns[32181] = 29'b0_111110110110_101_1_001111101101;
      patterns[32182] = 29'b0_111110110110_110_0_111110110110;
      patterns[32183] = 29'b0_111110110110_111_0_111110110110;
      patterns[32184] = 29'b0_111110110111_000_0_111110110111;
      patterns[32185] = 29'b0_111110110111_001_0_110111111110;
      patterns[32186] = 29'b0_111110110111_010_1_111101101110;
      patterns[32187] = 29'b0_111110110111_011_1_111011011101;
      patterns[32188] = 29'b0_111110110111_100_1_011111011011;
      patterns[32189] = 29'b0_111110110111_101_1_101111101101;
      patterns[32190] = 29'b0_111110110111_110_0_111110110111;
      patterns[32191] = 29'b0_111110110111_111_0_111110110111;
      patterns[32192] = 29'b0_111110111000_000_0_111110111000;
      patterns[32193] = 29'b0_111110111000_001_0_111000111110;
      patterns[32194] = 29'b0_111110111000_010_1_111101110000;
      patterns[32195] = 29'b0_111110111000_011_1_111011100001;
      patterns[32196] = 29'b0_111110111000_100_0_011111011100;
      patterns[32197] = 29'b0_111110111000_101_0_001111101110;
      patterns[32198] = 29'b0_111110111000_110_0_111110111000;
      patterns[32199] = 29'b0_111110111000_111_0_111110111000;
      patterns[32200] = 29'b0_111110111001_000_0_111110111001;
      patterns[32201] = 29'b0_111110111001_001_0_111001111110;
      patterns[32202] = 29'b0_111110111001_010_1_111101110010;
      patterns[32203] = 29'b0_111110111001_011_1_111011100101;
      patterns[32204] = 29'b0_111110111001_100_1_011111011100;
      patterns[32205] = 29'b0_111110111001_101_0_101111101110;
      patterns[32206] = 29'b0_111110111001_110_0_111110111001;
      patterns[32207] = 29'b0_111110111001_111_0_111110111001;
      patterns[32208] = 29'b0_111110111010_000_0_111110111010;
      patterns[32209] = 29'b0_111110111010_001_0_111010111110;
      patterns[32210] = 29'b0_111110111010_010_1_111101110100;
      patterns[32211] = 29'b0_111110111010_011_1_111011101001;
      patterns[32212] = 29'b0_111110111010_100_0_011111011101;
      patterns[32213] = 29'b0_111110111010_101_1_001111101110;
      patterns[32214] = 29'b0_111110111010_110_0_111110111010;
      patterns[32215] = 29'b0_111110111010_111_0_111110111010;
      patterns[32216] = 29'b0_111110111011_000_0_111110111011;
      patterns[32217] = 29'b0_111110111011_001_0_111011111110;
      patterns[32218] = 29'b0_111110111011_010_1_111101110110;
      patterns[32219] = 29'b0_111110111011_011_1_111011101101;
      patterns[32220] = 29'b0_111110111011_100_1_011111011101;
      patterns[32221] = 29'b0_111110111011_101_1_101111101110;
      patterns[32222] = 29'b0_111110111011_110_0_111110111011;
      patterns[32223] = 29'b0_111110111011_111_0_111110111011;
      patterns[32224] = 29'b0_111110111100_000_0_111110111100;
      patterns[32225] = 29'b0_111110111100_001_0_111100111110;
      patterns[32226] = 29'b0_111110111100_010_1_111101111000;
      patterns[32227] = 29'b0_111110111100_011_1_111011110001;
      patterns[32228] = 29'b0_111110111100_100_0_011111011110;
      patterns[32229] = 29'b0_111110111100_101_0_001111101111;
      patterns[32230] = 29'b0_111110111100_110_0_111110111100;
      patterns[32231] = 29'b0_111110111100_111_0_111110111100;
      patterns[32232] = 29'b0_111110111101_000_0_111110111101;
      patterns[32233] = 29'b0_111110111101_001_0_111101111110;
      patterns[32234] = 29'b0_111110111101_010_1_111101111010;
      patterns[32235] = 29'b0_111110111101_011_1_111011110101;
      patterns[32236] = 29'b0_111110111101_100_1_011111011110;
      patterns[32237] = 29'b0_111110111101_101_0_101111101111;
      patterns[32238] = 29'b0_111110111101_110_0_111110111101;
      patterns[32239] = 29'b0_111110111101_111_0_111110111101;
      patterns[32240] = 29'b0_111110111110_000_0_111110111110;
      patterns[32241] = 29'b0_111110111110_001_0_111110111110;
      patterns[32242] = 29'b0_111110111110_010_1_111101111100;
      patterns[32243] = 29'b0_111110111110_011_1_111011111001;
      patterns[32244] = 29'b0_111110111110_100_0_011111011111;
      patterns[32245] = 29'b0_111110111110_101_1_001111101111;
      patterns[32246] = 29'b0_111110111110_110_0_111110111110;
      patterns[32247] = 29'b0_111110111110_111_0_111110111110;
      patterns[32248] = 29'b0_111110111111_000_0_111110111111;
      patterns[32249] = 29'b0_111110111111_001_0_111111111110;
      patterns[32250] = 29'b0_111110111111_010_1_111101111110;
      patterns[32251] = 29'b0_111110111111_011_1_111011111101;
      patterns[32252] = 29'b0_111110111111_100_1_011111011111;
      patterns[32253] = 29'b0_111110111111_101_1_101111101111;
      patterns[32254] = 29'b0_111110111111_110_0_111110111111;
      patterns[32255] = 29'b0_111110111111_111_0_111110111111;
      patterns[32256] = 29'b0_111111000000_000_0_111111000000;
      patterns[32257] = 29'b0_111111000000_001_0_000000111111;
      patterns[32258] = 29'b0_111111000000_010_1_111110000000;
      patterns[32259] = 29'b0_111111000000_011_1_111100000001;
      patterns[32260] = 29'b0_111111000000_100_0_011111100000;
      patterns[32261] = 29'b0_111111000000_101_0_001111110000;
      patterns[32262] = 29'b0_111111000000_110_0_111111000000;
      patterns[32263] = 29'b0_111111000000_111_0_111111000000;
      patterns[32264] = 29'b0_111111000001_000_0_111111000001;
      patterns[32265] = 29'b0_111111000001_001_0_000001111111;
      patterns[32266] = 29'b0_111111000001_010_1_111110000010;
      patterns[32267] = 29'b0_111111000001_011_1_111100000101;
      patterns[32268] = 29'b0_111111000001_100_1_011111100000;
      patterns[32269] = 29'b0_111111000001_101_0_101111110000;
      patterns[32270] = 29'b0_111111000001_110_0_111111000001;
      patterns[32271] = 29'b0_111111000001_111_0_111111000001;
      patterns[32272] = 29'b0_111111000010_000_0_111111000010;
      patterns[32273] = 29'b0_111111000010_001_0_000010111111;
      patterns[32274] = 29'b0_111111000010_010_1_111110000100;
      patterns[32275] = 29'b0_111111000010_011_1_111100001001;
      patterns[32276] = 29'b0_111111000010_100_0_011111100001;
      patterns[32277] = 29'b0_111111000010_101_1_001111110000;
      patterns[32278] = 29'b0_111111000010_110_0_111111000010;
      patterns[32279] = 29'b0_111111000010_111_0_111111000010;
      patterns[32280] = 29'b0_111111000011_000_0_111111000011;
      patterns[32281] = 29'b0_111111000011_001_0_000011111111;
      patterns[32282] = 29'b0_111111000011_010_1_111110000110;
      patterns[32283] = 29'b0_111111000011_011_1_111100001101;
      patterns[32284] = 29'b0_111111000011_100_1_011111100001;
      patterns[32285] = 29'b0_111111000011_101_1_101111110000;
      patterns[32286] = 29'b0_111111000011_110_0_111111000011;
      patterns[32287] = 29'b0_111111000011_111_0_111111000011;
      patterns[32288] = 29'b0_111111000100_000_0_111111000100;
      patterns[32289] = 29'b0_111111000100_001_0_000100111111;
      patterns[32290] = 29'b0_111111000100_010_1_111110001000;
      patterns[32291] = 29'b0_111111000100_011_1_111100010001;
      patterns[32292] = 29'b0_111111000100_100_0_011111100010;
      patterns[32293] = 29'b0_111111000100_101_0_001111110001;
      patterns[32294] = 29'b0_111111000100_110_0_111111000100;
      patterns[32295] = 29'b0_111111000100_111_0_111111000100;
      patterns[32296] = 29'b0_111111000101_000_0_111111000101;
      patterns[32297] = 29'b0_111111000101_001_0_000101111111;
      patterns[32298] = 29'b0_111111000101_010_1_111110001010;
      patterns[32299] = 29'b0_111111000101_011_1_111100010101;
      patterns[32300] = 29'b0_111111000101_100_1_011111100010;
      patterns[32301] = 29'b0_111111000101_101_0_101111110001;
      patterns[32302] = 29'b0_111111000101_110_0_111111000101;
      patterns[32303] = 29'b0_111111000101_111_0_111111000101;
      patterns[32304] = 29'b0_111111000110_000_0_111111000110;
      patterns[32305] = 29'b0_111111000110_001_0_000110111111;
      patterns[32306] = 29'b0_111111000110_010_1_111110001100;
      patterns[32307] = 29'b0_111111000110_011_1_111100011001;
      patterns[32308] = 29'b0_111111000110_100_0_011111100011;
      patterns[32309] = 29'b0_111111000110_101_1_001111110001;
      patterns[32310] = 29'b0_111111000110_110_0_111111000110;
      patterns[32311] = 29'b0_111111000110_111_0_111111000110;
      patterns[32312] = 29'b0_111111000111_000_0_111111000111;
      patterns[32313] = 29'b0_111111000111_001_0_000111111111;
      patterns[32314] = 29'b0_111111000111_010_1_111110001110;
      patterns[32315] = 29'b0_111111000111_011_1_111100011101;
      patterns[32316] = 29'b0_111111000111_100_1_011111100011;
      patterns[32317] = 29'b0_111111000111_101_1_101111110001;
      patterns[32318] = 29'b0_111111000111_110_0_111111000111;
      patterns[32319] = 29'b0_111111000111_111_0_111111000111;
      patterns[32320] = 29'b0_111111001000_000_0_111111001000;
      patterns[32321] = 29'b0_111111001000_001_0_001000111111;
      patterns[32322] = 29'b0_111111001000_010_1_111110010000;
      patterns[32323] = 29'b0_111111001000_011_1_111100100001;
      patterns[32324] = 29'b0_111111001000_100_0_011111100100;
      patterns[32325] = 29'b0_111111001000_101_0_001111110010;
      patterns[32326] = 29'b0_111111001000_110_0_111111001000;
      patterns[32327] = 29'b0_111111001000_111_0_111111001000;
      patterns[32328] = 29'b0_111111001001_000_0_111111001001;
      patterns[32329] = 29'b0_111111001001_001_0_001001111111;
      patterns[32330] = 29'b0_111111001001_010_1_111110010010;
      patterns[32331] = 29'b0_111111001001_011_1_111100100101;
      patterns[32332] = 29'b0_111111001001_100_1_011111100100;
      patterns[32333] = 29'b0_111111001001_101_0_101111110010;
      patterns[32334] = 29'b0_111111001001_110_0_111111001001;
      patterns[32335] = 29'b0_111111001001_111_0_111111001001;
      patterns[32336] = 29'b0_111111001010_000_0_111111001010;
      patterns[32337] = 29'b0_111111001010_001_0_001010111111;
      patterns[32338] = 29'b0_111111001010_010_1_111110010100;
      patterns[32339] = 29'b0_111111001010_011_1_111100101001;
      patterns[32340] = 29'b0_111111001010_100_0_011111100101;
      patterns[32341] = 29'b0_111111001010_101_1_001111110010;
      patterns[32342] = 29'b0_111111001010_110_0_111111001010;
      patterns[32343] = 29'b0_111111001010_111_0_111111001010;
      patterns[32344] = 29'b0_111111001011_000_0_111111001011;
      patterns[32345] = 29'b0_111111001011_001_0_001011111111;
      patterns[32346] = 29'b0_111111001011_010_1_111110010110;
      patterns[32347] = 29'b0_111111001011_011_1_111100101101;
      patterns[32348] = 29'b0_111111001011_100_1_011111100101;
      patterns[32349] = 29'b0_111111001011_101_1_101111110010;
      patterns[32350] = 29'b0_111111001011_110_0_111111001011;
      patterns[32351] = 29'b0_111111001011_111_0_111111001011;
      patterns[32352] = 29'b0_111111001100_000_0_111111001100;
      patterns[32353] = 29'b0_111111001100_001_0_001100111111;
      patterns[32354] = 29'b0_111111001100_010_1_111110011000;
      patterns[32355] = 29'b0_111111001100_011_1_111100110001;
      patterns[32356] = 29'b0_111111001100_100_0_011111100110;
      patterns[32357] = 29'b0_111111001100_101_0_001111110011;
      patterns[32358] = 29'b0_111111001100_110_0_111111001100;
      patterns[32359] = 29'b0_111111001100_111_0_111111001100;
      patterns[32360] = 29'b0_111111001101_000_0_111111001101;
      patterns[32361] = 29'b0_111111001101_001_0_001101111111;
      patterns[32362] = 29'b0_111111001101_010_1_111110011010;
      patterns[32363] = 29'b0_111111001101_011_1_111100110101;
      patterns[32364] = 29'b0_111111001101_100_1_011111100110;
      patterns[32365] = 29'b0_111111001101_101_0_101111110011;
      patterns[32366] = 29'b0_111111001101_110_0_111111001101;
      patterns[32367] = 29'b0_111111001101_111_0_111111001101;
      patterns[32368] = 29'b0_111111001110_000_0_111111001110;
      patterns[32369] = 29'b0_111111001110_001_0_001110111111;
      patterns[32370] = 29'b0_111111001110_010_1_111110011100;
      patterns[32371] = 29'b0_111111001110_011_1_111100111001;
      patterns[32372] = 29'b0_111111001110_100_0_011111100111;
      patterns[32373] = 29'b0_111111001110_101_1_001111110011;
      patterns[32374] = 29'b0_111111001110_110_0_111111001110;
      patterns[32375] = 29'b0_111111001110_111_0_111111001110;
      patterns[32376] = 29'b0_111111001111_000_0_111111001111;
      patterns[32377] = 29'b0_111111001111_001_0_001111111111;
      patterns[32378] = 29'b0_111111001111_010_1_111110011110;
      patterns[32379] = 29'b0_111111001111_011_1_111100111101;
      patterns[32380] = 29'b0_111111001111_100_1_011111100111;
      patterns[32381] = 29'b0_111111001111_101_1_101111110011;
      patterns[32382] = 29'b0_111111001111_110_0_111111001111;
      patterns[32383] = 29'b0_111111001111_111_0_111111001111;
      patterns[32384] = 29'b0_111111010000_000_0_111111010000;
      patterns[32385] = 29'b0_111111010000_001_0_010000111111;
      patterns[32386] = 29'b0_111111010000_010_1_111110100000;
      patterns[32387] = 29'b0_111111010000_011_1_111101000001;
      patterns[32388] = 29'b0_111111010000_100_0_011111101000;
      patterns[32389] = 29'b0_111111010000_101_0_001111110100;
      patterns[32390] = 29'b0_111111010000_110_0_111111010000;
      patterns[32391] = 29'b0_111111010000_111_0_111111010000;
      patterns[32392] = 29'b0_111111010001_000_0_111111010001;
      patterns[32393] = 29'b0_111111010001_001_0_010001111111;
      patterns[32394] = 29'b0_111111010001_010_1_111110100010;
      patterns[32395] = 29'b0_111111010001_011_1_111101000101;
      patterns[32396] = 29'b0_111111010001_100_1_011111101000;
      patterns[32397] = 29'b0_111111010001_101_0_101111110100;
      patterns[32398] = 29'b0_111111010001_110_0_111111010001;
      patterns[32399] = 29'b0_111111010001_111_0_111111010001;
      patterns[32400] = 29'b0_111111010010_000_0_111111010010;
      patterns[32401] = 29'b0_111111010010_001_0_010010111111;
      patterns[32402] = 29'b0_111111010010_010_1_111110100100;
      patterns[32403] = 29'b0_111111010010_011_1_111101001001;
      patterns[32404] = 29'b0_111111010010_100_0_011111101001;
      patterns[32405] = 29'b0_111111010010_101_1_001111110100;
      patterns[32406] = 29'b0_111111010010_110_0_111111010010;
      patterns[32407] = 29'b0_111111010010_111_0_111111010010;
      patterns[32408] = 29'b0_111111010011_000_0_111111010011;
      patterns[32409] = 29'b0_111111010011_001_0_010011111111;
      patterns[32410] = 29'b0_111111010011_010_1_111110100110;
      patterns[32411] = 29'b0_111111010011_011_1_111101001101;
      patterns[32412] = 29'b0_111111010011_100_1_011111101001;
      patterns[32413] = 29'b0_111111010011_101_1_101111110100;
      patterns[32414] = 29'b0_111111010011_110_0_111111010011;
      patterns[32415] = 29'b0_111111010011_111_0_111111010011;
      patterns[32416] = 29'b0_111111010100_000_0_111111010100;
      patterns[32417] = 29'b0_111111010100_001_0_010100111111;
      patterns[32418] = 29'b0_111111010100_010_1_111110101000;
      patterns[32419] = 29'b0_111111010100_011_1_111101010001;
      patterns[32420] = 29'b0_111111010100_100_0_011111101010;
      patterns[32421] = 29'b0_111111010100_101_0_001111110101;
      patterns[32422] = 29'b0_111111010100_110_0_111111010100;
      patterns[32423] = 29'b0_111111010100_111_0_111111010100;
      patterns[32424] = 29'b0_111111010101_000_0_111111010101;
      patterns[32425] = 29'b0_111111010101_001_0_010101111111;
      patterns[32426] = 29'b0_111111010101_010_1_111110101010;
      patterns[32427] = 29'b0_111111010101_011_1_111101010101;
      patterns[32428] = 29'b0_111111010101_100_1_011111101010;
      patterns[32429] = 29'b0_111111010101_101_0_101111110101;
      patterns[32430] = 29'b0_111111010101_110_0_111111010101;
      patterns[32431] = 29'b0_111111010101_111_0_111111010101;
      patterns[32432] = 29'b0_111111010110_000_0_111111010110;
      patterns[32433] = 29'b0_111111010110_001_0_010110111111;
      patterns[32434] = 29'b0_111111010110_010_1_111110101100;
      patterns[32435] = 29'b0_111111010110_011_1_111101011001;
      patterns[32436] = 29'b0_111111010110_100_0_011111101011;
      patterns[32437] = 29'b0_111111010110_101_1_001111110101;
      patterns[32438] = 29'b0_111111010110_110_0_111111010110;
      patterns[32439] = 29'b0_111111010110_111_0_111111010110;
      patterns[32440] = 29'b0_111111010111_000_0_111111010111;
      patterns[32441] = 29'b0_111111010111_001_0_010111111111;
      patterns[32442] = 29'b0_111111010111_010_1_111110101110;
      patterns[32443] = 29'b0_111111010111_011_1_111101011101;
      patterns[32444] = 29'b0_111111010111_100_1_011111101011;
      patterns[32445] = 29'b0_111111010111_101_1_101111110101;
      patterns[32446] = 29'b0_111111010111_110_0_111111010111;
      patterns[32447] = 29'b0_111111010111_111_0_111111010111;
      patterns[32448] = 29'b0_111111011000_000_0_111111011000;
      patterns[32449] = 29'b0_111111011000_001_0_011000111111;
      patterns[32450] = 29'b0_111111011000_010_1_111110110000;
      patterns[32451] = 29'b0_111111011000_011_1_111101100001;
      patterns[32452] = 29'b0_111111011000_100_0_011111101100;
      patterns[32453] = 29'b0_111111011000_101_0_001111110110;
      patterns[32454] = 29'b0_111111011000_110_0_111111011000;
      patterns[32455] = 29'b0_111111011000_111_0_111111011000;
      patterns[32456] = 29'b0_111111011001_000_0_111111011001;
      patterns[32457] = 29'b0_111111011001_001_0_011001111111;
      patterns[32458] = 29'b0_111111011001_010_1_111110110010;
      patterns[32459] = 29'b0_111111011001_011_1_111101100101;
      patterns[32460] = 29'b0_111111011001_100_1_011111101100;
      patterns[32461] = 29'b0_111111011001_101_0_101111110110;
      patterns[32462] = 29'b0_111111011001_110_0_111111011001;
      patterns[32463] = 29'b0_111111011001_111_0_111111011001;
      patterns[32464] = 29'b0_111111011010_000_0_111111011010;
      patterns[32465] = 29'b0_111111011010_001_0_011010111111;
      patterns[32466] = 29'b0_111111011010_010_1_111110110100;
      patterns[32467] = 29'b0_111111011010_011_1_111101101001;
      patterns[32468] = 29'b0_111111011010_100_0_011111101101;
      patterns[32469] = 29'b0_111111011010_101_1_001111110110;
      patterns[32470] = 29'b0_111111011010_110_0_111111011010;
      patterns[32471] = 29'b0_111111011010_111_0_111111011010;
      patterns[32472] = 29'b0_111111011011_000_0_111111011011;
      patterns[32473] = 29'b0_111111011011_001_0_011011111111;
      patterns[32474] = 29'b0_111111011011_010_1_111110110110;
      patterns[32475] = 29'b0_111111011011_011_1_111101101101;
      patterns[32476] = 29'b0_111111011011_100_1_011111101101;
      patterns[32477] = 29'b0_111111011011_101_1_101111110110;
      patterns[32478] = 29'b0_111111011011_110_0_111111011011;
      patterns[32479] = 29'b0_111111011011_111_0_111111011011;
      patterns[32480] = 29'b0_111111011100_000_0_111111011100;
      patterns[32481] = 29'b0_111111011100_001_0_011100111111;
      patterns[32482] = 29'b0_111111011100_010_1_111110111000;
      patterns[32483] = 29'b0_111111011100_011_1_111101110001;
      patterns[32484] = 29'b0_111111011100_100_0_011111101110;
      patterns[32485] = 29'b0_111111011100_101_0_001111110111;
      patterns[32486] = 29'b0_111111011100_110_0_111111011100;
      patterns[32487] = 29'b0_111111011100_111_0_111111011100;
      patterns[32488] = 29'b0_111111011101_000_0_111111011101;
      patterns[32489] = 29'b0_111111011101_001_0_011101111111;
      patterns[32490] = 29'b0_111111011101_010_1_111110111010;
      patterns[32491] = 29'b0_111111011101_011_1_111101110101;
      patterns[32492] = 29'b0_111111011101_100_1_011111101110;
      patterns[32493] = 29'b0_111111011101_101_0_101111110111;
      patterns[32494] = 29'b0_111111011101_110_0_111111011101;
      patterns[32495] = 29'b0_111111011101_111_0_111111011101;
      patterns[32496] = 29'b0_111111011110_000_0_111111011110;
      patterns[32497] = 29'b0_111111011110_001_0_011110111111;
      patterns[32498] = 29'b0_111111011110_010_1_111110111100;
      patterns[32499] = 29'b0_111111011110_011_1_111101111001;
      patterns[32500] = 29'b0_111111011110_100_0_011111101111;
      patterns[32501] = 29'b0_111111011110_101_1_001111110111;
      patterns[32502] = 29'b0_111111011110_110_0_111111011110;
      patterns[32503] = 29'b0_111111011110_111_0_111111011110;
      patterns[32504] = 29'b0_111111011111_000_0_111111011111;
      patterns[32505] = 29'b0_111111011111_001_0_011111111111;
      patterns[32506] = 29'b0_111111011111_010_1_111110111110;
      patterns[32507] = 29'b0_111111011111_011_1_111101111101;
      patterns[32508] = 29'b0_111111011111_100_1_011111101111;
      patterns[32509] = 29'b0_111111011111_101_1_101111110111;
      patterns[32510] = 29'b0_111111011111_110_0_111111011111;
      patterns[32511] = 29'b0_111111011111_111_0_111111011111;
      patterns[32512] = 29'b0_111111100000_000_0_111111100000;
      patterns[32513] = 29'b0_111111100000_001_0_100000111111;
      patterns[32514] = 29'b0_111111100000_010_1_111111000000;
      patterns[32515] = 29'b0_111111100000_011_1_111110000001;
      patterns[32516] = 29'b0_111111100000_100_0_011111110000;
      patterns[32517] = 29'b0_111111100000_101_0_001111111000;
      patterns[32518] = 29'b0_111111100000_110_0_111111100000;
      patterns[32519] = 29'b0_111111100000_111_0_111111100000;
      patterns[32520] = 29'b0_111111100001_000_0_111111100001;
      patterns[32521] = 29'b0_111111100001_001_0_100001111111;
      patterns[32522] = 29'b0_111111100001_010_1_111111000010;
      patterns[32523] = 29'b0_111111100001_011_1_111110000101;
      patterns[32524] = 29'b0_111111100001_100_1_011111110000;
      patterns[32525] = 29'b0_111111100001_101_0_101111111000;
      patterns[32526] = 29'b0_111111100001_110_0_111111100001;
      patterns[32527] = 29'b0_111111100001_111_0_111111100001;
      patterns[32528] = 29'b0_111111100010_000_0_111111100010;
      patterns[32529] = 29'b0_111111100010_001_0_100010111111;
      patterns[32530] = 29'b0_111111100010_010_1_111111000100;
      patterns[32531] = 29'b0_111111100010_011_1_111110001001;
      patterns[32532] = 29'b0_111111100010_100_0_011111110001;
      patterns[32533] = 29'b0_111111100010_101_1_001111111000;
      patterns[32534] = 29'b0_111111100010_110_0_111111100010;
      patterns[32535] = 29'b0_111111100010_111_0_111111100010;
      patterns[32536] = 29'b0_111111100011_000_0_111111100011;
      patterns[32537] = 29'b0_111111100011_001_0_100011111111;
      patterns[32538] = 29'b0_111111100011_010_1_111111000110;
      patterns[32539] = 29'b0_111111100011_011_1_111110001101;
      patterns[32540] = 29'b0_111111100011_100_1_011111110001;
      patterns[32541] = 29'b0_111111100011_101_1_101111111000;
      patterns[32542] = 29'b0_111111100011_110_0_111111100011;
      patterns[32543] = 29'b0_111111100011_111_0_111111100011;
      patterns[32544] = 29'b0_111111100100_000_0_111111100100;
      patterns[32545] = 29'b0_111111100100_001_0_100100111111;
      patterns[32546] = 29'b0_111111100100_010_1_111111001000;
      patterns[32547] = 29'b0_111111100100_011_1_111110010001;
      patterns[32548] = 29'b0_111111100100_100_0_011111110010;
      patterns[32549] = 29'b0_111111100100_101_0_001111111001;
      patterns[32550] = 29'b0_111111100100_110_0_111111100100;
      patterns[32551] = 29'b0_111111100100_111_0_111111100100;
      patterns[32552] = 29'b0_111111100101_000_0_111111100101;
      patterns[32553] = 29'b0_111111100101_001_0_100101111111;
      patterns[32554] = 29'b0_111111100101_010_1_111111001010;
      patterns[32555] = 29'b0_111111100101_011_1_111110010101;
      patterns[32556] = 29'b0_111111100101_100_1_011111110010;
      patterns[32557] = 29'b0_111111100101_101_0_101111111001;
      patterns[32558] = 29'b0_111111100101_110_0_111111100101;
      patterns[32559] = 29'b0_111111100101_111_0_111111100101;
      patterns[32560] = 29'b0_111111100110_000_0_111111100110;
      patterns[32561] = 29'b0_111111100110_001_0_100110111111;
      patterns[32562] = 29'b0_111111100110_010_1_111111001100;
      patterns[32563] = 29'b0_111111100110_011_1_111110011001;
      patterns[32564] = 29'b0_111111100110_100_0_011111110011;
      patterns[32565] = 29'b0_111111100110_101_1_001111111001;
      patterns[32566] = 29'b0_111111100110_110_0_111111100110;
      patterns[32567] = 29'b0_111111100110_111_0_111111100110;
      patterns[32568] = 29'b0_111111100111_000_0_111111100111;
      patterns[32569] = 29'b0_111111100111_001_0_100111111111;
      patterns[32570] = 29'b0_111111100111_010_1_111111001110;
      patterns[32571] = 29'b0_111111100111_011_1_111110011101;
      patterns[32572] = 29'b0_111111100111_100_1_011111110011;
      patterns[32573] = 29'b0_111111100111_101_1_101111111001;
      patterns[32574] = 29'b0_111111100111_110_0_111111100111;
      patterns[32575] = 29'b0_111111100111_111_0_111111100111;
      patterns[32576] = 29'b0_111111101000_000_0_111111101000;
      patterns[32577] = 29'b0_111111101000_001_0_101000111111;
      patterns[32578] = 29'b0_111111101000_010_1_111111010000;
      patterns[32579] = 29'b0_111111101000_011_1_111110100001;
      patterns[32580] = 29'b0_111111101000_100_0_011111110100;
      patterns[32581] = 29'b0_111111101000_101_0_001111111010;
      patterns[32582] = 29'b0_111111101000_110_0_111111101000;
      patterns[32583] = 29'b0_111111101000_111_0_111111101000;
      patterns[32584] = 29'b0_111111101001_000_0_111111101001;
      patterns[32585] = 29'b0_111111101001_001_0_101001111111;
      patterns[32586] = 29'b0_111111101001_010_1_111111010010;
      patterns[32587] = 29'b0_111111101001_011_1_111110100101;
      patterns[32588] = 29'b0_111111101001_100_1_011111110100;
      patterns[32589] = 29'b0_111111101001_101_0_101111111010;
      patterns[32590] = 29'b0_111111101001_110_0_111111101001;
      patterns[32591] = 29'b0_111111101001_111_0_111111101001;
      patterns[32592] = 29'b0_111111101010_000_0_111111101010;
      patterns[32593] = 29'b0_111111101010_001_0_101010111111;
      patterns[32594] = 29'b0_111111101010_010_1_111111010100;
      patterns[32595] = 29'b0_111111101010_011_1_111110101001;
      patterns[32596] = 29'b0_111111101010_100_0_011111110101;
      patterns[32597] = 29'b0_111111101010_101_1_001111111010;
      patterns[32598] = 29'b0_111111101010_110_0_111111101010;
      patterns[32599] = 29'b0_111111101010_111_0_111111101010;
      patterns[32600] = 29'b0_111111101011_000_0_111111101011;
      patterns[32601] = 29'b0_111111101011_001_0_101011111111;
      patterns[32602] = 29'b0_111111101011_010_1_111111010110;
      patterns[32603] = 29'b0_111111101011_011_1_111110101101;
      patterns[32604] = 29'b0_111111101011_100_1_011111110101;
      patterns[32605] = 29'b0_111111101011_101_1_101111111010;
      patterns[32606] = 29'b0_111111101011_110_0_111111101011;
      patterns[32607] = 29'b0_111111101011_111_0_111111101011;
      patterns[32608] = 29'b0_111111101100_000_0_111111101100;
      patterns[32609] = 29'b0_111111101100_001_0_101100111111;
      patterns[32610] = 29'b0_111111101100_010_1_111111011000;
      patterns[32611] = 29'b0_111111101100_011_1_111110110001;
      patterns[32612] = 29'b0_111111101100_100_0_011111110110;
      patterns[32613] = 29'b0_111111101100_101_0_001111111011;
      patterns[32614] = 29'b0_111111101100_110_0_111111101100;
      patterns[32615] = 29'b0_111111101100_111_0_111111101100;
      patterns[32616] = 29'b0_111111101101_000_0_111111101101;
      patterns[32617] = 29'b0_111111101101_001_0_101101111111;
      patterns[32618] = 29'b0_111111101101_010_1_111111011010;
      patterns[32619] = 29'b0_111111101101_011_1_111110110101;
      patterns[32620] = 29'b0_111111101101_100_1_011111110110;
      patterns[32621] = 29'b0_111111101101_101_0_101111111011;
      patterns[32622] = 29'b0_111111101101_110_0_111111101101;
      patterns[32623] = 29'b0_111111101101_111_0_111111101101;
      patterns[32624] = 29'b0_111111101110_000_0_111111101110;
      patterns[32625] = 29'b0_111111101110_001_0_101110111111;
      patterns[32626] = 29'b0_111111101110_010_1_111111011100;
      patterns[32627] = 29'b0_111111101110_011_1_111110111001;
      patterns[32628] = 29'b0_111111101110_100_0_011111110111;
      patterns[32629] = 29'b0_111111101110_101_1_001111111011;
      patterns[32630] = 29'b0_111111101110_110_0_111111101110;
      patterns[32631] = 29'b0_111111101110_111_0_111111101110;
      patterns[32632] = 29'b0_111111101111_000_0_111111101111;
      patterns[32633] = 29'b0_111111101111_001_0_101111111111;
      patterns[32634] = 29'b0_111111101111_010_1_111111011110;
      patterns[32635] = 29'b0_111111101111_011_1_111110111101;
      patterns[32636] = 29'b0_111111101111_100_1_011111110111;
      patterns[32637] = 29'b0_111111101111_101_1_101111111011;
      patterns[32638] = 29'b0_111111101111_110_0_111111101111;
      patterns[32639] = 29'b0_111111101111_111_0_111111101111;
      patterns[32640] = 29'b0_111111110000_000_0_111111110000;
      patterns[32641] = 29'b0_111111110000_001_0_110000111111;
      patterns[32642] = 29'b0_111111110000_010_1_111111100000;
      patterns[32643] = 29'b0_111111110000_011_1_111111000001;
      patterns[32644] = 29'b0_111111110000_100_0_011111111000;
      patterns[32645] = 29'b0_111111110000_101_0_001111111100;
      patterns[32646] = 29'b0_111111110000_110_0_111111110000;
      patterns[32647] = 29'b0_111111110000_111_0_111111110000;
      patterns[32648] = 29'b0_111111110001_000_0_111111110001;
      patterns[32649] = 29'b0_111111110001_001_0_110001111111;
      patterns[32650] = 29'b0_111111110001_010_1_111111100010;
      patterns[32651] = 29'b0_111111110001_011_1_111111000101;
      patterns[32652] = 29'b0_111111110001_100_1_011111111000;
      patterns[32653] = 29'b0_111111110001_101_0_101111111100;
      patterns[32654] = 29'b0_111111110001_110_0_111111110001;
      patterns[32655] = 29'b0_111111110001_111_0_111111110001;
      patterns[32656] = 29'b0_111111110010_000_0_111111110010;
      patterns[32657] = 29'b0_111111110010_001_0_110010111111;
      patterns[32658] = 29'b0_111111110010_010_1_111111100100;
      patterns[32659] = 29'b0_111111110010_011_1_111111001001;
      patterns[32660] = 29'b0_111111110010_100_0_011111111001;
      patterns[32661] = 29'b0_111111110010_101_1_001111111100;
      patterns[32662] = 29'b0_111111110010_110_0_111111110010;
      patterns[32663] = 29'b0_111111110010_111_0_111111110010;
      patterns[32664] = 29'b0_111111110011_000_0_111111110011;
      patterns[32665] = 29'b0_111111110011_001_0_110011111111;
      patterns[32666] = 29'b0_111111110011_010_1_111111100110;
      patterns[32667] = 29'b0_111111110011_011_1_111111001101;
      patterns[32668] = 29'b0_111111110011_100_1_011111111001;
      patterns[32669] = 29'b0_111111110011_101_1_101111111100;
      patterns[32670] = 29'b0_111111110011_110_0_111111110011;
      patterns[32671] = 29'b0_111111110011_111_0_111111110011;
      patterns[32672] = 29'b0_111111110100_000_0_111111110100;
      patterns[32673] = 29'b0_111111110100_001_0_110100111111;
      patterns[32674] = 29'b0_111111110100_010_1_111111101000;
      patterns[32675] = 29'b0_111111110100_011_1_111111010001;
      patterns[32676] = 29'b0_111111110100_100_0_011111111010;
      patterns[32677] = 29'b0_111111110100_101_0_001111111101;
      patterns[32678] = 29'b0_111111110100_110_0_111111110100;
      patterns[32679] = 29'b0_111111110100_111_0_111111110100;
      patterns[32680] = 29'b0_111111110101_000_0_111111110101;
      patterns[32681] = 29'b0_111111110101_001_0_110101111111;
      patterns[32682] = 29'b0_111111110101_010_1_111111101010;
      patterns[32683] = 29'b0_111111110101_011_1_111111010101;
      patterns[32684] = 29'b0_111111110101_100_1_011111111010;
      patterns[32685] = 29'b0_111111110101_101_0_101111111101;
      patterns[32686] = 29'b0_111111110101_110_0_111111110101;
      patterns[32687] = 29'b0_111111110101_111_0_111111110101;
      patterns[32688] = 29'b0_111111110110_000_0_111111110110;
      patterns[32689] = 29'b0_111111110110_001_0_110110111111;
      patterns[32690] = 29'b0_111111110110_010_1_111111101100;
      patterns[32691] = 29'b0_111111110110_011_1_111111011001;
      patterns[32692] = 29'b0_111111110110_100_0_011111111011;
      patterns[32693] = 29'b0_111111110110_101_1_001111111101;
      patterns[32694] = 29'b0_111111110110_110_0_111111110110;
      patterns[32695] = 29'b0_111111110110_111_0_111111110110;
      patterns[32696] = 29'b0_111111110111_000_0_111111110111;
      patterns[32697] = 29'b0_111111110111_001_0_110111111111;
      patterns[32698] = 29'b0_111111110111_010_1_111111101110;
      patterns[32699] = 29'b0_111111110111_011_1_111111011101;
      patterns[32700] = 29'b0_111111110111_100_1_011111111011;
      patterns[32701] = 29'b0_111111110111_101_1_101111111101;
      patterns[32702] = 29'b0_111111110111_110_0_111111110111;
      patterns[32703] = 29'b0_111111110111_111_0_111111110111;
      patterns[32704] = 29'b0_111111111000_000_0_111111111000;
      patterns[32705] = 29'b0_111111111000_001_0_111000111111;
      patterns[32706] = 29'b0_111111111000_010_1_111111110000;
      patterns[32707] = 29'b0_111111111000_011_1_111111100001;
      patterns[32708] = 29'b0_111111111000_100_0_011111111100;
      patterns[32709] = 29'b0_111111111000_101_0_001111111110;
      patterns[32710] = 29'b0_111111111000_110_0_111111111000;
      patterns[32711] = 29'b0_111111111000_111_0_111111111000;
      patterns[32712] = 29'b0_111111111001_000_0_111111111001;
      patterns[32713] = 29'b0_111111111001_001_0_111001111111;
      patterns[32714] = 29'b0_111111111001_010_1_111111110010;
      patterns[32715] = 29'b0_111111111001_011_1_111111100101;
      patterns[32716] = 29'b0_111111111001_100_1_011111111100;
      patterns[32717] = 29'b0_111111111001_101_0_101111111110;
      patterns[32718] = 29'b0_111111111001_110_0_111111111001;
      patterns[32719] = 29'b0_111111111001_111_0_111111111001;
      patterns[32720] = 29'b0_111111111010_000_0_111111111010;
      patterns[32721] = 29'b0_111111111010_001_0_111010111111;
      patterns[32722] = 29'b0_111111111010_010_1_111111110100;
      patterns[32723] = 29'b0_111111111010_011_1_111111101001;
      patterns[32724] = 29'b0_111111111010_100_0_011111111101;
      patterns[32725] = 29'b0_111111111010_101_1_001111111110;
      patterns[32726] = 29'b0_111111111010_110_0_111111111010;
      patterns[32727] = 29'b0_111111111010_111_0_111111111010;
      patterns[32728] = 29'b0_111111111011_000_0_111111111011;
      patterns[32729] = 29'b0_111111111011_001_0_111011111111;
      patterns[32730] = 29'b0_111111111011_010_1_111111110110;
      patterns[32731] = 29'b0_111111111011_011_1_111111101101;
      patterns[32732] = 29'b0_111111111011_100_1_011111111101;
      patterns[32733] = 29'b0_111111111011_101_1_101111111110;
      patterns[32734] = 29'b0_111111111011_110_0_111111111011;
      patterns[32735] = 29'b0_111111111011_111_0_111111111011;
      patterns[32736] = 29'b0_111111111100_000_0_111111111100;
      patterns[32737] = 29'b0_111111111100_001_0_111100111111;
      patterns[32738] = 29'b0_111111111100_010_1_111111111000;
      patterns[32739] = 29'b0_111111111100_011_1_111111110001;
      patterns[32740] = 29'b0_111111111100_100_0_011111111110;
      patterns[32741] = 29'b0_111111111100_101_0_001111111111;
      patterns[32742] = 29'b0_111111111100_110_0_111111111100;
      patterns[32743] = 29'b0_111111111100_111_0_111111111100;
      patterns[32744] = 29'b0_111111111101_000_0_111111111101;
      patterns[32745] = 29'b0_111111111101_001_0_111101111111;
      patterns[32746] = 29'b0_111111111101_010_1_111111111010;
      patterns[32747] = 29'b0_111111111101_011_1_111111110101;
      patterns[32748] = 29'b0_111111111101_100_1_011111111110;
      patterns[32749] = 29'b0_111111111101_101_0_101111111111;
      patterns[32750] = 29'b0_111111111101_110_0_111111111101;
      patterns[32751] = 29'b0_111111111101_111_0_111111111101;
      patterns[32752] = 29'b0_111111111110_000_0_111111111110;
      patterns[32753] = 29'b0_111111111110_001_0_111110111111;
      patterns[32754] = 29'b0_111111111110_010_1_111111111100;
      patterns[32755] = 29'b0_111111111110_011_1_111111111001;
      patterns[32756] = 29'b0_111111111110_100_0_011111111111;
      patterns[32757] = 29'b0_111111111110_101_1_001111111111;
      patterns[32758] = 29'b0_111111111110_110_0_111111111110;
      patterns[32759] = 29'b0_111111111110_111_0_111111111110;
      patterns[32760] = 29'b0_111111111111_000_0_111111111111;
      patterns[32761] = 29'b0_111111111111_001_0_111111111111;
      patterns[32762] = 29'b0_111111111111_010_1_111111111110;
      patterns[32763] = 29'b0_111111111111_011_1_111111111101;
      patterns[32764] = 29'b0_111111111111_100_1_011111111111;
      patterns[32765] = 29'b0_111111111111_101_1_101111111111;
      patterns[32766] = 29'b0_111111111111_110_0_111111111111;
      patterns[32767] = 29'b0_111111111111_111_0_111111111111;
      patterns[32768] = 29'b1_000000000000_000_1_000000000000;
      patterns[32769] = 29'b1_000000000000_001_1_000000000000;
      patterns[32770] = 29'b1_000000000000_010_0_000000000001;
      patterns[32771] = 29'b1_000000000000_011_0_000000000010;
      patterns[32772] = 29'b1_000000000000_100_0_100000000000;
      patterns[32773] = 29'b1_000000000000_101_0_010000000000;
      patterns[32774] = 29'b1_000000000000_110_1_000000000000;
      patterns[32775] = 29'b1_000000000000_111_1_000000000000;
      patterns[32776] = 29'b1_000000000001_000_1_000000000001;
      patterns[32777] = 29'b1_000000000001_001_1_000001000000;
      patterns[32778] = 29'b1_000000000001_010_0_000000000011;
      patterns[32779] = 29'b1_000000000001_011_0_000000000110;
      patterns[32780] = 29'b1_000000000001_100_1_100000000000;
      patterns[32781] = 29'b1_000000000001_101_0_110000000000;
      patterns[32782] = 29'b1_000000000001_110_1_000000000001;
      patterns[32783] = 29'b1_000000000001_111_1_000000000001;
      patterns[32784] = 29'b1_000000000010_000_1_000000000010;
      patterns[32785] = 29'b1_000000000010_001_1_000010000000;
      patterns[32786] = 29'b1_000000000010_010_0_000000000101;
      patterns[32787] = 29'b1_000000000010_011_0_000000001010;
      patterns[32788] = 29'b1_000000000010_100_0_100000000001;
      patterns[32789] = 29'b1_000000000010_101_1_010000000000;
      patterns[32790] = 29'b1_000000000010_110_1_000000000010;
      patterns[32791] = 29'b1_000000000010_111_1_000000000010;
      patterns[32792] = 29'b1_000000000011_000_1_000000000011;
      patterns[32793] = 29'b1_000000000011_001_1_000011000000;
      patterns[32794] = 29'b1_000000000011_010_0_000000000111;
      patterns[32795] = 29'b1_000000000011_011_0_000000001110;
      patterns[32796] = 29'b1_000000000011_100_1_100000000001;
      patterns[32797] = 29'b1_000000000011_101_1_110000000000;
      patterns[32798] = 29'b1_000000000011_110_1_000000000011;
      patterns[32799] = 29'b1_000000000011_111_1_000000000011;
      patterns[32800] = 29'b1_000000000100_000_1_000000000100;
      patterns[32801] = 29'b1_000000000100_001_1_000100000000;
      patterns[32802] = 29'b1_000000000100_010_0_000000001001;
      patterns[32803] = 29'b1_000000000100_011_0_000000010010;
      patterns[32804] = 29'b1_000000000100_100_0_100000000010;
      patterns[32805] = 29'b1_000000000100_101_0_010000000001;
      patterns[32806] = 29'b1_000000000100_110_1_000000000100;
      patterns[32807] = 29'b1_000000000100_111_1_000000000100;
      patterns[32808] = 29'b1_000000000101_000_1_000000000101;
      patterns[32809] = 29'b1_000000000101_001_1_000101000000;
      patterns[32810] = 29'b1_000000000101_010_0_000000001011;
      patterns[32811] = 29'b1_000000000101_011_0_000000010110;
      patterns[32812] = 29'b1_000000000101_100_1_100000000010;
      patterns[32813] = 29'b1_000000000101_101_0_110000000001;
      patterns[32814] = 29'b1_000000000101_110_1_000000000101;
      patterns[32815] = 29'b1_000000000101_111_1_000000000101;
      patterns[32816] = 29'b1_000000000110_000_1_000000000110;
      patterns[32817] = 29'b1_000000000110_001_1_000110000000;
      patterns[32818] = 29'b1_000000000110_010_0_000000001101;
      patterns[32819] = 29'b1_000000000110_011_0_000000011010;
      patterns[32820] = 29'b1_000000000110_100_0_100000000011;
      patterns[32821] = 29'b1_000000000110_101_1_010000000001;
      patterns[32822] = 29'b1_000000000110_110_1_000000000110;
      patterns[32823] = 29'b1_000000000110_111_1_000000000110;
      patterns[32824] = 29'b1_000000000111_000_1_000000000111;
      patterns[32825] = 29'b1_000000000111_001_1_000111000000;
      patterns[32826] = 29'b1_000000000111_010_0_000000001111;
      patterns[32827] = 29'b1_000000000111_011_0_000000011110;
      patterns[32828] = 29'b1_000000000111_100_1_100000000011;
      patterns[32829] = 29'b1_000000000111_101_1_110000000001;
      patterns[32830] = 29'b1_000000000111_110_1_000000000111;
      patterns[32831] = 29'b1_000000000111_111_1_000000000111;
      patterns[32832] = 29'b1_000000001000_000_1_000000001000;
      patterns[32833] = 29'b1_000000001000_001_1_001000000000;
      patterns[32834] = 29'b1_000000001000_010_0_000000010001;
      patterns[32835] = 29'b1_000000001000_011_0_000000100010;
      patterns[32836] = 29'b1_000000001000_100_0_100000000100;
      patterns[32837] = 29'b1_000000001000_101_0_010000000010;
      patterns[32838] = 29'b1_000000001000_110_1_000000001000;
      patterns[32839] = 29'b1_000000001000_111_1_000000001000;
      patterns[32840] = 29'b1_000000001001_000_1_000000001001;
      patterns[32841] = 29'b1_000000001001_001_1_001001000000;
      patterns[32842] = 29'b1_000000001001_010_0_000000010011;
      patterns[32843] = 29'b1_000000001001_011_0_000000100110;
      patterns[32844] = 29'b1_000000001001_100_1_100000000100;
      patterns[32845] = 29'b1_000000001001_101_0_110000000010;
      patterns[32846] = 29'b1_000000001001_110_1_000000001001;
      patterns[32847] = 29'b1_000000001001_111_1_000000001001;
      patterns[32848] = 29'b1_000000001010_000_1_000000001010;
      patterns[32849] = 29'b1_000000001010_001_1_001010000000;
      patterns[32850] = 29'b1_000000001010_010_0_000000010101;
      patterns[32851] = 29'b1_000000001010_011_0_000000101010;
      patterns[32852] = 29'b1_000000001010_100_0_100000000101;
      patterns[32853] = 29'b1_000000001010_101_1_010000000010;
      patterns[32854] = 29'b1_000000001010_110_1_000000001010;
      patterns[32855] = 29'b1_000000001010_111_1_000000001010;
      patterns[32856] = 29'b1_000000001011_000_1_000000001011;
      patterns[32857] = 29'b1_000000001011_001_1_001011000000;
      patterns[32858] = 29'b1_000000001011_010_0_000000010111;
      patterns[32859] = 29'b1_000000001011_011_0_000000101110;
      patterns[32860] = 29'b1_000000001011_100_1_100000000101;
      patterns[32861] = 29'b1_000000001011_101_1_110000000010;
      patterns[32862] = 29'b1_000000001011_110_1_000000001011;
      patterns[32863] = 29'b1_000000001011_111_1_000000001011;
      patterns[32864] = 29'b1_000000001100_000_1_000000001100;
      patterns[32865] = 29'b1_000000001100_001_1_001100000000;
      patterns[32866] = 29'b1_000000001100_010_0_000000011001;
      patterns[32867] = 29'b1_000000001100_011_0_000000110010;
      patterns[32868] = 29'b1_000000001100_100_0_100000000110;
      patterns[32869] = 29'b1_000000001100_101_0_010000000011;
      patterns[32870] = 29'b1_000000001100_110_1_000000001100;
      patterns[32871] = 29'b1_000000001100_111_1_000000001100;
      patterns[32872] = 29'b1_000000001101_000_1_000000001101;
      patterns[32873] = 29'b1_000000001101_001_1_001101000000;
      patterns[32874] = 29'b1_000000001101_010_0_000000011011;
      patterns[32875] = 29'b1_000000001101_011_0_000000110110;
      patterns[32876] = 29'b1_000000001101_100_1_100000000110;
      patterns[32877] = 29'b1_000000001101_101_0_110000000011;
      patterns[32878] = 29'b1_000000001101_110_1_000000001101;
      patterns[32879] = 29'b1_000000001101_111_1_000000001101;
      patterns[32880] = 29'b1_000000001110_000_1_000000001110;
      patterns[32881] = 29'b1_000000001110_001_1_001110000000;
      patterns[32882] = 29'b1_000000001110_010_0_000000011101;
      patterns[32883] = 29'b1_000000001110_011_0_000000111010;
      patterns[32884] = 29'b1_000000001110_100_0_100000000111;
      patterns[32885] = 29'b1_000000001110_101_1_010000000011;
      patterns[32886] = 29'b1_000000001110_110_1_000000001110;
      patterns[32887] = 29'b1_000000001110_111_1_000000001110;
      patterns[32888] = 29'b1_000000001111_000_1_000000001111;
      patterns[32889] = 29'b1_000000001111_001_1_001111000000;
      patterns[32890] = 29'b1_000000001111_010_0_000000011111;
      patterns[32891] = 29'b1_000000001111_011_0_000000111110;
      patterns[32892] = 29'b1_000000001111_100_1_100000000111;
      patterns[32893] = 29'b1_000000001111_101_1_110000000011;
      patterns[32894] = 29'b1_000000001111_110_1_000000001111;
      patterns[32895] = 29'b1_000000001111_111_1_000000001111;
      patterns[32896] = 29'b1_000000010000_000_1_000000010000;
      patterns[32897] = 29'b1_000000010000_001_1_010000000000;
      patterns[32898] = 29'b1_000000010000_010_0_000000100001;
      patterns[32899] = 29'b1_000000010000_011_0_000001000010;
      patterns[32900] = 29'b1_000000010000_100_0_100000001000;
      patterns[32901] = 29'b1_000000010000_101_0_010000000100;
      patterns[32902] = 29'b1_000000010000_110_1_000000010000;
      patterns[32903] = 29'b1_000000010000_111_1_000000010000;
      patterns[32904] = 29'b1_000000010001_000_1_000000010001;
      patterns[32905] = 29'b1_000000010001_001_1_010001000000;
      patterns[32906] = 29'b1_000000010001_010_0_000000100011;
      patterns[32907] = 29'b1_000000010001_011_0_000001000110;
      patterns[32908] = 29'b1_000000010001_100_1_100000001000;
      patterns[32909] = 29'b1_000000010001_101_0_110000000100;
      patterns[32910] = 29'b1_000000010001_110_1_000000010001;
      patterns[32911] = 29'b1_000000010001_111_1_000000010001;
      patterns[32912] = 29'b1_000000010010_000_1_000000010010;
      patterns[32913] = 29'b1_000000010010_001_1_010010000000;
      patterns[32914] = 29'b1_000000010010_010_0_000000100101;
      patterns[32915] = 29'b1_000000010010_011_0_000001001010;
      patterns[32916] = 29'b1_000000010010_100_0_100000001001;
      patterns[32917] = 29'b1_000000010010_101_1_010000000100;
      patterns[32918] = 29'b1_000000010010_110_1_000000010010;
      patterns[32919] = 29'b1_000000010010_111_1_000000010010;
      patterns[32920] = 29'b1_000000010011_000_1_000000010011;
      patterns[32921] = 29'b1_000000010011_001_1_010011000000;
      patterns[32922] = 29'b1_000000010011_010_0_000000100111;
      patterns[32923] = 29'b1_000000010011_011_0_000001001110;
      patterns[32924] = 29'b1_000000010011_100_1_100000001001;
      patterns[32925] = 29'b1_000000010011_101_1_110000000100;
      patterns[32926] = 29'b1_000000010011_110_1_000000010011;
      patterns[32927] = 29'b1_000000010011_111_1_000000010011;
      patterns[32928] = 29'b1_000000010100_000_1_000000010100;
      patterns[32929] = 29'b1_000000010100_001_1_010100000000;
      patterns[32930] = 29'b1_000000010100_010_0_000000101001;
      patterns[32931] = 29'b1_000000010100_011_0_000001010010;
      patterns[32932] = 29'b1_000000010100_100_0_100000001010;
      patterns[32933] = 29'b1_000000010100_101_0_010000000101;
      patterns[32934] = 29'b1_000000010100_110_1_000000010100;
      patterns[32935] = 29'b1_000000010100_111_1_000000010100;
      patterns[32936] = 29'b1_000000010101_000_1_000000010101;
      patterns[32937] = 29'b1_000000010101_001_1_010101000000;
      patterns[32938] = 29'b1_000000010101_010_0_000000101011;
      patterns[32939] = 29'b1_000000010101_011_0_000001010110;
      patterns[32940] = 29'b1_000000010101_100_1_100000001010;
      patterns[32941] = 29'b1_000000010101_101_0_110000000101;
      patterns[32942] = 29'b1_000000010101_110_1_000000010101;
      patterns[32943] = 29'b1_000000010101_111_1_000000010101;
      patterns[32944] = 29'b1_000000010110_000_1_000000010110;
      patterns[32945] = 29'b1_000000010110_001_1_010110000000;
      patterns[32946] = 29'b1_000000010110_010_0_000000101101;
      patterns[32947] = 29'b1_000000010110_011_0_000001011010;
      patterns[32948] = 29'b1_000000010110_100_0_100000001011;
      patterns[32949] = 29'b1_000000010110_101_1_010000000101;
      patterns[32950] = 29'b1_000000010110_110_1_000000010110;
      patterns[32951] = 29'b1_000000010110_111_1_000000010110;
      patterns[32952] = 29'b1_000000010111_000_1_000000010111;
      patterns[32953] = 29'b1_000000010111_001_1_010111000000;
      patterns[32954] = 29'b1_000000010111_010_0_000000101111;
      patterns[32955] = 29'b1_000000010111_011_0_000001011110;
      patterns[32956] = 29'b1_000000010111_100_1_100000001011;
      patterns[32957] = 29'b1_000000010111_101_1_110000000101;
      patterns[32958] = 29'b1_000000010111_110_1_000000010111;
      patterns[32959] = 29'b1_000000010111_111_1_000000010111;
      patterns[32960] = 29'b1_000000011000_000_1_000000011000;
      patterns[32961] = 29'b1_000000011000_001_1_011000000000;
      patterns[32962] = 29'b1_000000011000_010_0_000000110001;
      patterns[32963] = 29'b1_000000011000_011_0_000001100010;
      patterns[32964] = 29'b1_000000011000_100_0_100000001100;
      patterns[32965] = 29'b1_000000011000_101_0_010000000110;
      patterns[32966] = 29'b1_000000011000_110_1_000000011000;
      patterns[32967] = 29'b1_000000011000_111_1_000000011000;
      patterns[32968] = 29'b1_000000011001_000_1_000000011001;
      patterns[32969] = 29'b1_000000011001_001_1_011001000000;
      patterns[32970] = 29'b1_000000011001_010_0_000000110011;
      patterns[32971] = 29'b1_000000011001_011_0_000001100110;
      patterns[32972] = 29'b1_000000011001_100_1_100000001100;
      patterns[32973] = 29'b1_000000011001_101_0_110000000110;
      patterns[32974] = 29'b1_000000011001_110_1_000000011001;
      patterns[32975] = 29'b1_000000011001_111_1_000000011001;
      patterns[32976] = 29'b1_000000011010_000_1_000000011010;
      patterns[32977] = 29'b1_000000011010_001_1_011010000000;
      patterns[32978] = 29'b1_000000011010_010_0_000000110101;
      patterns[32979] = 29'b1_000000011010_011_0_000001101010;
      patterns[32980] = 29'b1_000000011010_100_0_100000001101;
      patterns[32981] = 29'b1_000000011010_101_1_010000000110;
      patterns[32982] = 29'b1_000000011010_110_1_000000011010;
      patterns[32983] = 29'b1_000000011010_111_1_000000011010;
      patterns[32984] = 29'b1_000000011011_000_1_000000011011;
      patterns[32985] = 29'b1_000000011011_001_1_011011000000;
      patterns[32986] = 29'b1_000000011011_010_0_000000110111;
      patterns[32987] = 29'b1_000000011011_011_0_000001101110;
      patterns[32988] = 29'b1_000000011011_100_1_100000001101;
      patterns[32989] = 29'b1_000000011011_101_1_110000000110;
      patterns[32990] = 29'b1_000000011011_110_1_000000011011;
      patterns[32991] = 29'b1_000000011011_111_1_000000011011;
      patterns[32992] = 29'b1_000000011100_000_1_000000011100;
      patterns[32993] = 29'b1_000000011100_001_1_011100000000;
      patterns[32994] = 29'b1_000000011100_010_0_000000111001;
      patterns[32995] = 29'b1_000000011100_011_0_000001110010;
      patterns[32996] = 29'b1_000000011100_100_0_100000001110;
      patterns[32997] = 29'b1_000000011100_101_0_010000000111;
      patterns[32998] = 29'b1_000000011100_110_1_000000011100;
      patterns[32999] = 29'b1_000000011100_111_1_000000011100;
      patterns[33000] = 29'b1_000000011101_000_1_000000011101;
      patterns[33001] = 29'b1_000000011101_001_1_011101000000;
      patterns[33002] = 29'b1_000000011101_010_0_000000111011;
      patterns[33003] = 29'b1_000000011101_011_0_000001110110;
      patterns[33004] = 29'b1_000000011101_100_1_100000001110;
      patterns[33005] = 29'b1_000000011101_101_0_110000000111;
      patterns[33006] = 29'b1_000000011101_110_1_000000011101;
      patterns[33007] = 29'b1_000000011101_111_1_000000011101;
      patterns[33008] = 29'b1_000000011110_000_1_000000011110;
      patterns[33009] = 29'b1_000000011110_001_1_011110000000;
      patterns[33010] = 29'b1_000000011110_010_0_000000111101;
      patterns[33011] = 29'b1_000000011110_011_0_000001111010;
      patterns[33012] = 29'b1_000000011110_100_0_100000001111;
      patterns[33013] = 29'b1_000000011110_101_1_010000000111;
      patterns[33014] = 29'b1_000000011110_110_1_000000011110;
      patterns[33015] = 29'b1_000000011110_111_1_000000011110;
      patterns[33016] = 29'b1_000000011111_000_1_000000011111;
      patterns[33017] = 29'b1_000000011111_001_1_011111000000;
      patterns[33018] = 29'b1_000000011111_010_0_000000111111;
      patterns[33019] = 29'b1_000000011111_011_0_000001111110;
      patterns[33020] = 29'b1_000000011111_100_1_100000001111;
      patterns[33021] = 29'b1_000000011111_101_1_110000000111;
      patterns[33022] = 29'b1_000000011111_110_1_000000011111;
      patterns[33023] = 29'b1_000000011111_111_1_000000011111;
      patterns[33024] = 29'b1_000000100000_000_1_000000100000;
      patterns[33025] = 29'b1_000000100000_001_1_100000000000;
      patterns[33026] = 29'b1_000000100000_010_0_000001000001;
      patterns[33027] = 29'b1_000000100000_011_0_000010000010;
      patterns[33028] = 29'b1_000000100000_100_0_100000010000;
      patterns[33029] = 29'b1_000000100000_101_0_010000001000;
      patterns[33030] = 29'b1_000000100000_110_1_000000100000;
      patterns[33031] = 29'b1_000000100000_111_1_000000100000;
      patterns[33032] = 29'b1_000000100001_000_1_000000100001;
      patterns[33033] = 29'b1_000000100001_001_1_100001000000;
      patterns[33034] = 29'b1_000000100001_010_0_000001000011;
      patterns[33035] = 29'b1_000000100001_011_0_000010000110;
      patterns[33036] = 29'b1_000000100001_100_1_100000010000;
      patterns[33037] = 29'b1_000000100001_101_0_110000001000;
      patterns[33038] = 29'b1_000000100001_110_1_000000100001;
      patterns[33039] = 29'b1_000000100001_111_1_000000100001;
      patterns[33040] = 29'b1_000000100010_000_1_000000100010;
      patterns[33041] = 29'b1_000000100010_001_1_100010000000;
      patterns[33042] = 29'b1_000000100010_010_0_000001000101;
      patterns[33043] = 29'b1_000000100010_011_0_000010001010;
      patterns[33044] = 29'b1_000000100010_100_0_100000010001;
      patterns[33045] = 29'b1_000000100010_101_1_010000001000;
      patterns[33046] = 29'b1_000000100010_110_1_000000100010;
      patterns[33047] = 29'b1_000000100010_111_1_000000100010;
      patterns[33048] = 29'b1_000000100011_000_1_000000100011;
      patterns[33049] = 29'b1_000000100011_001_1_100011000000;
      patterns[33050] = 29'b1_000000100011_010_0_000001000111;
      patterns[33051] = 29'b1_000000100011_011_0_000010001110;
      patterns[33052] = 29'b1_000000100011_100_1_100000010001;
      patterns[33053] = 29'b1_000000100011_101_1_110000001000;
      patterns[33054] = 29'b1_000000100011_110_1_000000100011;
      patterns[33055] = 29'b1_000000100011_111_1_000000100011;
      patterns[33056] = 29'b1_000000100100_000_1_000000100100;
      patterns[33057] = 29'b1_000000100100_001_1_100100000000;
      patterns[33058] = 29'b1_000000100100_010_0_000001001001;
      patterns[33059] = 29'b1_000000100100_011_0_000010010010;
      patterns[33060] = 29'b1_000000100100_100_0_100000010010;
      patterns[33061] = 29'b1_000000100100_101_0_010000001001;
      patterns[33062] = 29'b1_000000100100_110_1_000000100100;
      patterns[33063] = 29'b1_000000100100_111_1_000000100100;
      patterns[33064] = 29'b1_000000100101_000_1_000000100101;
      patterns[33065] = 29'b1_000000100101_001_1_100101000000;
      patterns[33066] = 29'b1_000000100101_010_0_000001001011;
      patterns[33067] = 29'b1_000000100101_011_0_000010010110;
      patterns[33068] = 29'b1_000000100101_100_1_100000010010;
      patterns[33069] = 29'b1_000000100101_101_0_110000001001;
      patterns[33070] = 29'b1_000000100101_110_1_000000100101;
      patterns[33071] = 29'b1_000000100101_111_1_000000100101;
      patterns[33072] = 29'b1_000000100110_000_1_000000100110;
      patterns[33073] = 29'b1_000000100110_001_1_100110000000;
      patterns[33074] = 29'b1_000000100110_010_0_000001001101;
      patterns[33075] = 29'b1_000000100110_011_0_000010011010;
      patterns[33076] = 29'b1_000000100110_100_0_100000010011;
      patterns[33077] = 29'b1_000000100110_101_1_010000001001;
      patterns[33078] = 29'b1_000000100110_110_1_000000100110;
      patterns[33079] = 29'b1_000000100110_111_1_000000100110;
      patterns[33080] = 29'b1_000000100111_000_1_000000100111;
      patterns[33081] = 29'b1_000000100111_001_1_100111000000;
      patterns[33082] = 29'b1_000000100111_010_0_000001001111;
      patterns[33083] = 29'b1_000000100111_011_0_000010011110;
      patterns[33084] = 29'b1_000000100111_100_1_100000010011;
      patterns[33085] = 29'b1_000000100111_101_1_110000001001;
      patterns[33086] = 29'b1_000000100111_110_1_000000100111;
      patterns[33087] = 29'b1_000000100111_111_1_000000100111;
      patterns[33088] = 29'b1_000000101000_000_1_000000101000;
      patterns[33089] = 29'b1_000000101000_001_1_101000000000;
      patterns[33090] = 29'b1_000000101000_010_0_000001010001;
      patterns[33091] = 29'b1_000000101000_011_0_000010100010;
      patterns[33092] = 29'b1_000000101000_100_0_100000010100;
      patterns[33093] = 29'b1_000000101000_101_0_010000001010;
      patterns[33094] = 29'b1_000000101000_110_1_000000101000;
      patterns[33095] = 29'b1_000000101000_111_1_000000101000;
      patterns[33096] = 29'b1_000000101001_000_1_000000101001;
      patterns[33097] = 29'b1_000000101001_001_1_101001000000;
      patterns[33098] = 29'b1_000000101001_010_0_000001010011;
      patterns[33099] = 29'b1_000000101001_011_0_000010100110;
      patterns[33100] = 29'b1_000000101001_100_1_100000010100;
      patterns[33101] = 29'b1_000000101001_101_0_110000001010;
      patterns[33102] = 29'b1_000000101001_110_1_000000101001;
      patterns[33103] = 29'b1_000000101001_111_1_000000101001;
      patterns[33104] = 29'b1_000000101010_000_1_000000101010;
      patterns[33105] = 29'b1_000000101010_001_1_101010000000;
      patterns[33106] = 29'b1_000000101010_010_0_000001010101;
      patterns[33107] = 29'b1_000000101010_011_0_000010101010;
      patterns[33108] = 29'b1_000000101010_100_0_100000010101;
      patterns[33109] = 29'b1_000000101010_101_1_010000001010;
      patterns[33110] = 29'b1_000000101010_110_1_000000101010;
      patterns[33111] = 29'b1_000000101010_111_1_000000101010;
      patterns[33112] = 29'b1_000000101011_000_1_000000101011;
      patterns[33113] = 29'b1_000000101011_001_1_101011000000;
      patterns[33114] = 29'b1_000000101011_010_0_000001010111;
      patterns[33115] = 29'b1_000000101011_011_0_000010101110;
      patterns[33116] = 29'b1_000000101011_100_1_100000010101;
      patterns[33117] = 29'b1_000000101011_101_1_110000001010;
      patterns[33118] = 29'b1_000000101011_110_1_000000101011;
      patterns[33119] = 29'b1_000000101011_111_1_000000101011;
      patterns[33120] = 29'b1_000000101100_000_1_000000101100;
      patterns[33121] = 29'b1_000000101100_001_1_101100000000;
      patterns[33122] = 29'b1_000000101100_010_0_000001011001;
      patterns[33123] = 29'b1_000000101100_011_0_000010110010;
      patterns[33124] = 29'b1_000000101100_100_0_100000010110;
      patterns[33125] = 29'b1_000000101100_101_0_010000001011;
      patterns[33126] = 29'b1_000000101100_110_1_000000101100;
      patterns[33127] = 29'b1_000000101100_111_1_000000101100;
      patterns[33128] = 29'b1_000000101101_000_1_000000101101;
      patterns[33129] = 29'b1_000000101101_001_1_101101000000;
      patterns[33130] = 29'b1_000000101101_010_0_000001011011;
      patterns[33131] = 29'b1_000000101101_011_0_000010110110;
      patterns[33132] = 29'b1_000000101101_100_1_100000010110;
      patterns[33133] = 29'b1_000000101101_101_0_110000001011;
      patterns[33134] = 29'b1_000000101101_110_1_000000101101;
      patterns[33135] = 29'b1_000000101101_111_1_000000101101;
      patterns[33136] = 29'b1_000000101110_000_1_000000101110;
      patterns[33137] = 29'b1_000000101110_001_1_101110000000;
      patterns[33138] = 29'b1_000000101110_010_0_000001011101;
      patterns[33139] = 29'b1_000000101110_011_0_000010111010;
      patterns[33140] = 29'b1_000000101110_100_0_100000010111;
      patterns[33141] = 29'b1_000000101110_101_1_010000001011;
      patterns[33142] = 29'b1_000000101110_110_1_000000101110;
      patterns[33143] = 29'b1_000000101110_111_1_000000101110;
      patterns[33144] = 29'b1_000000101111_000_1_000000101111;
      patterns[33145] = 29'b1_000000101111_001_1_101111000000;
      patterns[33146] = 29'b1_000000101111_010_0_000001011111;
      patterns[33147] = 29'b1_000000101111_011_0_000010111110;
      patterns[33148] = 29'b1_000000101111_100_1_100000010111;
      patterns[33149] = 29'b1_000000101111_101_1_110000001011;
      patterns[33150] = 29'b1_000000101111_110_1_000000101111;
      patterns[33151] = 29'b1_000000101111_111_1_000000101111;
      patterns[33152] = 29'b1_000000110000_000_1_000000110000;
      patterns[33153] = 29'b1_000000110000_001_1_110000000000;
      patterns[33154] = 29'b1_000000110000_010_0_000001100001;
      patterns[33155] = 29'b1_000000110000_011_0_000011000010;
      patterns[33156] = 29'b1_000000110000_100_0_100000011000;
      patterns[33157] = 29'b1_000000110000_101_0_010000001100;
      patterns[33158] = 29'b1_000000110000_110_1_000000110000;
      patterns[33159] = 29'b1_000000110000_111_1_000000110000;
      patterns[33160] = 29'b1_000000110001_000_1_000000110001;
      patterns[33161] = 29'b1_000000110001_001_1_110001000000;
      patterns[33162] = 29'b1_000000110001_010_0_000001100011;
      patterns[33163] = 29'b1_000000110001_011_0_000011000110;
      patterns[33164] = 29'b1_000000110001_100_1_100000011000;
      patterns[33165] = 29'b1_000000110001_101_0_110000001100;
      patterns[33166] = 29'b1_000000110001_110_1_000000110001;
      patterns[33167] = 29'b1_000000110001_111_1_000000110001;
      patterns[33168] = 29'b1_000000110010_000_1_000000110010;
      patterns[33169] = 29'b1_000000110010_001_1_110010000000;
      patterns[33170] = 29'b1_000000110010_010_0_000001100101;
      patterns[33171] = 29'b1_000000110010_011_0_000011001010;
      patterns[33172] = 29'b1_000000110010_100_0_100000011001;
      patterns[33173] = 29'b1_000000110010_101_1_010000001100;
      patterns[33174] = 29'b1_000000110010_110_1_000000110010;
      patterns[33175] = 29'b1_000000110010_111_1_000000110010;
      patterns[33176] = 29'b1_000000110011_000_1_000000110011;
      patterns[33177] = 29'b1_000000110011_001_1_110011000000;
      patterns[33178] = 29'b1_000000110011_010_0_000001100111;
      patterns[33179] = 29'b1_000000110011_011_0_000011001110;
      patterns[33180] = 29'b1_000000110011_100_1_100000011001;
      patterns[33181] = 29'b1_000000110011_101_1_110000001100;
      patterns[33182] = 29'b1_000000110011_110_1_000000110011;
      patterns[33183] = 29'b1_000000110011_111_1_000000110011;
      patterns[33184] = 29'b1_000000110100_000_1_000000110100;
      patterns[33185] = 29'b1_000000110100_001_1_110100000000;
      patterns[33186] = 29'b1_000000110100_010_0_000001101001;
      patterns[33187] = 29'b1_000000110100_011_0_000011010010;
      patterns[33188] = 29'b1_000000110100_100_0_100000011010;
      patterns[33189] = 29'b1_000000110100_101_0_010000001101;
      patterns[33190] = 29'b1_000000110100_110_1_000000110100;
      patterns[33191] = 29'b1_000000110100_111_1_000000110100;
      patterns[33192] = 29'b1_000000110101_000_1_000000110101;
      patterns[33193] = 29'b1_000000110101_001_1_110101000000;
      patterns[33194] = 29'b1_000000110101_010_0_000001101011;
      patterns[33195] = 29'b1_000000110101_011_0_000011010110;
      patterns[33196] = 29'b1_000000110101_100_1_100000011010;
      patterns[33197] = 29'b1_000000110101_101_0_110000001101;
      patterns[33198] = 29'b1_000000110101_110_1_000000110101;
      patterns[33199] = 29'b1_000000110101_111_1_000000110101;
      patterns[33200] = 29'b1_000000110110_000_1_000000110110;
      patterns[33201] = 29'b1_000000110110_001_1_110110000000;
      patterns[33202] = 29'b1_000000110110_010_0_000001101101;
      patterns[33203] = 29'b1_000000110110_011_0_000011011010;
      patterns[33204] = 29'b1_000000110110_100_0_100000011011;
      patterns[33205] = 29'b1_000000110110_101_1_010000001101;
      patterns[33206] = 29'b1_000000110110_110_1_000000110110;
      patterns[33207] = 29'b1_000000110110_111_1_000000110110;
      patterns[33208] = 29'b1_000000110111_000_1_000000110111;
      patterns[33209] = 29'b1_000000110111_001_1_110111000000;
      patterns[33210] = 29'b1_000000110111_010_0_000001101111;
      patterns[33211] = 29'b1_000000110111_011_0_000011011110;
      patterns[33212] = 29'b1_000000110111_100_1_100000011011;
      patterns[33213] = 29'b1_000000110111_101_1_110000001101;
      patterns[33214] = 29'b1_000000110111_110_1_000000110111;
      patterns[33215] = 29'b1_000000110111_111_1_000000110111;
      patterns[33216] = 29'b1_000000111000_000_1_000000111000;
      patterns[33217] = 29'b1_000000111000_001_1_111000000000;
      patterns[33218] = 29'b1_000000111000_010_0_000001110001;
      patterns[33219] = 29'b1_000000111000_011_0_000011100010;
      patterns[33220] = 29'b1_000000111000_100_0_100000011100;
      patterns[33221] = 29'b1_000000111000_101_0_010000001110;
      patterns[33222] = 29'b1_000000111000_110_1_000000111000;
      patterns[33223] = 29'b1_000000111000_111_1_000000111000;
      patterns[33224] = 29'b1_000000111001_000_1_000000111001;
      patterns[33225] = 29'b1_000000111001_001_1_111001000000;
      patterns[33226] = 29'b1_000000111001_010_0_000001110011;
      patterns[33227] = 29'b1_000000111001_011_0_000011100110;
      patterns[33228] = 29'b1_000000111001_100_1_100000011100;
      patterns[33229] = 29'b1_000000111001_101_0_110000001110;
      patterns[33230] = 29'b1_000000111001_110_1_000000111001;
      patterns[33231] = 29'b1_000000111001_111_1_000000111001;
      patterns[33232] = 29'b1_000000111010_000_1_000000111010;
      patterns[33233] = 29'b1_000000111010_001_1_111010000000;
      patterns[33234] = 29'b1_000000111010_010_0_000001110101;
      patterns[33235] = 29'b1_000000111010_011_0_000011101010;
      patterns[33236] = 29'b1_000000111010_100_0_100000011101;
      patterns[33237] = 29'b1_000000111010_101_1_010000001110;
      patterns[33238] = 29'b1_000000111010_110_1_000000111010;
      patterns[33239] = 29'b1_000000111010_111_1_000000111010;
      patterns[33240] = 29'b1_000000111011_000_1_000000111011;
      patterns[33241] = 29'b1_000000111011_001_1_111011000000;
      patterns[33242] = 29'b1_000000111011_010_0_000001110111;
      patterns[33243] = 29'b1_000000111011_011_0_000011101110;
      patterns[33244] = 29'b1_000000111011_100_1_100000011101;
      patterns[33245] = 29'b1_000000111011_101_1_110000001110;
      patterns[33246] = 29'b1_000000111011_110_1_000000111011;
      patterns[33247] = 29'b1_000000111011_111_1_000000111011;
      patterns[33248] = 29'b1_000000111100_000_1_000000111100;
      patterns[33249] = 29'b1_000000111100_001_1_111100000000;
      patterns[33250] = 29'b1_000000111100_010_0_000001111001;
      patterns[33251] = 29'b1_000000111100_011_0_000011110010;
      patterns[33252] = 29'b1_000000111100_100_0_100000011110;
      patterns[33253] = 29'b1_000000111100_101_0_010000001111;
      patterns[33254] = 29'b1_000000111100_110_1_000000111100;
      patterns[33255] = 29'b1_000000111100_111_1_000000111100;
      patterns[33256] = 29'b1_000000111101_000_1_000000111101;
      patterns[33257] = 29'b1_000000111101_001_1_111101000000;
      patterns[33258] = 29'b1_000000111101_010_0_000001111011;
      patterns[33259] = 29'b1_000000111101_011_0_000011110110;
      patterns[33260] = 29'b1_000000111101_100_1_100000011110;
      patterns[33261] = 29'b1_000000111101_101_0_110000001111;
      patterns[33262] = 29'b1_000000111101_110_1_000000111101;
      patterns[33263] = 29'b1_000000111101_111_1_000000111101;
      patterns[33264] = 29'b1_000000111110_000_1_000000111110;
      patterns[33265] = 29'b1_000000111110_001_1_111110000000;
      patterns[33266] = 29'b1_000000111110_010_0_000001111101;
      patterns[33267] = 29'b1_000000111110_011_0_000011111010;
      patterns[33268] = 29'b1_000000111110_100_0_100000011111;
      patterns[33269] = 29'b1_000000111110_101_1_010000001111;
      patterns[33270] = 29'b1_000000111110_110_1_000000111110;
      patterns[33271] = 29'b1_000000111110_111_1_000000111110;
      patterns[33272] = 29'b1_000000111111_000_1_000000111111;
      patterns[33273] = 29'b1_000000111111_001_1_111111000000;
      patterns[33274] = 29'b1_000000111111_010_0_000001111111;
      patterns[33275] = 29'b1_000000111111_011_0_000011111110;
      patterns[33276] = 29'b1_000000111111_100_1_100000011111;
      patterns[33277] = 29'b1_000000111111_101_1_110000001111;
      patterns[33278] = 29'b1_000000111111_110_1_000000111111;
      patterns[33279] = 29'b1_000000111111_111_1_000000111111;
      patterns[33280] = 29'b1_000001000000_000_1_000001000000;
      patterns[33281] = 29'b1_000001000000_001_1_000000000001;
      patterns[33282] = 29'b1_000001000000_010_0_000010000001;
      patterns[33283] = 29'b1_000001000000_011_0_000100000010;
      patterns[33284] = 29'b1_000001000000_100_0_100000100000;
      patterns[33285] = 29'b1_000001000000_101_0_010000010000;
      patterns[33286] = 29'b1_000001000000_110_1_000001000000;
      patterns[33287] = 29'b1_000001000000_111_1_000001000000;
      patterns[33288] = 29'b1_000001000001_000_1_000001000001;
      patterns[33289] = 29'b1_000001000001_001_1_000001000001;
      patterns[33290] = 29'b1_000001000001_010_0_000010000011;
      patterns[33291] = 29'b1_000001000001_011_0_000100000110;
      patterns[33292] = 29'b1_000001000001_100_1_100000100000;
      patterns[33293] = 29'b1_000001000001_101_0_110000010000;
      patterns[33294] = 29'b1_000001000001_110_1_000001000001;
      patterns[33295] = 29'b1_000001000001_111_1_000001000001;
      patterns[33296] = 29'b1_000001000010_000_1_000001000010;
      patterns[33297] = 29'b1_000001000010_001_1_000010000001;
      patterns[33298] = 29'b1_000001000010_010_0_000010000101;
      patterns[33299] = 29'b1_000001000010_011_0_000100001010;
      patterns[33300] = 29'b1_000001000010_100_0_100000100001;
      patterns[33301] = 29'b1_000001000010_101_1_010000010000;
      patterns[33302] = 29'b1_000001000010_110_1_000001000010;
      patterns[33303] = 29'b1_000001000010_111_1_000001000010;
      patterns[33304] = 29'b1_000001000011_000_1_000001000011;
      patterns[33305] = 29'b1_000001000011_001_1_000011000001;
      patterns[33306] = 29'b1_000001000011_010_0_000010000111;
      patterns[33307] = 29'b1_000001000011_011_0_000100001110;
      patterns[33308] = 29'b1_000001000011_100_1_100000100001;
      patterns[33309] = 29'b1_000001000011_101_1_110000010000;
      patterns[33310] = 29'b1_000001000011_110_1_000001000011;
      patterns[33311] = 29'b1_000001000011_111_1_000001000011;
      patterns[33312] = 29'b1_000001000100_000_1_000001000100;
      patterns[33313] = 29'b1_000001000100_001_1_000100000001;
      patterns[33314] = 29'b1_000001000100_010_0_000010001001;
      patterns[33315] = 29'b1_000001000100_011_0_000100010010;
      patterns[33316] = 29'b1_000001000100_100_0_100000100010;
      patterns[33317] = 29'b1_000001000100_101_0_010000010001;
      patterns[33318] = 29'b1_000001000100_110_1_000001000100;
      patterns[33319] = 29'b1_000001000100_111_1_000001000100;
      patterns[33320] = 29'b1_000001000101_000_1_000001000101;
      patterns[33321] = 29'b1_000001000101_001_1_000101000001;
      patterns[33322] = 29'b1_000001000101_010_0_000010001011;
      patterns[33323] = 29'b1_000001000101_011_0_000100010110;
      patterns[33324] = 29'b1_000001000101_100_1_100000100010;
      patterns[33325] = 29'b1_000001000101_101_0_110000010001;
      patterns[33326] = 29'b1_000001000101_110_1_000001000101;
      patterns[33327] = 29'b1_000001000101_111_1_000001000101;
      patterns[33328] = 29'b1_000001000110_000_1_000001000110;
      patterns[33329] = 29'b1_000001000110_001_1_000110000001;
      patterns[33330] = 29'b1_000001000110_010_0_000010001101;
      patterns[33331] = 29'b1_000001000110_011_0_000100011010;
      patterns[33332] = 29'b1_000001000110_100_0_100000100011;
      patterns[33333] = 29'b1_000001000110_101_1_010000010001;
      patterns[33334] = 29'b1_000001000110_110_1_000001000110;
      patterns[33335] = 29'b1_000001000110_111_1_000001000110;
      patterns[33336] = 29'b1_000001000111_000_1_000001000111;
      patterns[33337] = 29'b1_000001000111_001_1_000111000001;
      patterns[33338] = 29'b1_000001000111_010_0_000010001111;
      patterns[33339] = 29'b1_000001000111_011_0_000100011110;
      patterns[33340] = 29'b1_000001000111_100_1_100000100011;
      patterns[33341] = 29'b1_000001000111_101_1_110000010001;
      patterns[33342] = 29'b1_000001000111_110_1_000001000111;
      patterns[33343] = 29'b1_000001000111_111_1_000001000111;
      patterns[33344] = 29'b1_000001001000_000_1_000001001000;
      patterns[33345] = 29'b1_000001001000_001_1_001000000001;
      patterns[33346] = 29'b1_000001001000_010_0_000010010001;
      patterns[33347] = 29'b1_000001001000_011_0_000100100010;
      patterns[33348] = 29'b1_000001001000_100_0_100000100100;
      patterns[33349] = 29'b1_000001001000_101_0_010000010010;
      patterns[33350] = 29'b1_000001001000_110_1_000001001000;
      patterns[33351] = 29'b1_000001001000_111_1_000001001000;
      patterns[33352] = 29'b1_000001001001_000_1_000001001001;
      patterns[33353] = 29'b1_000001001001_001_1_001001000001;
      patterns[33354] = 29'b1_000001001001_010_0_000010010011;
      patterns[33355] = 29'b1_000001001001_011_0_000100100110;
      patterns[33356] = 29'b1_000001001001_100_1_100000100100;
      patterns[33357] = 29'b1_000001001001_101_0_110000010010;
      patterns[33358] = 29'b1_000001001001_110_1_000001001001;
      patterns[33359] = 29'b1_000001001001_111_1_000001001001;
      patterns[33360] = 29'b1_000001001010_000_1_000001001010;
      patterns[33361] = 29'b1_000001001010_001_1_001010000001;
      patterns[33362] = 29'b1_000001001010_010_0_000010010101;
      patterns[33363] = 29'b1_000001001010_011_0_000100101010;
      patterns[33364] = 29'b1_000001001010_100_0_100000100101;
      patterns[33365] = 29'b1_000001001010_101_1_010000010010;
      patterns[33366] = 29'b1_000001001010_110_1_000001001010;
      patterns[33367] = 29'b1_000001001010_111_1_000001001010;
      patterns[33368] = 29'b1_000001001011_000_1_000001001011;
      patterns[33369] = 29'b1_000001001011_001_1_001011000001;
      patterns[33370] = 29'b1_000001001011_010_0_000010010111;
      patterns[33371] = 29'b1_000001001011_011_0_000100101110;
      patterns[33372] = 29'b1_000001001011_100_1_100000100101;
      patterns[33373] = 29'b1_000001001011_101_1_110000010010;
      patterns[33374] = 29'b1_000001001011_110_1_000001001011;
      patterns[33375] = 29'b1_000001001011_111_1_000001001011;
      patterns[33376] = 29'b1_000001001100_000_1_000001001100;
      patterns[33377] = 29'b1_000001001100_001_1_001100000001;
      patterns[33378] = 29'b1_000001001100_010_0_000010011001;
      patterns[33379] = 29'b1_000001001100_011_0_000100110010;
      patterns[33380] = 29'b1_000001001100_100_0_100000100110;
      patterns[33381] = 29'b1_000001001100_101_0_010000010011;
      patterns[33382] = 29'b1_000001001100_110_1_000001001100;
      patterns[33383] = 29'b1_000001001100_111_1_000001001100;
      patterns[33384] = 29'b1_000001001101_000_1_000001001101;
      patterns[33385] = 29'b1_000001001101_001_1_001101000001;
      patterns[33386] = 29'b1_000001001101_010_0_000010011011;
      patterns[33387] = 29'b1_000001001101_011_0_000100110110;
      patterns[33388] = 29'b1_000001001101_100_1_100000100110;
      patterns[33389] = 29'b1_000001001101_101_0_110000010011;
      patterns[33390] = 29'b1_000001001101_110_1_000001001101;
      patterns[33391] = 29'b1_000001001101_111_1_000001001101;
      patterns[33392] = 29'b1_000001001110_000_1_000001001110;
      patterns[33393] = 29'b1_000001001110_001_1_001110000001;
      patterns[33394] = 29'b1_000001001110_010_0_000010011101;
      patterns[33395] = 29'b1_000001001110_011_0_000100111010;
      patterns[33396] = 29'b1_000001001110_100_0_100000100111;
      patterns[33397] = 29'b1_000001001110_101_1_010000010011;
      patterns[33398] = 29'b1_000001001110_110_1_000001001110;
      patterns[33399] = 29'b1_000001001110_111_1_000001001110;
      patterns[33400] = 29'b1_000001001111_000_1_000001001111;
      patterns[33401] = 29'b1_000001001111_001_1_001111000001;
      patterns[33402] = 29'b1_000001001111_010_0_000010011111;
      patterns[33403] = 29'b1_000001001111_011_0_000100111110;
      patterns[33404] = 29'b1_000001001111_100_1_100000100111;
      patterns[33405] = 29'b1_000001001111_101_1_110000010011;
      patterns[33406] = 29'b1_000001001111_110_1_000001001111;
      patterns[33407] = 29'b1_000001001111_111_1_000001001111;
      patterns[33408] = 29'b1_000001010000_000_1_000001010000;
      patterns[33409] = 29'b1_000001010000_001_1_010000000001;
      patterns[33410] = 29'b1_000001010000_010_0_000010100001;
      patterns[33411] = 29'b1_000001010000_011_0_000101000010;
      patterns[33412] = 29'b1_000001010000_100_0_100000101000;
      patterns[33413] = 29'b1_000001010000_101_0_010000010100;
      patterns[33414] = 29'b1_000001010000_110_1_000001010000;
      patterns[33415] = 29'b1_000001010000_111_1_000001010000;
      patterns[33416] = 29'b1_000001010001_000_1_000001010001;
      patterns[33417] = 29'b1_000001010001_001_1_010001000001;
      patterns[33418] = 29'b1_000001010001_010_0_000010100011;
      patterns[33419] = 29'b1_000001010001_011_0_000101000110;
      patterns[33420] = 29'b1_000001010001_100_1_100000101000;
      patterns[33421] = 29'b1_000001010001_101_0_110000010100;
      patterns[33422] = 29'b1_000001010001_110_1_000001010001;
      patterns[33423] = 29'b1_000001010001_111_1_000001010001;
      patterns[33424] = 29'b1_000001010010_000_1_000001010010;
      patterns[33425] = 29'b1_000001010010_001_1_010010000001;
      patterns[33426] = 29'b1_000001010010_010_0_000010100101;
      patterns[33427] = 29'b1_000001010010_011_0_000101001010;
      patterns[33428] = 29'b1_000001010010_100_0_100000101001;
      patterns[33429] = 29'b1_000001010010_101_1_010000010100;
      patterns[33430] = 29'b1_000001010010_110_1_000001010010;
      patterns[33431] = 29'b1_000001010010_111_1_000001010010;
      patterns[33432] = 29'b1_000001010011_000_1_000001010011;
      patterns[33433] = 29'b1_000001010011_001_1_010011000001;
      patterns[33434] = 29'b1_000001010011_010_0_000010100111;
      patterns[33435] = 29'b1_000001010011_011_0_000101001110;
      patterns[33436] = 29'b1_000001010011_100_1_100000101001;
      patterns[33437] = 29'b1_000001010011_101_1_110000010100;
      patterns[33438] = 29'b1_000001010011_110_1_000001010011;
      patterns[33439] = 29'b1_000001010011_111_1_000001010011;
      patterns[33440] = 29'b1_000001010100_000_1_000001010100;
      patterns[33441] = 29'b1_000001010100_001_1_010100000001;
      patterns[33442] = 29'b1_000001010100_010_0_000010101001;
      patterns[33443] = 29'b1_000001010100_011_0_000101010010;
      patterns[33444] = 29'b1_000001010100_100_0_100000101010;
      patterns[33445] = 29'b1_000001010100_101_0_010000010101;
      patterns[33446] = 29'b1_000001010100_110_1_000001010100;
      patterns[33447] = 29'b1_000001010100_111_1_000001010100;
      patterns[33448] = 29'b1_000001010101_000_1_000001010101;
      patterns[33449] = 29'b1_000001010101_001_1_010101000001;
      patterns[33450] = 29'b1_000001010101_010_0_000010101011;
      patterns[33451] = 29'b1_000001010101_011_0_000101010110;
      patterns[33452] = 29'b1_000001010101_100_1_100000101010;
      patterns[33453] = 29'b1_000001010101_101_0_110000010101;
      patterns[33454] = 29'b1_000001010101_110_1_000001010101;
      patterns[33455] = 29'b1_000001010101_111_1_000001010101;
      patterns[33456] = 29'b1_000001010110_000_1_000001010110;
      patterns[33457] = 29'b1_000001010110_001_1_010110000001;
      patterns[33458] = 29'b1_000001010110_010_0_000010101101;
      patterns[33459] = 29'b1_000001010110_011_0_000101011010;
      patterns[33460] = 29'b1_000001010110_100_0_100000101011;
      patterns[33461] = 29'b1_000001010110_101_1_010000010101;
      patterns[33462] = 29'b1_000001010110_110_1_000001010110;
      patterns[33463] = 29'b1_000001010110_111_1_000001010110;
      patterns[33464] = 29'b1_000001010111_000_1_000001010111;
      patterns[33465] = 29'b1_000001010111_001_1_010111000001;
      patterns[33466] = 29'b1_000001010111_010_0_000010101111;
      patterns[33467] = 29'b1_000001010111_011_0_000101011110;
      patterns[33468] = 29'b1_000001010111_100_1_100000101011;
      patterns[33469] = 29'b1_000001010111_101_1_110000010101;
      patterns[33470] = 29'b1_000001010111_110_1_000001010111;
      patterns[33471] = 29'b1_000001010111_111_1_000001010111;
      patterns[33472] = 29'b1_000001011000_000_1_000001011000;
      patterns[33473] = 29'b1_000001011000_001_1_011000000001;
      patterns[33474] = 29'b1_000001011000_010_0_000010110001;
      patterns[33475] = 29'b1_000001011000_011_0_000101100010;
      patterns[33476] = 29'b1_000001011000_100_0_100000101100;
      patterns[33477] = 29'b1_000001011000_101_0_010000010110;
      patterns[33478] = 29'b1_000001011000_110_1_000001011000;
      patterns[33479] = 29'b1_000001011000_111_1_000001011000;
      patterns[33480] = 29'b1_000001011001_000_1_000001011001;
      patterns[33481] = 29'b1_000001011001_001_1_011001000001;
      patterns[33482] = 29'b1_000001011001_010_0_000010110011;
      patterns[33483] = 29'b1_000001011001_011_0_000101100110;
      patterns[33484] = 29'b1_000001011001_100_1_100000101100;
      patterns[33485] = 29'b1_000001011001_101_0_110000010110;
      patterns[33486] = 29'b1_000001011001_110_1_000001011001;
      patterns[33487] = 29'b1_000001011001_111_1_000001011001;
      patterns[33488] = 29'b1_000001011010_000_1_000001011010;
      patterns[33489] = 29'b1_000001011010_001_1_011010000001;
      patterns[33490] = 29'b1_000001011010_010_0_000010110101;
      patterns[33491] = 29'b1_000001011010_011_0_000101101010;
      patterns[33492] = 29'b1_000001011010_100_0_100000101101;
      patterns[33493] = 29'b1_000001011010_101_1_010000010110;
      patterns[33494] = 29'b1_000001011010_110_1_000001011010;
      patterns[33495] = 29'b1_000001011010_111_1_000001011010;
      patterns[33496] = 29'b1_000001011011_000_1_000001011011;
      patterns[33497] = 29'b1_000001011011_001_1_011011000001;
      patterns[33498] = 29'b1_000001011011_010_0_000010110111;
      patterns[33499] = 29'b1_000001011011_011_0_000101101110;
      patterns[33500] = 29'b1_000001011011_100_1_100000101101;
      patterns[33501] = 29'b1_000001011011_101_1_110000010110;
      patterns[33502] = 29'b1_000001011011_110_1_000001011011;
      patterns[33503] = 29'b1_000001011011_111_1_000001011011;
      patterns[33504] = 29'b1_000001011100_000_1_000001011100;
      patterns[33505] = 29'b1_000001011100_001_1_011100000001;
      patterns[33506] = 29'b1_000001011100_010_0_000010111001;
      patterns[33507] = 29'b1_000001011100_011_0_000101110010;
      patterns[33508] = 29'b1_000001011100_100_0_100000101110;
      patterns[33509] = 29'b1_000001011100_101_0_010000010111;
      patterns[33510] = 29'b1_000001011100_110_1_000001011100;
      patterns[33511] = 29'b1_000001011100_111_1_000001011100;
      patterns[33512] = 29'b1_000001011101_000_1_000001011101;
      patterns[33513] = 29'b1_000001011101_001_1_011101000001;
      patterns[33514] = 29'b1_000001011101_010_0_000010111011;
      patterns[33515] = 29'b1_000001011101_011_0_000101110110;
      patterns[33516] = 29'b1_000001011101_100_1_100000101110;
      patterns[33517] = 29'b1_000001011101_101_0_110000010111;
      patterns[33518] = 29'b1_000001011101_110_1_000001011101;
      patterns[33519] = 29'b1_000001011101_111_1_000001011101;
      patterns[33520] = 29'b1_000001011110_000_1_000001011110;
      patterns[33521] = 29'b1_000001011110_001_1_011110000001;
      patterns[33522] = 29'b1_000001011110_010_0_000010111101;
      patterns[33523] = 29'b1_000001011110_011_0_000101111010;
      patterns[33524] = 29'b1_000001011110_100_0_100000101111;
      patterns[33525] = 29'b1_000001011110_101_1_010000010111;
      patterns[33526] = 29'b1_000001011110_110_1_000001011110;
      patterns[33527] = 29'b1_000001011110_111_1_000001011110;
      patterns[33528] = 29'b1_000001011111_000_1_000001011111;
      patterns[33529] = 29'b1_000001011111_001_1_011111000001;
      patterns[33530] = 29'b1_000001011111_010_0_000010111111;
      patterns[33531] = 29'b1_000001011111_011_0_000101111110;
      patterns[33532] = 29'b1_000001011111_100_1_100000101111;
      patterns[33533] = 29'b1_000001011111_101_1_110000010111;
      patterns[33534] = 29'b1_000001011111_110_1_000001011111;
      patterns[33535] = 29'b1_000001011111_111_1_000001011111;
      patterns[33536] = 29'b1_000001100000_000_1_000001100000;
      patterns[33537] = 29'b1_000001100000_001_1_100000000001;
      patterns[33538] = 29'b1_000001100000_010_0_000011000001;
      patterns[33539] = 29'b1_000001100000_011_0_000110000010;
      patterns[33540] = 29'b1_000001100000_100_0_100000110000;
      patterns[33541] = 29'b1_000001100000_101_0_010000011000;
      patterns[33542] = 29'b1_000001100000_110_1_000001100000;
      patterns[33543] = 29'b1_000001100000_111_1_000001100000;
      patterns[33544] = 29'b1_000001100001_000_1_000001100001;
      patterns[33545] = 29'b1_000001100001_001_1_100001000001;
      patterns[33546] = 29'b1_000001100001_010_0_000011000011;
      patterns[33547] = 29'b1_000001100001_011_0_000110000110;
      patterns[33548] = 29'b1_000001100001_100_1_100000110000;
      patterns[33549] = 29'b1_000001100001_101_0_110000011000;
      patterns[33550] = 29'b1_000001100001_110_1_000001100001;
      patterns[33551] = 29'b1_000001100001_111_1_000001100001;
      patterns[33552] = 29'b1_000001100010_000_1_000001100010;
      patterns[33553] = 29'b1_000001100010_001_1_100010000001;
      patterns[33554] = 29'b1_000001100010_010_0_000011000101;
      patterns[33555] = 29'b1_000001100010_011_0_000110001010;
      patterns[33556] = 29'b1_000001100010_100_0_100000110001;
      patterns[33557] = 29'b1_000001100010_101_1_010000011000;
      patterns[33558] = 29'b1_000001100010_110_1_000001100010;
      patterns[33559] = 29'b1_000001100010_111_1_000001100010;
      patterns[33560] = 29'b1_000001100011_000_1_000001100011;
      patterns[33561] = 29'b1_000001100011_001_1_100011000001;
      patterns[33562] = 29'b1_000001100011_010_0_000011000111;
      patterns[33563] = 29'b1_000001100011_011_0_000110001110;
      patterns[33564] = 29'b1_000001100011_100_1_100000110001;
      patterns[33565] = 29'b1_000001100011_101_1_110000011000;
      patterns[33566] = 29'b1_000001100011_110_1_000001100011;
      patterns[33567] = 29'b1_000001100011_111_1_000001100011;
      patterns[33568] = 29'b1_000001100100_000_1_000001100100;
      patterns[33569] = 29'b1_000001100100_001_1_100100000001;
      patterns[33570] = 29'b1_000001100100_010_0_000011001001;
      patterns[33571] = 29'b1_000001100100_011_0_000110010010;
      patterns[33572] = 29'b1_000001100100_100_0_100000110010;
      patterns[33573] = 29'b1_000001100100_101_0_010000011001;
      patterns[33574] = 29'b1_000001100100_110_1_000001100100;
      patterns[33575] = 29'b1_000001100100_111_1_000001100100;
      patterns[33576] = 29'b1_000001100101_000_1_000001100101;
      patterns[33577] = 29'b1_000001100101_001_1_100101000001;
      patterns[33578] = 29'b1_000001100101_010_0_000011001011;
      patterns[33579] = 29'b1_000001100101_011_0_000110010110;
      patterns[33580] = 29'b1_000001100101_100_1_100000110010;
      patterns[33581] = 29'b1_000001100101_101_0_110000011001;
      patterns[33582] = 29'b1_000001100101_110_1_000001100101;
      patterns[33583] = 29'b1_000001100101_111_1_000001100101;
      patterns[33584] = 29'b1_000001100110_000_1_000001100110;
      patterns[33585] = 29'b1_000001100110_001_1_100110000001;
      patterns[33586] = 29'b1_000001100110_010_0_000011001101;
      patterns[33587] = 29'b1_000001100110_011_0_000110011010;
      patterns[33588] = 29'b1_000001100110_100_0_100000110011;
      patterns[33589] = 29'b1_000001100110_101_1_010000011001;
      patterns[33590] = 29'b1_000001100110_110_1_000001100110;
      patterns[33591] = 29'b1_000001100110_111_1_000001100110;
      patterns[33592] = 29'b1_000001100111_000_1_000001100111;
      patterns[33593] = 29'b1_000001100111_001_1_100111000001;
      patterns[33594] = 29'b1_000001100111_010_0_000011001111;
      patterns[33595] = 29'b1_000001100111_011_0_000110011110;
      patterns[33596] = 29'b1_000001100111_100_1_100000110011;
      patterns[33597] = 29'b1_000001100111_101_1_110000011001;
      patterns[33598] = 29'b1_000001100111_110_1_000001100111;
      patterns[33599] = 29'b1_000001100111_111_1_000001100111;
      patterns[33600] = 29'b1_000001101000_000_1_000001101000;
      patterns[33601] = 29'b1_000001101000_001_1_101000000001;
      patterns[33602] = 29'b1_000001101000_010_0_000011010001;
      patterns[33603] = 29'b1_000001101000_011_0_000110100010;
      patterns[33604] = 29'b1_000001101000_100_0_100000110100;
      patterns[33605] = 29'b1_000001101000_101_0_010000011010;
      patterns[33606] = 29'b1_000001101000_110_1_000001101000;
      patterns[33607] = 29'b1_000001101000_111_1_000001101000;
      patterns[33608] = 29'b1_000001101001_000_1_000001101001;
      patterns[33609] = 29'b1_000001101001_001_1_101001000001;
      patterns[33610] = 29'b1_000001101001_010_0_000011010011;
      patterns[33611] = 29'b1_000001101001_011_0_000110100110;
      patterns[33612] = 29'b1_000001101001_100_1_100000110100;
      patterns[33613] = 29'b1_000001101001_101_0_110000011010;
      patterns[33614] = 29'b1_000001101001_110_1_000001101001;
      patterns[33615] = 29'b1_000001101001_111_1_000001101001;
      patterns[33616] = 29'b1_000001101010_000_1_000001101010;
      patterns[33617] = 29'b1_000001101010_001_1_101010000001;
      patterns[33618] = 29'b1_000001101010_010_0_000011010101;
      patterns[33619] = 29'b1_000001101010_011_0_000110101010;
      patterns[33620] = 29'b1_000001101010_100_0_100000110101;
      patterns[33621] = 29'b1_000001101010_101_1_010000011010;
      patterns[33622] = 29'b1_000001101010_110_1_000001101010;
      patterns[33623] = 29'b1_000001101010_111_1_000001101010;
      patterns[33624] = 29'b1_000001101011_000_1_000001101011;
      patterns[33625] = 29'b1_000001101011_001_1_101011000001;
      patterns[33626] = 29'b1_000001101011_010_0_000011010111;
      patterns[33627] = 29'b1_000001101011_011_0_000110101110;
      patterns[33628] = 29'b1_000001101011_100_1_100000110101;
      patterns[33629] = 29'b1_000001101011_101_1_110000011010;
      patterns[33630] = 29'b1_000001101011_110_1_000001101011;
      patterns[33631] = 29'b1_000001101011_111_1_000001101011;
      patterns[33632] = 29'b1_000001101100_000_1_000001101100;
      patterns[33633] = 29'b1_000001101100_001_1_101100000001;
      patterns[33634] = 29'b1_000001101100_010_0_000011011001;
      patterns[33635] = 29'b1_000001101100_011_0_000110110010;
      patterns[33636] = 29'b1_000001101100_100_0_100000110110;
      patterns[33637] = 29'b1_000001101100_101_0_010000011011;
      patterns[33638] = 29'b1_000001101100_110_1_000001101100;
      patterns[33639] = 29'b1_000001101100_111_1_000001101100;
      patterns[33640] = 29'b1_000001101101_000_1_000001101101;
      patterns[33641] = 29'b1_000001101101_001_1_101101000001;
      patterns[33642] = 29'b1_000001101101_010_0_000011011011;
      patterns[33643] = 29'b1_000001101101_011_0_000110110110;
      patterns[33644] = 29'b1_000001101101_100_1_100000110110;
      patterns[33645] = 29'b1_000001101101_101_0_110000011011;
      patterns[33646] = 29'b1_000001101101_110_1_000001101101;
      patterns[33647] = 29'b1_000001101101_111_1_000001101101;
      patterns[33648] = 29'b1_000001101110_000_1_000001101110;
      patterns[33649] = 29'b1_000001101110_001_1_101110000001;
      patterns[33650] = 29'b1_000001101110_010_0_000011011101;
      patterns[33651] = 29'b1_000001101110_011_0_000110111010;
      patterns[33652] = 29'b1_000001101110_100_0_100000110111;
      patterns[33653] = 29'b1_000001101110_101_1_010000011011;
      patterns[33654] = 29'b1_000001101110_110_1_000001101110;
      patterns[33655] = 29'b1_000001101110_111_1_000001101110;
      patterns[33656] = 29'b1_000001101111_000_1_000001101111;
      patterns[33657] = 29'b1_000001101111_001_1_101111000001;
      patterns[33658] = 29'b1_000001101111_010_0_000011011111;
      patterns[33659] = 29'b1_000001101111_011_0_000110111110;
      patterns[33660] = 29'b1_000001101111_100_1_100000110111;
      patterns[33661] = 29'b1_000001101111_101_1_110000011011;
      patterns[33662] = 29'b1_000001101111_110_1_000001101111;
      patterns[33663] = 29'b1_000001101111_111_1_000001101111;
      patterns[33664] = 29'b1_000001110000_000_1_000001110000;
      patterns[33665] = 29'b1_000001110000_001_1_110000000001;
      patterns[33666] = 29'b1_000001110000_010_0_000011100001;
      patterns[33667] = 29'b1_000001110000_011_0_000111000010;
      patterns[33668] = 29'b1_000001110000_100_0_100000111000;
      patterns[33669] = 29'b1_000001110000_101_0_010000011100;
      patterns[33670] = 29'b1_000001110000_110_1_000001110000;
      patterns[33671] = 29'b1_000001110000_111_1_000001110000;
      patterns[33672] = 29'b1_000001110001_000_1_000001110001;
      patterns[33673] = 29'b1_000001110001_001_1_110001000001;
      patterns[33674] = 29'b1_000001110001_010_0_000011100011;
      patterns[33675] = 29'b1_000001110001_011_0_000111000110;
      patterns[33676] = 29'b1_000001110001_100_1_100000111000;
      patterns[33677] = 29'b1_000001110001_101_0_110000011100;
      patterns[33678] = 29'b1_000001110001_110_1_000001110001;
      patterns[33679] = 29'b1_000001110001_111_1_000001110001;
      patterns[33680] = 29'b1_000001110010_000_1_000001110010;
      patterns[33681] = 29'b1_000001110010_001_1_110010000001;
      patterns[33682] = 29'b1_000001110010_010_0_000011100101;
      patterns[33683] = 29'b1_000001110010_011_0_000111001010;
      patterns[33684] = 29'b1_000001110010_100_0_100000111001;
      patterns[33685] = 29'b1_000001110010_101_1_010000011100;
      patterns[33686] = 29'b1_000001110010_110_1_000001110010;
      patterns[33687] = 29'b1_000001110010_111_1_000001110010;
      patterns[33688] = 29'b1_000001110011_000_1_000001110011;
      patterns[33689] = 29'b1_000001110011_001_1_110011000001;
      patterns[33690] = 29'b1_000001110011_010_0_000011100111;
      patterns[33691] = 29'b1_000001110011_011_0_000111001110;
      patterns[33692] = 29'b1_000001110011_100_1_100000111001;
      patterns[33693] = 29'b1_000001110011_101_1_110000011100;
      patterns[33694] = 29'b1_000001110011_110_1_000001110011;
      patterns[33695] = 29'b1_000001110011_111_1_000001110011;
      patterns[33696] = 29'b1_000001110100_000_1_000001110100;
      patterns[33697] = 29'b1_000001110100_001_1_110100000001;
      patterns[33698] = 29'b1_000001110100_010_0_000011101001;
      patterns[33699] = 29'b1_000001110100_011_0_000111010010;
      patterns[33700] = 29'b1_000001110100_100_0_100000111010;
      patterns[33701] = 29'b1_000001110100_101_0_010000011101;
      patterns[33702] = 29'b1_000001110100_110_1_000001110100;
      patterns[33703] = 29'b1_000001110100_111_1_000001110100;
      patterns[33704] = 29'b1_000001110101_000_1_000001110101;
      patterns[33705] = 29'b1_000001110101_001_1_110101000001;
      patterns[33706] = 29'b1_000001110101_010_0_000011101011;
      patterns[33707] = 29'b1_000001110101_011_0_000111010110;
      patterns[33708] = 29'b1_000001110101_100_1_100000111010;
      patterns[33709] = 29'b1_000001110101_101_0_110000011101;
      patterns[33710] = 29'b1_000001110101_110_1_000001110101;
      patterns[33711] = 29'b1_000001110101_111_1_000001110101;
      patterns[33712] = 29'b1_000001110110_000_1_000001110110;
      patterns[33713] = 29'b1_000001110110_001_1_110110000001;
      patterns[33714] = 29'b1_000001110110_010_0_000011101101;
      patterns[33715] = 29'b1_000001110110_011_0_000111011010;
      patterns[33716] = 29'b1_000001110110_100_0_100000111011;
      patterns[33717] = 29'b1_000001110110_101_1_010000011101;
      patterns[33718] = 29'b1_000001110110_110_1_000001110110;
      patterns[33719] = 29'b1_000001110110_111_1_000001110110;
      patterns[33720] = 29'b1_000001110111_000_1_000001110111;
      patterns[33721] = 29'b1_000001110111_001_1_110111000001;
      patterns[33722] = 29'b1_000001110111_010_0_000011101111;
      patterns[33723] = 29'b1_000001110111_011_0_000111011110;
      patterns[33724] = 29'b1_000001110111_100_1_100000111011;
      patterns[33725] = 29'b1_000001110111_101_1_110000011101;
      patterns[33726] = 29'b1_000001110111_110_1_000001110111;
      patterns[33727] = 29'b1_000001110111_111_1_000001110111;
      patterns[33728] = 29'b1_000001111000_000_1_000001111000;
      patterns[33729] = 29'b1_000001111000_001_1_111000000001;
      patterns[33730] = 29'b1_000001111000_010_0_000011110001;
      patterns[33731] = 29'b1_000001111000_011_0_000111100010;
      patterns[33732] = 29'b1_000001111000_100_0_100000111100;
      patterns[33733] = 29'b1_000001111000_101_0_010000011110;
      patterns[33734] = 29'b1_000001111000_110_1_000001111000;
      patterns[33735] = 29'b1_000001111000_111_1_000001111000;
      patterns[33736] = 29'b1_000001111001_000_1_000001111001;
      patterns[33737] = 29'b1_000001111001_001_1_111001000001;
      patterns[33738] = 29'b1_000001111001_010_0_000011110011;
      patterns[33739] = 29'b1_000001111001_011_0_000111100110;
      patterns[33740] = 29'b1_000001111001_100_1_100000111100;
      patterns[33741] = 29'b1_000001111001_101_0_110000011110;
      patterns[33742] = 29'b1_000001111001_110_1_000001111001;
      patterns[33743] = 29'b1_000001111001_111_1_000001111001;
      patterns[33744] = 29'b1_000001111010_000_1_000001111010;
      patterns[33745] = 29'b1_000001111010_001_1_111010000001;
      patterns[33746] = 29'b1_000001111010_010_0_000011110101;
      patterns[33747] = 29'b1_000001111010_011_0_000111101010;
      patterns[33748] = 29'b1_000001111010_100_0_100000111101;
      patterns[33749] = 29'b1_000001111010_101_1_010000011110;
      patterns[33750] = 29'b1_000001111010_110_1_000001111010;
      patterns[33751] = 29'b1_000001111010_111_1_000001111010;
      patterns[33752] = 29'b1_000001111011_000_1_000001111011;
      patterns[33753] = 29'b1_000001111011_001_1_111011000001;
      patterns[33754] = 29'b1_000001111011_010_0_000011110111;
      patterns[33755] = 29'b1_000001111011_011_0_000111101110;
      patterns[33756] = 29'b1_000001111011_100_1_100000111101;
      patterns[33757] = 29'b1_000001111011_101_1_110000011110;
      patterns[33758] = 29'b1_000001111011_110_1_000001111011;
      patterns[33759] = 29'b1_000001111011_111_1_000001111011;
      patterns[33760] = 29'b1_000001111100_000_1_000001111100;
      patterns[33761] = 29'b1_000001111100_001_1_111100000001;
      patterns[33762] = 29'b1_000001111100_010_0_000011111001;
      patterns[33763] = 29'b1_000001111100_011_0_000111110010;
      patterns[33764] = 29'b1_000001111100_100_0_100000111110;
      patterns[33765] = 29'b1_000001111100_101_0_010000011111;
      patterns[33766] = 29'b1_000001111100_110_1_000001111100;
      patterns[33767] = 29'b1_000001111100_111_1_000001111100;
      patterns[33768] = 29'b1_000001111101_000_1_000001111101;
      patterns[33769] = 29'b1_000001111101_001_1_111101000001;
      patterns[33770] = 29'b1_000001111101_010_0_000011111011;
      patterns[33771] = 29'b1_000001111101_011_0_000111110110;
      patterns[33772] = 29'b1_000001111101_100_1_100000111110;
      patterns[33773] = 29'b1_000001111101_101_0_110000011111;
      patterns[33774] = 29'b1_000001111101_110_1_000001111101;
      patterns[33775] = 29'b1_000001111101_111_1_000001111101;
      patterns[33776] = 29'b1_000001111110_000_1_000001111110;
      patterns[33777] = 29'b1_000001111110_001_1_111110000001;
      patterns[33778] = 29'b1_000001111110_010_0_000011111101;
      patterns[33779] = 29'b1_000001111110_011_0_000111111010;
      patterns[33780] = 29'b1_000001111110_100_0_100000111111;
      patterns[33781] = 29'b1_000001111110_101_1_010000011111;
      patterns[33782] = 29'b1_000001111110_110_1_000001111110;
      patterns[33783] = 29'b1_000001111110_111_1_000001111110;
      patterns[33784] = 29'b1_000001111111_000_1_000001111111;
      patterns[33785] = 29'b1_000001111111_001_1_111111000001;
      patterns[33786] = 29'b1_000001111111_010_0_000011111111;
      patterns[33787] = 29'b1_000001111111_011_0_000111111110;
      patterns[33788] = 29'b1_000001111111_100_1_100000111111;
      patterns[33789] = 29'b1_000001111111_101_1_110000011111;
      patterns[33790] = 29'b1_000001111111_110_1_000001111111;
      patterns[33791] = 29'b1_000001111111_111_1_000001111111;
      patterns[33792] = 29'b1_000010000000_000_1_000010000000;
      patterns[33793] = 29'b1_000010000000_001_1_000000000010;
      patterns[33794] = 29'b1_000010000000_010_0_000100000001;
      patterns[33795] = 29'b1_000010000000_011_0_001000000010;
      patterns[33796] = 29'b1_000010000000_100_0_100001000000;
      patterns[33797] = 29'b1_000010000000_101_0_010000100000;
      patterns[33798] = 29'b1_000010000000_110_1_000010000000;
      patterns[33799] = 29'b1_000010000000_111_1_000010000000;
      patterns[33800] = 29'b1_000010000001_000_1_000010000001;
      patterns[33801] = 29'b1_000010000001_001_1_000001000010;
      patterns[33802] = 29'b1_000010000001_010_0_000100000011;
      patterns[33803] = 29'b1_000010000001_011_0_001000000110;
      patterns[33804] = 29'b1_000010000001_100_1_100001000000;
      patterns[33805] = 29'b1_000010000001_101_0_110000100000;
      patterns[33806] = 29'b1_000010000001_110_1_000010000001;
      patterns[33807] = 29'b1_000010000001_111_1_000010000001;
      patterns[33808] = 29'b1_000010000010_000_1_000010000010;
      patterns[33809] = 29'b1_000010000010_001_1_000010000010;
      patterns[33810] = 29'b1_000010000010_010_0_000100000101;
      patterns[33811] = 29'b1_000010000010_011_0_001000001010;
      patterns[33812] = 29'b1_000010000010_100_0_100001000001;
      patterns[33813] = 29'b1_000010000010_101_1_010000100000;
      patterns[33814] = 29'b1_000010000010_110_1_000010000010;
      patterns[33815] = 29'b1_000010000010_111_1_000010000010;
      patterns[33816] = 29'b1_000010000011_000_1_000010000011;
      patterns[33817] = 29'b1_000010000011_001_1_000011000010;
      patterns[33818] = 29'b1_000010000011_010_0_000100000111;
      patterns[33819] = 29'b1_000010000011_011_0_001000001110;
      patterns[33820] = 29'b1_000010000011_100_1_100001000001;
      patterns[33821] = 29'b1_000010000011_101_1_110000100000;
      patterns[33822] = 29'b1_000010000011_110_1_000010000011;
      patterns[33823] = 29'b1_000010000011_111_1_000010000011;
      patterns[33824] = 29'b1_000010000100_000_1_000010000100;
      patterns[33825] = 29'b1_000010000100_001_1_000100000010;
      patterns[33826] = 29'b1_000010000100_010_0_000100001001;
      patterns[33827] = 29'b1_000010000100_011_0_001000010010;
      patterns[33828] = 29'b1_000010000100_100_0_100001000010;
      patterns[33829] = 29'b1_000010000100_101_0_010000100001;
      patterns[33830] = 29'b1_000010000100_110_1_000010000100;
      patterns[33831] = 29'b1_000010000100_111_1_000010000100;
      patterns[33832] = 29'b1_000010000101_000_1_000010000101;
      patterns[33833] = 29'b1_000010000101_001_1_000101000010;
      patterns[33834] = 29'b1_000010000101_010_0_000100001011;
      patterns[33835] = 29'b1_000010000101_011_0_001000010110;
      patterns[33836] = 29'b1_000010000101_100_1_100001000010;
      patterns[33837] = 29'b1_000010000101_101_0_110000100001;
      patterns[33838] = 29'b1_000010000101_110_1_000010000101;
      patterns[33839] = 29'b1_000010000101_111_1_000010000101;
      patterns[33840] = 29'b1_000010000110_000_1_000010000110;
      patterns[33841] = 29'b1_000010000110_001_1_000110000010;
      patterns[33842] = 29'b1_000010000110_010_0_000100001101;
      patterns[33843] = 29'b1_000010000110_011_0_001000011010;
      patterns[33844] = 29'b1_000010000110_100_0_100001000011;
      patterns[33845] = 29'b1_000010000110_101_1_010000100001;
      patterns[33846] = 29'b1_000010000110_110_1_000010000110;
      patterns[33847] = 29'b1_000010000110_111_1_000010000110;
      patterns[33848] = 29'b1_000010000111_000_1_000010000111;
      patterns[33849] = 29'b1_000010000111_001_1_000111000010;
      patterns[33850] = 29'b1_000010000111_010_0_000100001111;
      patterns[33851] = 29'b1_000010000111_011_0_001000011110;
      patterns[33852] = 29'b1_000010000111_100_1_100001000011;
      patterns[33853] = 29'b1_000010000111_101_1_110000100001;
      patterns[33854] = 29'b1_000010000111_110_1_000010000111;
      patterns[33855] = 29'b1_000010000111_111_1_000010000111;
      patterns[33856] = 29'b1_000010001000_000_1_000010001000;
      patterns[33857] = 29'b1_000010001000_001_1_001000000010;
      patterns[33858] = 29'b1_000010001000_010_0_000100010001;
      patterns[33859] = 29'b1_000010001000_011_0_001000100010;
      patterns[33860] = 29'b1_000010001000_100_0_100001000100;
      patterns[33861] = 29'b1_000010001000_101_0_010000100010;
      patterns[33862] = 29'b1_000010001000_110_1_000010001000;
      patterns[33863] = 29'b1_000010001000_111_1_000010001000;
      patterns[33864] = 29'b1_000010001001_000_1_000010001001;
      patterns[33865] = 29'b1_000010001001_001_1_001001000010;
      patterns[33866] = 29'b1_000010001001_010_0_000100010011;
      patterns[33867] = 29'b1_000010001001_011_0_001000100110;
      patterns[33868] = 29'b1_000010001001_100_1_100001000100;
      patterns[33869] = 29'b1_000010001001_101_0_110000100010;
      patterns[33870] = 29'b1_000010001001_110_1_000010001001;
      patterns[33871] = 29'b1_000010001001_111_1_000010001001;
      patterns[33872] = 29'b1_000010001010_000_1_000010001010;
      patterns[33873] = 29'b1_000010001010_001_1_001010000010;
      patterns[33874] = 29'b1_000010001010_010_0_000100010101;
      patterns[33875] = 29'b1_000010001010_011_0_001000101010;
      patterns[33876] = 29'b1_000010001010_100_0_100001000101;
      patterns[33877] = 29'b1_000010001010_101_1_010000100010;
      patterns[33878] = 29'b1_000010001010_110_1_000010001010;
      patterns[33879] = 29'b1_000010001010_111_1_000010001010;
      patterns[33880] = 29'b1_000010001011_000_1_000010001011;
      patterns[33881] = 29'b1_000010001011_001_1_001011000010;
      patterns[33882] = 29'b1_000010001011_010_0_000100010111;
      patterns[33883] = 29'b1_000010001011_011_0_001000101110;
      patterns[33884] = 29'b1_000010001011_100_1_100001000101;
      patterns[33885] = 29'b1_000010001011_101_1_110000100010;
      patterns[33886] = 29'b1_000010001011_110_1_000010001011;
      patterns[33887] = 29'b1_000010001011_111_1_000010001011;
      patterns[33888] = 29'b1_000010001100_000_1_000010001100;
      patterns[33889] = 29'b1_000010001100_001_1_001100000010;
      patterns[33890] = 29'b1_000010001100_010_0_000100011001;
      patterns[33891] = 29'b1_000010001100_011_0_001000110010;
      patterns[33892] = 29'b1_000010001100_100_0_100001000110;
      patterns[33893] = 29'b1_000010001100_101_0_010000100011;
      patterns[33894] = 29'b1_000010001100_110_1_000010001100;
      patterns[33895] = 29'b1_000010001100_111_1_000010001100;
      patterns[33896] = 29'b1_000010001101_000_1_000010001101;
      patterns[33897] = 29'b1_000010001101_001_1_001101000010;
      patterns[33898] = 29'b1_000010001101_010_0_000100011011;
      patterns[33899] = 29'b1_000010001101_011_0_001000110110;
      patterns[33900] = 29'b1_000010001101_100_1_100001000110;
      patterns[33901] = 29'b1_000010001101_101_0_110000100011;
      patterns[33902] = 29'b1_000010001101_110_1_000010001101;
      patterns[33903] = 29'b1_000010001101_111_1_000010001101;
      patterns[33904] = 29'b1_000010001110_000_1_000010001110;
      patterns[33905] = 29'b1_000010001110_001_1_001110000010;
      patterns[33906] = 29'b1_000010001110_010_0_000100011101;
      patterns[33907] = 29'b1_000010001110_011_0_001000111010;
      patterns[33908] = 29'b1_000010001110_100_0_100001000111;
      patterns[33909] = 29'b1_000010001110_101_1_010000100011;
      patterns[33910] = 29'b1_000010001110_110_1_000010001110;
      patterns[33911] = 29'b1_000010001110_111_1_000010001110;
      patterns[33912] = 29'b1_000010001111_000_1_000010001111;
      patterns[33913] = 29'b1_000010001111_001_1_001111000010;
      patterns[33914] = 29'b1_000010001111_010_0_000100011111;
      patterns[33915] = 29'b1_000010001111_011_0_001000111110;
      patterns[33916] = 29'b1_000010001111_100_1_100001000111;
      patterns[33917] = 29'b1_000010001111_101_1_110000100011;
      patterns[33918] = 29'b1_000010001111_110_1_000010001111;
      patterns[33919] = 29'b1_000010001111_111_1_000010001111;
      patterns[33920] = 29'b1_000010010000_000_1_000010010000;
      patterns[33921] = 29'b1_000010010000_001_1_010000000010;
      patterns[33922] = 29'b1_000010010000_010_0_000100100001;
      patterns[33923] = 29'b1_000010010000_011_0_001001000010;
      patterns[33924] = 29'b1_000010010000_100_0_100001001000;
      patterns[33925] = 29'b1_000010010000_101_0_010000100100;
      patterns[33926] = 29'b1_000010010000_110_1_000010010000;
      patterns[33927] = 29'b1_000010010000_111_1_000010010000;
      patterns[33928] = 29'b1_000010010001_000_1_000010010001;
      patterns[33929] = 29'b1_000010010001_001_1_010001000010;
      patterns[33930] = 29'b1_000010010001_010_0_000100100011;
      patterns[33931] = 29'b1_000010010001_011_0_001001000110;
      patterns[33932] = 29'b1_000010010001_100_1_100001001000;
      patterns[33933] = 29'b1_000010010001_101_0_110000100100;
      patterns[33934] = 29'b1_000010010001_110_1_000010010001;
      patterns[33935] = 29'b1_000010010001_111_1_000010010001;
      patterns[33936] = 29'b1_000010010010_000_1_000010010010;
      patterns[33937] = 29'b1_000010010010_001_1_010010000010;
      patterns[33938] = 29'b1_000010010010_010_0_000100100101;
      patterns[33939] = 29'b1_000010010010_011_0_001001001010;
      patterns[33940] = 29'b1_000010010010_100_0_100001001001;
      patterns[33941] = 29'b1_000010010010_101_1_010000100100;
      patterns[33942] = 29'b1_000010010010_110_1_000010010010;
      patterns[33943] = 29'b1_000010010010_111_1_000010010010;
      patterns[33944] = 29'b1_000010010011_000_1_000010010011;
      patterns[33945] = 29'b1_000010010011_001_1_010011000010;
      patterns[33946] = 29'b1_000010010011_010_0_000100100111;
      patterns[33947] = 29'b1_000010010011_011_0_001001001110;
      patterns[33948] = 29'b1_000010010011_100_1_100001001001;
      patterns[33949] = 29'b1_000010010011_101_1_110000100100;
      patterns[33950] = 29'b1_000010010011_110_1_000010010011;
      patterns[33951] = 29'b1_000010010011_111_1_000010010011;
      patterns[33952] = 29'b1_000010010100_000_1_000010010100;
      patterns[33953] = 29'b1_000010010100_001_1_010100000010;
      patterns[33954] = 29'b1_000010010100_010_0_000100101001;
      patterns[33955] = 29'b1_000010010100_011_0_001001010010;
      patterns[33956] = 29'b1_000010010100_100_0_100001001010;
      patterns[33957] = 29'b1_000010010100_101_0_010000100101;
      patterns[33958] = 29'b1_000010010100_110_1_000010010100;
      patterns[33959] = 29'b1_000010010100_111_1_000010010100;
      patterns[33960] = 29'b1_000010010101_000_1_000010010101;
      patterns[33961] = 29'b1_000010010101_001_1_010101000010;
      patterns[33962] = 29'b1_000010010101_010_0_000100101011;
      patterns[33963] = 29'b1_000010010101_011_0_001001010110;
      patterns[33964] = 29'b1_000010010101_100_1_100001001010;
      patterns[33965] = 29'b1_000010010101_101_0_110000100101;
      patterns[33966] = 29'b1_000010010101_110_1_000010010101;
      patterns[33967] = 29'b1_000010010101_111_1_000010010101;
      patterns[33968] = 29'b1_000010010110_000_1_000010010110;
      patterns[33969] = 29'b1_000010010110_001_1_010110000010;
      patterns[33970] = 29'b1_000010010110_010_0_000100101101;
      patterns[33971] = 29'b1_000010010110_011_0_001001011010;
      patterns[33972] = 29'b1_000010010110_100_0_100001001011;
      patterns[33973] = 29'b1_000010010110_101_1_010000100101;
      patterns[33974] = 29'b1_000010010110_110_1_000010010110;
      patterns[33975] = 29'b1_000010010110_111_1_000010010110;
      patterns[33976] = 29'b1_000010010111_000_1_000010010111;
      patterns[33977] = 29'b1_000010010111_001_1_010111000010;
      patterns[33978] = 29'b1_000010010111_010_0_000100101111;
      patterns[33979] = 29'b1_000010010111_011_0_001001011110;
      patterns[33980] = 29'b1_000010010111_100_1_100001001011;
      patterns[33981] = 29'b1_000010010111_101_1_110000100101;
      patterns[33982] = 29'b1_000010010111_110_1_000010010111;
      patterns[33983] = 29'b1_000010010111_111_1_000010010111;
      patterns[33984] = 29'b1_000010011000_000_1_000010011000;
      patterns[33985] = 29'b1_000010011000_001_1_011000000010;
      patterns[33986] = 29'b1_000010011000_010_0_000100110001;
      patterns[33987] = 29'b1_000010011000_011_0_001001100010;
      patterns[33988] = 29'b1_000010011000_100_0_100001001100;
      patterns[33989] = 29'b1_000010011000_101_0_010000100110;
      patterns[33990] = 29'b1_000010011000_110_1_000010011000;
      patterns[33991] = 29'b1_000010011000_111_1_000010011000;
      patterns[33992] = 29'b1_000010011001_000_1_000010011001;
      patterns[33993] = 29'b1_000010011001_001_1_011001000010;
      patterns[33994] = 29'b1_000010011001_010_0_000100110011;
      patterns[33995] = 29'b1_000010011001_011_0_001001100110;
      patterns[33996] = 29'b1_000010011001_100_1_100001001100;
      patterns[33997] = 29'b1_000010011001_101_0_110000100110;
      patterns[33998] = 29'b1_000010011001_110_1_000010011001;
      patterns[33999] = 29'b1_000010011001_111_1_000010011001;
      patterns[34000] = 29'b1_000010011010_000_1_000010011010;
      patterns[34001] = 29'b1_000010011010_001_1_011010000010;
      patterns[34002] = 29'b1_000010011010_010_0_000100110101;
      patterns[34003] = 29'b1_000010011010_011_0_001001101010;
      patterns[34004] = 29'b1_000010011010_100_0_100001001101;
      patterns[34005] = 29'b1_000010011010_101_1_010000100110;
      patterns[34006] = 29'b1_000010011010_110_1_000010011010;
      patterns[34007] = 29'b1_000010011010_111_1_000010011010;
      patterns[34008] = 29'b1_000010011011_000_1_000010011011;
      patterns[34009] = 29'b1_000010011011_001_1_011011000010;
      patterns[34010] = 29'b1_000010011011_010_0_000100110111;
      patterns[34011] = 29'b1_000010011011_011_0_001001101110;
      patterns[34012] = 29'b1_000010011011_100_1_100001001101;
      patterns[34013] = 29'b1_000010011011_101_1_110000100110;
      patterns[34014] = 29'b1_000010011011_110_1_000010011011;
      patterns[34015] = 29'b1_000010011011_111_1_000010011011;
      patterns[34016] = 29'b1_000010011100_000_1_000010011100;
      patterns[34017] = 29'b1_000010011100_001_1_011100000010;
      patterns[34018] = 29'b1_000010011100_010_0_000100111001;
      patterns[34019] = 29'b1_000010011100_011_0_001001110010;
      patterns[34020] = 29'b1_000010011100_100_0_100001001110;
      patterns[34021] = 29'b1_000010011100_101_0_010000100111;
      patterns[34022] = 29'b1_000010011100_110_1_000010011100;
      patterns[34023] = 29'b1_000010011100_111_1_000010011100;
      patterns[34024] = 29'b1_000010011101_000_1_000010011101;
      patterns[34025] = 29'b1_000010011101_001_1_011101000010;
      patterns[34026] = 29'b1_000010011101_010_0_000100111011;
      patterns[34027] = 29'b1_000010011101_011_0_001001110110;
      patterns[34028] = 29'b1_000010011101_100_1_100001001110;
      patterns[34029] = 29'b1_000010011101_101_0_110000100111;
      patterns[34030] = 29'b1_000010011101_110_1_000010011101;
      patterns[34031] = 29'b1_000010011101_111_1_000010011101;
      patterns[34032] = 29'b1_000010011110_000_1_000010011110;
      patterns[34033] = 29'b1_000010011110_001_1_011110000010;
      patterns[34034] = 29'b1_000010011110_010_0_000100111101;
      patterns[34035] = 29'b1_000010011110_011_0_001001111010;
      patterns[34036] = 29'b1_000010011110_100_0_100001001111;
      patterns[34037] = 29'b1_000010011110_101_1_010000100111;
      patterns[34038] = 29'b1_000010011110_110_1_000010011110;
      patterns[34039] = 29'b1_000010011110_111_1_000010011110;
      patterns[34040] = 29'b1_000010011111_000_1_000010011111;
      patterns[34041] = 29'b1_000010011111_001_1_011111000010;
      patterns[34042] = 29'b1_000010011111_010_0_000100111111;
      patterns[34043] = 29'b1_000010011111_011_0_001001111110;
      patterns[34044] = 29'b1_000010011111_100_1_100001001111;
      patterns[34045] = 29'b1_000010011111_101_1_110000100111;
      patterns[34046] = 29'b1_000010011111_110_1_000010011111;
      patterns[34047] = 29'b1_000010011111_111_1_000010011111;
      patterns[34048] = 29'b1_000010100000_000_1_000010100000;
      patterns[34049] = 29'b1_000010100000_001_1_100000000010;
      patterns[34050] = 29'b1_000010100000_010_0_000101000001;
      patterns[34051] = 29'b1_000010100000_011_0_001010000010;
      patterns[34052] = 29'b1_000010100000_100_0_100001010000;
      patterns[34053] = 29'b1_000010100000_101_0_010000101000;
      patterns[34054] = 29'b1_000010100000_110_1_000010100000;
      patterns[34055] = 29'b1_000010100000_111_1_000010100000;
      patterns[34056] = 29'b1_000010100001_000_1_000010100001;
      patterns[34057] = 29'b1_000010100001_001_1_100001000010;
      patterns[34058] = 29'b1_000010100001_010_0_000101000011;
      patterns[34059] = 29'b1_000010100001_011_0_001010000110;
      patterns[34060] = 29'b1_000010100001_100_1_100001010000;
      patterns[34061] = 29'b1_000010100001_101_0_110000101000;
      patterns[34062] = 29'b1_000010100001_110_1_000010100001;
      patterns[34063] = 29'b1_000010100001_111_1_000010100001;
      patterns[34064] = 29'b1_000010100010_000_1_000010100010;
      patterns[34065] = 29'b1_000010100010_001_1_100010000010;
      patterns[34066] = 29'b1_000010100010_010_0_000101000101;
      patterns[34067] = 29'b1_000010100010_011_0_001010001010;
      patterns[34068] = 29'b1_000010100010_100_0_100001010001;
      patterns[34069] = 29'b1_000010100010_101_1_010000101000;
      patterns[34070] = 29'b1_000010100010_110_1_000010100010;
      patterns[34071] = 29'b1_000010100010_111_1_000010100010;
      patterns[34072] = 29'b1_000010100011_000_1_000010100011;
      patterns[34073] = 29'b1_000010100011_001_1_100011000010;
      patterns[34074] = 29'b1_000010100011_010_0_000101000111;
      patterns[34075] = 29'b1_000010100011_011_0_001010001110;
      patterns[34076] = 29'b1_000010100011_100_1_100001010001;
      patterns[34077] = 29'b1_000010100011_101_1_110000101000;
      patterns[34078] = 29'b1_000010100011_110_1_000010100011;
      patterns[34079] = 29'b1_000010100011_111_1_000010100011;
      patterns[34080] = 29'b1_000010100100_000_1_000010100100;
      patterns[34081] = 29'b1_000010100100_001_1_100100000010;
      patterns[34082] = 29'b1_000010100100_010_0_000101001001;
      patterns[34083] = 29'b1_000010100100_011_0_001010010010;
      patterns[34084] = 29'b1_000010100100_100_0_100001010010;
      patterns[34085] = 29'b1_000010100100_101_0_010000101001;
      patterns[34086] = 29'b1_000010100100_110_1_000010100100;
      patterns[34087] = 29'b1_000010100100_111_1_000010100100;
      patterns[34088] = 29'b1_000010100101_000_1_000010100101;
      patterns[34089] = 29'b1_000010100101_001_1_100101000010;
      patterns[34090] = 29'b1_000010100101_010_0_000101001011;
      patterns[34091] = 29'b1_000010100101_011_0_001010010110;
      patterns[34092] = 29'b1_000010100101_100_1_100001010010;
      patterns[34093] = 29'b1_000010100101_101_0_110000101001;
      patterns[34094] = 29'b1_000010100101_110_1_000010100101;
      patterns[34095] = 29'b1_000010100101_111_1_000010100101;
      patterns[34096] = 29'b1_000010100110_000_1_000010100110;
      patterns[34097] = 29'b1_000010100110_001_1_100110000010;
      patterns[34098] = 29'b1_000010100110_010_0_000101001101;
      patterns[34099] = 29'b1_000010100110_011_0_001010011010;
      patterns[34100] = 29'b1_000010100110_100_0_100001010011;
      patterns[34101] = 29'b1_000010100110_101_1_010000101001;
      patterns[34102] = 29'b1_000010100110_110_1_000010100110;
      patterns[34103] = 29'b1_000010100110_111_1_000010100110;
      patterns[34104] = 29'b1_000010100111_000_1_000010100111;
      patterns[34105] = 29'b1_000010100111_001_1_100111000010;
      patterns[34106] = 29'b1_000010100111_010_0_000101001111;
      patterns[34107] = 29'b1_000010100111_011_0_001010011110;
      patterns[34108] = 29'b1_000010100111_100_1_100001010011;
      patterns[34109] = 29'b1_000010100111_101_1_110000101001;
      patterns[34110] = 29'b1_000010100111_110_1_000010100111;
      patterns[34111] = 29'b1_000010100111_111_1_000010100111;
      patterns[34112] = 29'b1_000010101000_000_1_000010101000;
      patterns[34113] = 29'b1_000010101000_001_1_101000000010;
      patterns[34114] = 29'b1_000010101000_010_0_000101010001;
      patterns[34115] = 29'b1_000010101000_011_0_001010100010;
      patterns[34116] = 29'b1_000010101000_100_0_100001010100;
      patterns[34117] = 29'b1_000010101000_101_0_010000101010;
      patterns[34118] = 29'b1_000010101000_110_1_000010101000;
      patterns[34119] = 29'b1_000010101000_111_1_000010101000;
      patterns[34120] = 29'b1_000010101001_000_1_000010101001;
      patterns[34121] = 29'b1_000010101001_001_1_101001000010;
      patterns[34122] = 29'b1_000010101001_010_0_000101010011;
      patterns[34123] = 29'b1_000010101001_011_0_001010100110;
      patterns[34124] = 29'b1_000010101001_100_1_100001010100;
      patterns[34125] = 29'b1_000010101001_101_0_110000101010;
      patterns[34126] = 29'b1_000010101001_110_1_000010101001;
      patterns[34127] = 29'b1_000010101001_111_1_000010101001;
      patterns[34128] = 29'b1_000010101010_000_1_000010101010;
      patterns[34129] = 29'b1_000010101010_001_1_101010000010;
      patterns[34130] = 29'b1_000010101010_010_0_000101010101;
      patterns[34131] = 29'b1_000010101010_011_0_001010101010;
      patterns[34132] = 29'b1_000010101010_100_0_100001010101;
      patterns[34133] = 29'b1_000010101010_101_1_010000101010;
      patterns[34134] = 29'b1_000010101010_110_1_000010101010;
      patterns[34135] = 29'b1_000010101010_111_1_000010101010;
      patterns[34136] = 29'b1_000010101011_000_1_000010101011;
      patterns[34137] = 29'b1_000010101011_001_1_101011000010;
      patterns[34138] = 29'b1_000010101011_010_0_000101010111;
      patterns[34139] = 29'b1_000010101011_011_0_001010101110;
      patterns[34140] = 29'b1_000010101011_100_1_100001010101;
      patterns[34141] = 29'b1_000010101011_101_1_110000101010;
      patterns[34142] = 29'b1_000010101011_110_1_000010101011;
      patterns[34143] = 29'b1_000010101011_111_1_000010101011;
      patterns[34144] = 29'b1_000010101100_000_1_000010101100;
      patterns[34145] = 29'b1_000010101100_001_1_101100000010;
      patterns[34146] = 29'b1_000010101100_010_0_000101011001;
      patterns[34147] = 29'b1_000010101100_011_0_001010110010;
      patterns[34148] = 29'b1_000010101100_100_0_100001010110;
      patterns[34149] = 29'b1_000010101100_101_0_010000101011;
      patterns[34150] = 29'b1_000010101100_110_1_000010101100;
      patterns[34151] = 29'b1_000010101100_111_1_000010101100;
      patterns[34152] = 29'b1_000010101101_000_1_000010101101;
      patterns[34153] = 29'b1_000010101101_001_1_101101000010;
      patterns[34154] = 29'b1_000010101101_010_0_000101011011;
      patterns[34155] = 29'b1_000010101101_011_0_001010110110;
      patterns[34156] = 29'b1_000010101101_100_1_100001010110;
      patterns[34157] = 29'b1_000010101101_101_0_110000101011;
      patterns[34158] = 29'b1_000010101101_110_1_000010101101;
      patterns[34159] = 29'b1_000010101101_111_1_000010101101;
      patterns[34160] = 29'b1_000010101110_000_1_000010101110;
      patterns[34161] = 29'b1_000010101110_001_1_101110000010;
      patterns[34162] = 29'b1_000010101110_010_0_000101011101;
      patterns[34163] = 29'b1_000010101110_011_0_001010111010;
      patterns[34164] = 29'b1_000010101110_100_0_100001010111;
      patterns[34165] = 29'b1_000010101110_101_1_010000101011;
      patterns[34166] = 29'b1_000010101110_110_1_000010101110;
      patterns[34167] = 29'b1_000010101110_111_1_000010101110;
      patterns[34168] = 29'b1_000010101111_000_1_000010101111;
      patterns[34169] = 29'b1_000010101111_001_1_101111000010;
      patterns[34170] = 29'b1_000010101111_010_0_000101011111;
      patterns[34171] = 29'b1_000010101111_011_0_001010111110;
      patterns[34172] = 29'b1_000010101111_100_1_100001010111;
      patterns[34173] = 29'b1_000010101111_101_1_110000101011;
      patterns[34174] = 29'b1_000010101111_110_1_000010101111;
      patterns[34175] = 29'b1_000010101111_111_1_000010101111;
      patterns[34176] = 29'b1_000010110000_000_1_000010110000;
      patterns[34177] = 29'b1_000010110000_001_1_110000000010;
      patterns[34178] = 29'b1_000010110000_010_0_000101100001;
      patterns[34179] = 29'b1_000010110000_011_0_001011000010;
      patterns[34180] = 29'b1_000010110000_100_0_100001011000;
      patterns[34181] = 29'b1_000010110000_101_0_010000101100;
      patterns[34182] = 29'b1_000010110000_110_1_000010110000;
      patterns[34183] = 29'b1_000010110000_111_1_000010110000;
      patterns[34184] = 29'b1_000010110001_000_1_000010110001;
      patterns[34185] = 29'b1_000010110001_001_1_110001000010;
      patterns[34186] = 29'b1_000010110001_010_0_000101100011;
      patterns[34187] = 29'b1_000010110001_011_0_001011000110;
      patterns[34188] = 29'b1_000010110001_100_1_100001011000;
      patterns[34189] = 29'b1_000010110001_101_0_110000101100;
      patterns[34190] = 29'b1_000010110001_110_1_000010110001;
      patterns[34191] = 29'b1_000010110001_111_1_000010110001;
      patterns[34192] = 29'b1_000010110010_000_1_000010110010;
      patterns[34193] = 29'b1_000010110010_001_1_110010000010;
      patterns[34194] = 29'b1_000010110010_010_0_000101100101;
      patterns[34195] = 29'b1_000010110010_011_0_001011001010;
      patterns[34196] = 29'b1_000010110010_100_0_100001011001;
      patterns[34197] = 29'b1_000010110010_101_1_010000101100;
      patterns[34198] = 29'b1_000010110010_110_1_000010110010;
      patterns[34199] = 29'b1_000010110010_111_1_000010110010;
      patterns[34200] = 29'b1_000010110011_000_1_000010110011;
      patterns[34201] = 29'b1_000010110011_001_1_110011000010;
      patterns[34202] = 29'b1_000010110011_010_0_000101100111;
      patterns[34203] = 29'b1_000010110011_011_0_001011001110;
      patterns[34204] = 29'b1_000010110011_100_1_100001011001;
      patterns[34205] = 29'b1_000010110011_101_1_110000101100;
      patterns[34206] = 29'b1_000010110011_110_1_000010110011;
      patterns[34207] = 29'b1_000010110011_111_1_000010110011;
      patterns[34208] = 29'b1_000010110100_000_1_000010110100;
      patterns[34209] = 29'b1_000010110100_001_1_110100000010;
      patterns[34210] = 29'b1_000010110100_010_0_000101101001;
      patterns[34211] = 29'b1_000010110100_011_0_001011010010;
      patterns[34212] = 29'b1_000010110100_100_0_100001011010;
      patterns[34213] = 29'b1_000010110100_101_0_010000101101;
      patterns[34214] = 29'b1_000010110100_110_1_000010110100;
      patterns[34215] = 29'b1_000010110100_111_1_000010110100;
      patterns[34216] = 29'b1_000010110101_000_1_000010110101;
      patterns[34217] = 29'b1_000010110101_001_1_110101000010;
      patterns[34218] = 29'b1_000010110101_010_0_000101101011;
      patterns[34219] = 29'b1_000010110101_011_0_001011010110;
      patterns[34220] = 29'b1_000010110101_100_1_100001011010;
      patterns[34221] = 29'b1_000010110101_101_0_110000101101;
      patterns[34222] = 29'b1_000010110101_110_1_000010110101;
      patterns[34223] = 29'b1_000010110101_111_1_000010110101;
      patterns[34224] = 29'b1_000010110110_000_1_000010110110;
      patterns[34225] = 29'b1_000010110110_001_1_110110000010;
      patterns[34226] = 29'b1_000010110110_010_0_000101101101;
      patterns[34227] = 29'b1_000010110110_011_0_001011011010;
      patterns[34228] = 29'b1_000010110110_100_0_100001011011;
      patterns[34229] = 29'b1_000010110110_101_1_010000101101;
      patterns[34230] = 29'b1_000010110110_110_1_000010110110;
      patterns[34231] = 29'b1_000010110110_111_1_000010110110;
      patterns[34232] = 29'b1_000010110111_000_1_000010110111;
      patterns[34233] = 29'b1_000010110111_001_1_110111000010;
      patterns[34234] = 29'b1_000010110111_010_0_000101101111;
      patterns[34235] = 29'b1_000010110111_011_0_001011011110;
      patterns[34236] = 29'b1_000010110111_100_1_100001011011;
      patterns[34237] = 29'b1_000010110111_101_1_110000101101;
      patterns[34238] = 29'b1_000010110111_110_1_000010110111;
      patterns[34239] = 29'b1_000010110111_111_1_000010110111;
      patterns[34240] = 29'b1_000010111000_000_1_000010111000;
      patterns[34241] = 29'b1_000010111000_001_1_111000000010;
      patterns[34242] = 29'b1_000010111000_010_0_000101110001;
      patterns[34243] = 29'b1_000010111000_011_0_001011100010;
      patterns[34244] = 29'b1_000010111000_100_0_100001011100;
      patterns[34245] = 29'b1_000010111000_101_0_010000101110;
      patterns[34246] = 29'b1_000010111000_110_1_000010111000;
      patterns[34247] = 29'b1_000010111000_111_1_000010111000;
      patterns[34248] = 29'b1_000010111001_000_1_000010111001;
      patterns[34249] = 29'b1_000010111001_001_1_111001000010;
      patterns[34250] = 29'b1_000010111001_010_0_000101110011;
      patterns[34251] = 29'b1_000010111001_011_0_001011100110;
      patterns[34252] = 29'b1_000010111001_100_1_100001011100;
      patterns[34253] = 29'b1_000010111001_101_0_110000101110;
      patterns[34254] = 29'b1_000010111001_110_1_000010111001;
      patterns[34255] = 29'b1_000010111001_111_1_000010111001;
      patterns[34256] = 29'b1_000010111010_000_1_000010111010;
      patterns[34257] = 29'b1_000010111010_001_1_111010000010;
      patterns[34258] = 29'b1_000010111010_010_0_000101110101;
      patterns[34259] = 29'b1_000010111010_011_0_001011101010;
      patterns[34260] = 29'b1_000010111010_100_0_100001011101;
      patterns[34261] = 29'b1_000010111010_101_1_010000101110;
      patterns[34262] = 29'b1_000010111010_110_1_000010111010;
      patterns[34263] = 29'b1_000010111010_111_1_000010111010;
      patterns[34264] = 29'b1_000010111011_000_1_000010111011;
      patterns[34265] = 29'b1_000010111011_001_1_111011000010;
      patterns[34266] = 29'b1_000010111011_010_0_000101110111;
      patterns[34267] = 29'b1_000010111011_011_0_001011101110;
      patterns[34268] = 29'b1_000010111011_100_1_100001011101;
      patterns[34269] = 29'b1_000010111011_101_1_110000101110;
      patterns[34270] = 29'b1_000010111011_110_1_000010111011;
      patterns[34271] = 29'b1_000010111011_111_1_000010111011;
      patterns[34272] = 29'b1_000010111100_000_1_000010111100;
      patterns[34273] = 29'b1_000010111100_001_1_111100000010;
      patterns[34274] = 29'b1_000010111100_010_0_000101111001;
      patterns[34275] = 29'b1_000010111100_011_0_001011110010;
      patterns[34276] = 29'b1_000010111100_100_0_100001011110;
      patterns[34277] = 29'b1_000010111100_101_0_010000101111;
      patterns[34278] = 29'b1_000010111100_110_1_000010111100;
      patterns[34279] = 29'b1_000010111100_111_1_000010111100;
      patterns[34280] = 29'b1_000010111101_000_1_000010111101;
      patterns[34281] = 29'b1_000010111101_001_1_111101000010;
      patterns[34282] = 29'b1_000010111101_010_0_000101111011;
      patterns[34283] = 29'b1_000010111101_011_0_001011110110;
      patterns[34284] = 29'b1_000010111101_100_1_100001011110;
      patterns[34285] = 29'b1_000010111101_101_0_110000101111;
      patterns[34286] = 29'b1_000010111101_110_1_000010111101;
      patterns[34287] = 29'b1_000010111101_111_1_000010111101;
      patterns[34288] = 29'b1_000010111110_000_1_000010111110;
      patterns[34289] = 29'b1_000010111110_001_1_111110000010;
      patterns[34290] = 29'b1_000010111110_010_0_000101111101;
      patterns[34291] = 29'b1_000010111110_011_0_001011111010;
      patterns[34292] = 29'b1_000010111110_100_0_100001011111;
      patterns[34293] = 29'b1_000010111110_101_1_010000101111;
      patterns[34294] = 29'b1_000010111110_110_1_000010111110;
      patterns[34295] = 29'b1_000010111110_111_1_000010111110;
      patterns[34296] = 29'b1_000010111111_000_1_000010111111;
      patterns[34297] = 29'b1_000010111111_001_1_111111000010;
      patterns[34298] = 29'b1_000010111111_010_0_000101111111;
      patterns[34299] = 29'b1_000010111111_011_0_001011111110;
      patterns[34300] = 29'b1_000010111111_100_1_100001011111;
      patterns[34301] = 29'b1_000010111111_101_1_110000101111;
      patterns[34302] = 29'b1_000010111111_110_1_000010111111;
      patterns[34303] = 29'b1_000010111111_111_1_000010111111;
      patterns[34304] = 29'b1_000011000000_000_1_000011000000;
      patterns[34305] = 29'b1_000011000000_001_1_000000000011;
      patterns[34306] = 29'b1_000011000000_010_0_000110000001;
      patterns[34307] = 29'b1_000011000000_011_0_001100000010;
      patterns[34308] = 29'b1_000011000000_100_0_100001100000;
      patterns[34309] = 29'b1_000011000000_101_0_010000110000;
      patterns[34310] = 29'b1_000011000000_110_1_000011000000;
      patterns[34311] = 29'b1_000011000000_111_1_000011000000;
      patterns[34312] = 29'b1_000011000001_000_1_000011000001;
      patterns[34313] = 29'b1_000011000001_001_1_000001000011;
      patterns[34314] = 29'b1_000011000001_010_0_000110000011;
      patterns[34315] = 29'b1_000011000001_011_0_001100000110;
      patterns[34316] = 29'b1_000011000001_100_1_100001100000;
      patterns[34317] = 29'b1_000011000001_101_0_110000110000;
      patterns[34318] = 29'b1_000011000001_110_1_000011000001;
      patterns[34319] = 29'b1_000011000001_111_1_000011000001;
      patterns[34320] = 29'b1_000011000010_000_1_000011000010;
      patterns[34321] = 29'b1_000011000010_001_1_000010000011;
      patterns[34322] = 29'b1_000011000010_010_0_000110000101;
      patterns[34323] = 29'b1_000011000010_011_0_001100001010;
      patterns[34324] = 29'b1_000011000010_100_0_100001100001;
      patterns[34325] = 29'b1_000011000010_101_1_010000110000;
      patterns[34326] = 29'b1_000011000010_110_1_000011000010;
      patterns[34327] = 29'b1_000011000010_111_1_000011000010;
      patterns[34328] = 29'b1_000011000011_000_1_000011000011;
      patterns[34329] = 29'b1_000011000011_001_1_000011000011;
      patterns[34330] = 29'b1_000011000011_010_0_000110000111;
      patterns[34331] = 29'b1_000011000011_011_0_001100001110;
      patterns[34332] = 29'b1_000011000011_100_1_100001100001;
      patterns[34333] = 29'b1_000011000011_101_1_110000110000;
      patterns[34334] = 29'b1_000011000011_110_1_000011000011;
      patterns[34335] = 29'b1_000011000011_111_1_000011000011;
      patterns[34336] = 29'b1_000011000100_000_1_000011000100;
      patterns[34337] = 29'b1_000011000100_001_1_000100000011;
      patterns[34338] = 29'b1_000011000100_010_0_000110001001;
      patterns[34339] = 29'b1_000011000100_011_0_001100010010;
      patterns[34340] = 29'b1_000011000100_100_0_100001100010;
      patterns[34341] = 29'b1_000011000100_101_0_010000110001;
      patterns[34342] = 29'b1_000011000100_110_1_000011000100;
      patterns[34343] = 29'b1_000011000100_111_1_000011000100;
      patterns[34344] = 29'b1_000011000101_000_1_000011000101;
      patterns[34345] = 29'b1_000011000101_001_1_000101000011;
      patterns[34346] = 29'b1_000011000101_010_0_000110001011;
      patterns[34347] = 29'b1_000011000101_011_0_001100010110;
      patterns[34348] = 29'b1_000011000101_100_1_100001100010;
      patterns[34349] = 29'b1_000011000101_101_0_110000110001;
      patterns[34350] = 29'b1_000011000101_110_1_000011000101;
      patterns[34351] = 29'b1_000011000101_111_1_000011000101;
      patterns[34352] = 29'b1_000011000110_000_1_000011000110;
      patterns[34353] = 29'b1_000011000110_001_1_000110000011;
      patterns[34354] = 29'b1_000011000110_010_0_000110001101;
      patterns[34355] = 29'b1_000011000110_011_0_001100011010;
      patterns[34356] = 29'b1_000011000110_100_0_100001100011;
      patterns[34357] = 29'b1_000011000110_101_1_010000110001;
      patterns[34358] = 29'b1_000011000110_110_1_000011000110;
      patterns[34359] = 29'b1_000011000110_111_1_000011000110;
      patterns[34360] = 29'b1_000011000111_000_1_000011000111;
      patterns[34361] = 29'b1_000011000111_001_1_000111000011;
      patterns[34362] = 29'b1_000011000111_010_0_000110001111;
      patterns[34363] = 29'b1_000011000111_011_0_001100011110;
      patterns[34364] = 29'b1_000011000111_100_1_100001100011;
      patterns[34365] = 29'b1_000011000111_101_1_110000110001;
      patterns[34366] = 29'b1_000011000111_110_1_000011000111;
      patterns[34367] = 29'b1_000011000111_111_1_000011000111;
      patterns[34368] = 29'b1_000011001000_000_1_000011001000;
      patterns[34369] = 29'b1_000011001000_001_1_001000000011;
      patterns[34370] = 29'b1_000011001000_010_0_000110010001;
      patterns[34371] = 29'b1_000011001000_011_0_001100100010;
      patterns[34372] = 29'b1_000011001000_100_0_100001100100;
      patterns[34373] = 29'b1_000011001000_101_0_010000110010;
      patterns[34374] = 29'b1_000011001000_110_1_000011001000;
      patterns[34375] = 29'b1_000011001000_111_1_000011001000;
      patterns[34376] = 29'b1_000011001001_000_1_000011001001;
      patterns[34377] = 29'b1_000011001001_001_1_001001000011;
      patterns[34378] = 29'b1_000011001001_010_0_000110010011;
      patterns[34379] = 29'b1_000011001001_011_0_001100100110;
      patterns[34380] = 29'b1_000011001001_100_1_100001100100;
      patterns[34381] = 29'b1_000011001001_101_0_110000110010;
      patterns[34382] = 29'b1_000011001001_110_1_000011001001;
      patterns[34383] = 29'b1_000011001001_111_1_000011001001;
      patterns[34384] = 29'b1_000011001010_000_1_000011001010;
      patterns[34385] = 29'b1_000011001010_001_1_001010000011;
      patterns[34386] = 29'b1_000011001010_010_0_000110010101;
      patterns[34387] = 29'b1_000011001010_011_0_001100101010;
      patterns[34388] = 29'b1_000011001010_100_0_100001100101;
      patterns[34389] = 29'b1_000011001010_101_1_010000110010;
      patterns[34390] = 29'b1_000011001010_110_1_000011001010;
      patterns[34391] = 29'b1_000011001010_111_1_000011001010;
      patterns[34392] = 29'b1_000011001011_000_1_000011001011;
      patterns[34393] = 29'b1_000011001011_001_1_001011000011;
      patterns[34394] = 29'b1_000011001011_010_0_000110010111;
      patterns[34395] = 29'b1_000011001011_011_0_001100101110;
      patterns[34396] = 29'b1_000011001011_100_1_100001100101;
      patterns[34397] = 29'b1_000011001011_101_1_110000110010;
      patterns[34398] = 29'b1_000011001011_110_1_000011001011;
      patterns[34399] = 29'b1_000011001011_111_1_000011001011;
      patterns[34400] = 29'b1_000011001100_000_1_000011001100;
      patterns[34401] = 29'b1_000011001100_001_1_001100000011;
      patterns[34402] = 29'b1_000011001100_010_0_000110011001;
      patterns[34403] = 29'b1_000011001100_011_0_001100110010;
      patterns[34404] = 29'b1_000011001100_100_0_100001100110;
      patterns[34405] = 29'b1_000011001100_101_0_010000110011;
      patterns[34406] = 29'b1_000011001100_110_1_000011001100;
      patterns[34407] = 29'b1_000011001100_111_1_000011001100;
      patterns[34408] = 29'b1_000011001101_000_1_000011001101;
      patterns[34409] = 29'b1_000011001101_001_1_001101000011;
      patterns[34410] = 29'b1_000011001101_010_0_000110011011;
      patterns[34411] = 29'b1_000011001101_011_0_001100110110;
      patterns[34412] = 29'b1_000011001101_100_1_100001100110;
      patterns[34413] = 29'b1_000011001101_101_0_110000110011;
      patterns[34414] = 29'b1_000011001101_110_1_000011001101;
      patterns[34415] = 29'b1_000011001101_111_1_000011001101;
      patterns[34416] = 29'b1_000011001110_000_1_000011001110;
      patterns[34417] = 29'b1_000011001110_001_1_001110000011;
      patterns[34418] = 29'b1_000011001110_010_0_000110011101;
      patterns[34419] = 29'b1_000011001110_011_0_001100111010;
      patterns[34420] = 29'b1_000011001110_100_0_100001100111;
      patterns[34421] = 29'b1_000011001110_101_1_010000110011;
      patterns[34422] = 29'b1_000011001110_110_1_000011001110;
      patterns[34423] = 29'b1_000011001110_111_1_000011001110;
      patterns[34424] = 29'b1_000011001111_000_1_000011001111;
      patterns[34425] = 29'b1_000011001111_001_1_001111000011;
      patterns[34426] = 29'b1_000011001111_010_0_000110011111;
      patterns[34427] = 29'b1_000011001111_011_0_001100111110;
      patterns[34428] = 29'b1_000011001111_100_1_100001100111;
      patterns[34429] = 29'b1_000011001111_101_1_110000110011;
      patterns[34430] = 29'b1_000011001111_110_1_000011001111;
      patterns[34431] = 29'b1_000011001111_111_1_000011001111;
      patterns[34432] = 29'b1_000011010000_000_1_000011010000;
      patterns[34433] = 29'b1_000011010000_001_1_010000000011;
      patterns[34434] = 29'b1_000011010000_010_0_000110100001;
      patterns[34435] = 29'b1_000011010000_011_0_001101000010;
      patterns[34436] = 29'b1_000011010000_100_0_100001101000;
      patterns[34437] = 29'b1_000011010000_101_0_010000110100;
      patterns[34438] = 29'b1_000011010000_110_1_000011010000;
      patterns[34439] = 29'b1_000011010000_111_1_000011010000;
      patterns[34440] = 29'b1_000011010001_000_1_000011010001;
      patterns[34441] = 29'b1_000011010001_001_1_010001000011;
      patterns[34442] = 29'b1_000011010001_010_0_000110100011;
      patterns[34443] = 29'b1_000011010001_011_0_001101000110;
      patterns[34444] = 29'b1_000011010001_100_1_100001101000;
      patterns[34445] = 29'b1_000011010001_101_0_110000110100;
      patterns[34446] = 29'b1_000011010001_110_1_000011010001;
      patterns[34447] = 29'b1_000011010001_111_1_000011010001;
      patterns[34448] = 29'b1_000011010010_000_1_000011010010;
      patterns[34449] = 29'b1_000011010010_001_1_010010000011;
      patterns[34450] = 29'b1_000011010010_010_0_000110100101;
      patterns[34451] = 29'b1_000011010010_011_0_001101001010;
      patterns[34452] = 29'b1_000011010010_100_0_100001101001;
      patterns[34453] = 29'b1_000011010010_101_1_010000110100;
      patterns[34454] = 29'b1_000011010010_110_1_000011010010;
      patterns[34455] = 29'b1_000011010010_111_1_000011010010;
      patterns[34456] = 29'b1_000011010011_000_1_000011010011;
      patterns[34457] = 29'b1_000011010011_001_1_010011000011;
      patterns[34458] = 29'b1_000011010011_010_0_000110100111;
      patterns[34459] = 29'b1_000011010011_011_0_001101001110;
      patterns[34460] = 29'b1_000011010011_100_1_100001101001;
      patterns[34461] = 29'b1_000011010011_101_1_110000110100;
      patterns[34462] = 29'b1_000011010011_110_1_000011010011;
      patterns[34463] = 29'b1_000011010011_111_1_000011010011;
      patterns[34464] = 29'b1_000011010100_000_1_000011010100;
      patterns[34465] = 29'b1_000011010100_001_1_010100000011;
      patterns[34466] = 29'b1_000011010100_010_0_000110101001;
      patterns[34467] = 29'b1_000011010100_011_0_001101010010;
      patterns[34468] = 29'b1_000011010100_100_0_100001101010;
      patterns[34469] = 29'b1_000011010100_101_0_010000110101;
      patterns[34470] = 29'b1_000011010100_110_1_000011010100;
      patterns[34471] = 29'b1_000011010100_111_1_000011010100;
      patterns[34472] = 29'b1_000011010101_000_1_000011010101;
      patterns[34473] = 29'b1_000011010101_001_1_010101000011;
      patterns[34474] = 29'b1_000011010101_010_0_000110101011;
      patterns[34475] = 29'b1_000011010101_011_0_001101010110;
      patterns[34476] = 29'b1_000011010101_100_1_100001101010;
      patterns[34477] = 29'b1_000011010101_101_0_110000110101;
      patterns[34478] = 29'b1_000011010101_110_1_000011010101;
      patterns[34479] = 29'b1_000011010101_111_1_000011010101;
      patterns[34480] = 29'b1_000011010110_000_1_000011010110;
      patterns[34481] = 29'b1_000011010110_001_1_010110000011;
      patterns[34482] = 29'b1_000011010110_010_0_000110101101;
      patterns[34483] = 29'b1_000011010110_011_0_001101011010;
      patterns[34484] = 29'b1_000011010110_100_0_100001101011;
      patterns[34485] = 29'b1_000011010110_101_1_010000110101;
      patterns[34486] = 29'b1_000011010110_110_1_000011010110;
      patterns[34487] = 29'b1_000011010110_111_1_000011010110;
      patterns[34488] = 29'b1_000011010111_000_1_000011010111;
      patterns[34489] = 29'b1_000011010111_001_1_010111000011;
      patterns[34490] = 29'b1_000011010111_010_0_000110101111;
      patterns[34491] = 29'b1_000011010111_011_0_001101011110;
      patterns[34492] = 29'b1_000011010111_100_1_100001101011;
      patterns[34493] = 29'b1_000011010111_101_1_110000110101;
      patterns[34494] = 29'b1_000011010111_110_1_000011010111;
      patterns[34495] = 29'b1_000011010111_111_1_000011010111;
      patterns[34496] = 29'b1_000011011000_000_1_000011011000;
      patterns[34497] = 29'b1_000011011000_001_1_011000000011;
      patterns[34498] = 29'b1_000011011000_010_0_000110110001;
      patterns[34499] = 29'b1_000011011000_011_0_001101100010;
      patterns[34500] = 29'b1_000011011000_100_0_100001101100;
      patterns[34501] = 29'b1_000011011000_101_0_010000110110;
      patterns[34502] = 29'b1_000011011000_110_1_000011011000;
      patterns[34503] = 29'b1_000011011000_111_1_000011011000;
      patterns[34504] = 29'b1_000011011001_000_1_000011011001;
      patterns[34505] = 29'b1_000011011001_001_1_011001000011;
      patterns[34506] = 29'b1_000011011001_010_0_000110110011;
      patterns[34507] = 29'b1_000011011001_011_0_001101100110;
      patterns[34508] = 29'b1_000011011001_100_1_100001101100;
      patterns[34509] = 29'b1_000011011001_101_0_110000110110;
      patterns[34510] = 29'b1_000011011001_110_1_000011011001;
      patterns[34511] = 29'b1_000011011001_111_1_000011011001;
      patterns[34512] = 29'b1_000011011010_000_1_000011011010;
      patterns[34513] = 29'b1_000011011010_001_1_011010000011;
      patterns[34514] = 29'b1_000011011010_010_0_000110110101;
      patterns[34515] = 29'b1_000011011010_011_0_001101101010;
      patterns[34516] = 29'b1_000011011010_100_0_100001101101;
      patterns[34517] = 29'b1_000011011010_101_1_010000110110;
      patterns[34518] = 29'b1_000011011010_110_1_000011011010;
      patterns[34519] = 29'b1_000011011010_111_1_000011011010;
      patterns[34520] = 29'b1_000011011011_000_1_000011011011;
      patterns[34521] = 29'b1_000011011011_001_1_011011000011;
      patterns[34522] = 29'b1_000011011011_010_0_000110110111;
      patterns[34523] = 29'b1_000011011011_011_0_001101101110;
      patterns[34524] = 29'b1_000011011011_100_1_100001101101;
      patterns[34525] = 29'b1_000011011011_101_1_110000110110;
      patterns[34526] = 29'b1_000011011011_110_1_000011011011;
      patterns[34527] = 29'b1_000011011011_111_1_000011011011;
      patterns[34528] = 29'b1_000011011100_000_1_000011011100;
      patterns[34529] = 29'b1_000011011100_001_1_011100000011;
      patterns[34530] = 29'b1_000011011100_010_0_000110111001;
      patterns[34531] = 29'b1_000011011100_011_0_001101110010;
      patterns[34532] = 29'b1_000011011100_100_0_100001101110;
      patterns[34533] = 29'b1_000011011100_101_0_010000110111;
      patterns[34534] = 29'b1_000011011100_110_1_000011011100;
      patterns[34535] = 29'b1_000011011100_111_1_000011011100;
      patterns[34536] = 29'b1_000011011101_000_1_000011011101;
      patterns[34537] = 29'b1_000011011101_001_1_011101000011;
      patterns[34538] = 29'b1_000011011101_010_0_000110111011;
      patterns[34539] = 29'b1_000011011101_011_0_001101110110;
      patterns[34540] = 29'b1_000011011101_100_1_100001101110;
      patterns[34541] = 29'b1_000011011101_101_0_110000110111;
      patterns[34542] = 29'b1_000011011101_110_1_000011011101;
      patterns[34543] = 29'b1_000011011101_111_1_000011011101;
      patterns[34544] = 29'b1_000011011110_000_1_000011011110;
      patterns[34545] = 29'b1_000011011110_001_1_011110000011;
      patterns[34546] = 29'b1_000011011110_010_0_000110111101;
      patterns[34547] = 29'b1_000011011110_011_0_001101111010;
      patterns[34548] = 29'b1_000011011110_100_0_100001101111;
      patterns[34549] = 29'b1_000011011110_101_1_010000110111;
      patterns[34550] = 29'b1_000011011110_110_1_000011011110;
      patterns[34551] = 29'b1_000011011110_111_1_000011011110;
      patterns[34552] = 29'b1_000011011111_000_1_000011011111;
      patterns[34553] = 29'b1_000011011111_001_1_011111000011;
      patterns[34554] = 29'b1_000011011111_010_0_000110111111;
      patterns[34555] = 29'b1_000011011111_011_0_001101111110;
      patterns[34556] = 29'b1_000011011111_100_1_100001101111;
      patterns[34557] = 29'b1_000011011111_101_1_110000110111;
      patterns[34558] = 29'b1_000011011111_110_1_000011011111;
      patterns[34559] = 29'b1_000011011111_111_1_000011011111;
      patterns[34560] = 29'b1_000011100000_000_1_000011100000;
      patterns[34561] = 29'b1_000011100000_001_1_100000000011;
      patterns[34562] = 29'b1_000011100000_010_0_000111000001;
      patterns[34563] = 29'b1_000011100000_011_0_001110000010;
      patterns[34564] = 29'b1_000011100000_100_0_100001110000;
      patterns[34565] = 29'b1_000011100000_101_0_010000111000;
      patterns[34566] = 29'b1_000011100000_110_1_000011100000;
      patterns[34567] = 29'b1_000011100000_111_1_000011100000;
      patterns[34568] = 29'b1_000011100001_000_1_000011100001;
      patterns[34569] = 29'b1_000011100001_001_1_100001000011;
      patterns[34570] = 29'b1_000011100001_010_0_000111000011;
      patterns[34571] = 29'b1_000011100001_011_0_001110000110;
      patterns[34572] = 29'b1_000011100001_100_1_100001110000;
      patterns[34573] = 29'b1_000011100001_101_0_110000111000;
      patterns[34574] = 29'b1_000011100001_110_1_000011100001;
      patterns[34575] = 29'b1_000011100001_111_1_000011100001;
      patterns[34576] = 29'b1_000011100010_000_1_000011100010;
      patterns[34577] = 29'b1_000011100010_001_1_100010000011;
      patterns[34578] = 29'b1_000011100010_010_0_000111000101;
      patterns[34579] = 29'b1_000011100010_011_0_001110001010;
      patterns[34580] = 29'b1_000011100010_100_0_100001110001;
      patterns[34581] = 29'b1_000011100010_101_1_010000111000;
      patterns[34582] = 29'b1_000011100010_110_1_000011100010;
      patterns[34583] = 29'b1_000011100010_111_1_000011100010;
      patterns[34584] = 29'b1_000011100011_000_1_000011100011;
      patterns[34585] = 29'b1_000011100011_001_1_100011000011;
      patterns[34586] = 29'b1_000011100011_010_0_000111000111;
      patterns[34587] = 29'b1_000011100011_011_0_001110001110;
      patterns[34588] = 29'b1_000011100011_100_1_100001110001;
      patterns[34589] = 29'b1_000011100011_101_1_110000111000;
      patterns[34590] = 29'b1_000011100011_110_1_000011100011;
      patterns[34591] = 29'b1_000011100011_111_1_000011100011;
      patterns[34592] = 29'b1_000011100100_000_1_000011100100;
      patterns[34593] = 29'b1_000011100100_001_1_100100000011;
      patterns[34594] = 29'b1_000011100100_010_0_000111001001;
      patterns[34595] = 29'b1_000011100100_011_0_001110010010;
      patterns[34596] = 29'b1_000011100100_100_0_100001110010;
      patterns[34597] = 29'b1_000011100100_101_0_010000111001;
      patterns[34598] = 29'b1_000011100100_110_1_000011100100;
      patterns[34599] = 29'b1_000011100100_111_1_000011100100;
      patterns[34600] = 29'b1_000011100101_000_1_000011100101;
      patterns[34601] = 29'b1_000011100101_001_1_100101000011;
      patterns[34602] = 29'b1_000011100101_010_0_000111001011;
      patterns[34603] = 29'b1_000011100101_011_0_001110010110;
      patterns[34604] = 29'b1_000011100101_100_1_100001110010;
      patterns[34605] = 29'b1_000011100101_101_0_110000111001;
      patterns[34606] = 29'b1_000011100101_110_1_000011100101;
      patterns[34607] = 29'b1_000011100101_111_1_000011100101;
      patterns[34608] = 29'b1_000011100110_000_1_000011100110;
      patterns[34609] = 29'b1_000011100110_001_1_100110000011;
      patterns[34610] = 29'b1_000011100110_010_0_000111001101;
      patterns[34611] = 29'b1_000011100110_011_0_001110011010;
      patterns[34612] = 29'b1_000011100110_100_0_100001110011;
      patterns[34613] = 29'b1_000011100110_101_1_010000111001;
      patterns[34614] = 29'b1_000011100110_110_1_000011100110;
      patterns[34615] = 29'b1_000011100110_111_1_000011100110;
      patterns[34616] = 29'b1_000011100111_000_1_000011100111;
      patterns[34617] = 29'b1_000011100111_001_1_100111000011;
      patterns[34618] = 29'b1_000011100111_010_0_000111001111;
      patterns[34619] = 29'b1_000011100111_011_0_001110011110;
      patterns[34620] = 29'b1_000011100111_100_1_100001110011;
      patterns[34621] = 29'b1_000011100111_101_1_110000111001;
      patterns[34622] = 29'b1_000011100111_110_1_000011100111;
      patterns[34623] = 29'b1_000011100111_111_1_000011100111;
      patterns[34624] = 29'b1_000011101000_000_1_000011101000;
      patterns[34625] = 29'b1_000011101000_001_1_101000000011;
      patterns[34626] = 29'b1_000011101000_010_0_000111010001;
      patterns[34627] = 29'b1_000011101000_011_0_001110100010;
      patterns[34628] = 29'b1_000011101000_100_0_100001110100;
      patterns[34629] = 29'b1_000011101000_101_0_010000111010;
      patterns[34630] = 29'b1_000011101000_110_1_000011101000;
      patterns[34631] = 29'b1_000011101000_111_1_000011101000;
      patterns[34632] = 29'b1_000011101001_000_1_000011101001;
      patterns[34633] = 29'b1_000011101001_001_1_101001000011;
      patterns[34634] = 29'b1_000011101001_010_0_000111010011;
      patterns[34635] = 29'b1_000011101001_011_0_001110100110;
      patterns[34636] = 29'b1_000011101001_100_1_100001110100;
      patterns[34637] = 29'b1_000011101001_101_0_110000111010;
      patterns[34638] = 29'b1_000011101001_110_1_000011101001;
      patterns[34639] = 29'b1_000011101001_111_1_000011101001;
      patterns[34640] = 29'b1_000011101010_000_1_000011101010;
      patterns[34641] = 29'b1_000011101010_001_1_101010000011;
      patterns[34642] = 29'b1_000011101010_010_0_000111010101;
      patterns[34643] = 29'b1_000011101010_011_0_001110101010;
      patterns[34644] = 29'b1_000011101010_100_0_100001110101;
      patterns[34645] = 29'b1_000011101010_101_1_010000111010;
      patterns[34646] = 29'b1_000011101010_110_1_000011101010;
      patterns[34647] = 29'b1_000011101010_111_1_000011101010;
      patterns[34648] = 29'b1_000011101011_000_1_000011101011;
      patterns[34649] = 29'b1_000011101011_001_1_101011000011;
      patterns[34650] = 29'b1_000011101011_010_0_000111010111;
      patterns[34651] = 29'b1_000011101011_011_0_001110101110;
      patterns[34652] = 29'b1_000011101011_100_1_100001110101;
      patterns[34653] = 29'b1_000011101011_101_1_110000111010;
      patterns[34654] = 29'b1_000011101011_110_1_000011101011;
      patterns[34655] = 29'b1_000011101011_111_1_000011101011;
      patterns[34656] = 29'b1_000011101100_000_1_000011101100;
      patterns[34657] = 29'b1_000011101100_001_1_101100000011;
      patterns[34658] = 29'b1_000011101100_010_0_000111011001;
      patterns[34659] = 29'b1_000011101100_011_0_001110110010;
      patterns[34660] = 29'b1_000011101100_100_0_100001110110;
      patterns[34661] = 29'b1_000011101100_101_0_010000111011;
      patterns[34662] = 29'b1_000011101100_110_1_000011101100;
      patterns[34663] = 29'b1_000011101100_111_1_000011101100;
      patterns[34664] = 29'b1_000011101101_000_1_000011101101;
      patterns[34665] = 29'b1_000011101101_001_1_101101000011;
      patterns[34666] = 29'b1_000011101101_010_0_000111011011;
      patterns[34667] = 29'b1_000011101101_011_0_001110110110;
      patterns[34668] = 29'b1_000011101101_100_1_100001110110;
      patterns[34669] = 29'b1_000011101101_101_0_110000111011;
      patterns[34670] = 29'b1_000011101101_110_1_000011101101;
      patterns[34671] = 29'b1_000011101101_111_1_000011101101;
      patterns[34672] = 29'b1_000011101110_000_1_000011101110;
      patterns[34673] = 29'b1_000011101110_001_1_101110000011;
      patterns[34674] = 29'b1_000011101110_010_0_000111011101;
      patterns[34675] = 29'b1_000011101110_011_0_001110111010;
      patterns[34676] = 29'b1_000011101110_100_0_100001110111;
      patterns[34677] = 29'b1_000011101110_101_1_010000111011;
      patterns[34678] = 29'b1_000011101110_110_1_000011101110;
      patterns[34679] = 29'b1_000011101110_111_1_000011101110;
      patterns[34680] = 29'b1_000011101111_000_1_000011101111;
      patterns[34681] = 29'b1_000011101111_001_1_101111000011;
      patterns[34682] = 29'b1_000011101111_010_0_000111011111;
      patterns[34683] = 29'b1_000011101111_011_0_001110111110;
      patterns[34684] = 29'b1_000011101111_100_1_100001110111;
      patterns[34685] = 29'b1_000011101111_101_1_110000111011;
      patterns[34686] = 29'b1_000011101111_110_1_000011101111;
      patterns[34687] = 29'b1_000011101111_111_1_000011101111;
      patterns[34688] = 29'b1_000011110000_000_1_000011110000;
      patterns[34689] = 29'b1_000011110000_001_1_110000000011;
      patterns[34690] = 29'b1_000011110000_010_0_000111100001;
      patterns[34691] = 29'b1_000011110000_011_0_001111000010;
      patterns[34692] = 29'b1_000011110000_100_0_100001111000;
      patterns[34693] = 29'b1_000011110000_101_0_010000111100;
      patterns[34694] = 29'b1_000011110000_110_1_000011110000;
      patterns[34695] = 29'b1_000011110000_111_1_000011110000;
      patterns[34696] = 29'b1_000011110001_000_1_000011110001;
      patterns[34697] = 29'b1_000011110001_001_1_110001000011;
      patterns[34698] = 29'b1_000011110001_010_0_000111100011;
      patterns[34699] = 29'b1_000011110001_011_0_001111000110;
      patterns[34700] = 29'b1_000011110001_100_1_100001111000;
      patterns[34701] = 29'b1_000011110001_101_0_110000111100;
      patterns[34702] = 29'b1_000011110001_110_1_000011110001;
      patterns[34703] = 29'b1_000011110001_111_1_000011110001;
      patterns[34704] = 29'b1_000011110010_000_1_000011110010;
      patterns[34705] = 29'b1_000011110010_001_1_110010000011;
      patterns[34706] = 29'b1_000011110010_010_0_000111100101;
      patterns[34707] = 29'b1_000011110010_011_0_001111001010;
      patterns[34708] = 29'b1_000011110010_100_0_100001111001;
      patterns[34709] = 29'b1_000011110010_101_1_010000111100;
      patterns[34710] = 29'b1_000011110010_110_1_000011110010;
      patterns[34711] = 29'b1_000011110010_111_1_000011110010;
      patterns[34712] = 29'b1_000011110011_000_1_000011110011;
      patterns[34713] = 29'b1_000011110011_001_1_110011000011;
      patterns[34714] = 29'b1_000011110011_010_0_000111100111;
      patterns[34715] = 29'b1_000011110011_011_0_001111001110;
      patterns[34716] = 29'b1_000011110011_100_1_100001111001;
      patterns[34717] = 29'b1_000011110011_101_1_110000111100;
      patterns[34718] = 29'b1_000011110011_110_1_000011110011;
      patterns[34719] = 29'b1_000011110011_111_1_000011110011;
      patterns[34720] = 29'b1_000011110100_000_1_000011110100;
      patterns[34721] = 29'b1_000011110100_001_1_110100000011;
      patterns[34722] = 29'b1_000011110100_010_0_000111101001;
      patterns[34723] = 29'b1_000011110100_011_0_001111010010;
      patterns[34724] = 29'b1_000011110100_100_0_100001111010;
      patterns[34725] = 29'b1_000011110100_101_0_010000111101;
      patterns[34726] = 29'b1_000011110100_110_1_000011110100;
      patterns[34727] = 29'b1_000011110100_111_1_000011110100;
      patterns[34728] = 29'b1_000011110101_000_1_000011110101;
      patterns[34729] = 29'b1_000011110101_001_1_110101000011;
      patterns[34730] = 29'b1_000011110101_010_0_000111101011;
      patterns[34731] = 29'b1_000011110101_011_0_001111010110;
      patterns[34732] = 29'b1_000011110101_100_1_100001111010;
      patterns[34733] = 29'b1_000011110101_101_0_110000111101;
      patterns[34734] = 29'b1_000011110101_110_1_000011110101;
      patterns[34735] = 29'b1_000011110101_111_1_000011110101;
      patterns[34736] = 29'b1_000011110110_000_1_000011110110;
      patterns[34737] = 29'b1_000011110110_001_1_110110000011;
      patterns[34738] = 29'b1_000011110110_010_0_000111101101;
      patterns[34739] = 29'b1_000011110110_011_0_001111011010;
      patterns[34740] = 29'b1_000011110110_100_0_100001111011;
      patterns[34741] = 29'b1_000011110110_101_1_010000111101;
      patterns[34742] = 29'b1_000011110110_110_1_000011110110;
      patterns[34743] = 29'b1_000011110110_111_1_000011110110;
      patterns[34744] = 29'b1_000011110111_000_1_000011110111;
      patterns[34745] = 29'b1_000011110111_001_1_110111000011;
      patterns[34746] = 29'b1_000011110111_010_0_000111101111;
      patterns[34747] = 29'b1_000011110111_011_0_001111011110;
      patterns[34748] = 29'b1_000011110111_100_1_100001111011;
      patterns[34749] = 29'b1_000011110111_101_1_110000111101;
      patterns[34750] = 29'b1_000011110111_110_1_000011110111;
      patterns[34751] = 29'b1_000011110111_111_1_000011110111;
      patterns[34752] = 29'b1_000011111000_000_1_000011111000;
      patterns[34753] = 29'b1_000011111000_001_1_111000000011;
      patterns[34754] = 29'b1_000011111000_010_0_000111110001;
      patterns[34755] = 29'b1_000011111000_011_0_001111100010;
      patterns[34756] = 29'b1_000011111000_100_0_100001111100;
      patterns[34757] = 29'b1_000011111000_101_0_010000111110;
      patterns[34758] = 29'b1_000011111000_110_1_000011111000;
      patterns[34759] = 29'b1_000011111000_111_1_000011111000;
      patterns[34760] = 29'b1_000011111001_000_1_000011111001;
      patterns[34761] = 29'b1_000011111001_001_1_111001000011;
      patterns[34762] = 29'b1_000011111001_010_0_000111110011;
      patterns[34763] = 29'b1_000011111001_011_0_001111100110;
      patterns[34764] = 29'b1_000011111001_100_1_100001111100;
      patterns[34765] = 29'b1_000011111001_101_0_110000111110;
      patterns[34766] = 29'b1_000011111001_110_1_000011111001;
      patterns[34767] = 29'b1_000011111001_111_1_000011111001;
      patterns[34768] = 29'b1_000011111010_000_1_000011111010;
      patterns[34769] = 29'b1_000011111010_001_1_111010000011;
      patterns[34770] = 29'b1_000011111010_010_0_000111110101;
      patterns[34771] = 29'b1_000011111010_011_0_001111101010;
      patterns[34772] = 29'b1_000011111010_100_0_100001111101;
      patterns[34773] = 29'b1_000011111010_101_1_010000111110;
      patterns[34774] = 29'b1_000011111010_110_1_000011111010;
      patterns[34775] = 29'b1_000011111010_111_1_000011111010;
      patterns[34776] = 29'b1_000011111011_000_1_000011111011;
      patterns[34777] = 29'b1_000011111011_001_1_111011000011;
      patterns[34778] = 29'b1_000011111011_010_0_000111110111;
      patterns[34779] = 29'b1_000011111011_011_0_001111101110;
      patterns[34780] = 29'b1_000011111011_100_1_100001111101;
      patterns[34781] = 29'b1_000011111011_101_1_110000111110;
      patterns[34782] = 29'b1_000011111011_110_1_000011111011;
      patterns[34783] = 29'b1_000011111011_111_1_000011111011;
      patterns[34784] = 29'b1_000011111100_000_1_000011111100;
      patterns[34785] = 29'b1_000011111100_001_1_111100000011;
      patterns[34786] = 29'b1_000011111100_010_0_000111111001;
      patterns[34787] = 29'b1_000011111100_011_0_001111110010;
      patterns[34788] = 29'b1_000011111100_100_0_100001111110;
      patterns[34789] = 29'b1_000011111100_101_0_010000111111;
      patterns[34790] = 29'b1_000011111100_110_1_000011111100;
      patterns[34791] = 29'b1_000011111100_111_1_000011111100;
      patterns[34792] = 29'b1_000011111101_000_1_000011111101;
      patterns[34793] = 29'b1_000011111101_001_1_111101000011;
      patterns[34794] = 29'b1_000011111101_010_0_000111111011;
      patterns[34795] = 29'b1_000011111101_011_0_001111110110;
      patterns[34796] = 29'b1_000011111101_100_1_100001111110;
      patterns[34797] = 29'b1_000011111101_101_0_110000111111;
      patterns[34798] = 29'b1_000011111101_110_1_000011111101;
      patterns[34799] = 29'b1_000011111101_111_1_000011111101;
      patterns[34800] = 29'b1_000011111110_000_1_000011111110;
      patterns[34801] = 29'b1_000011111110_001_1_111110000011;
      patterns[34802] = 29'b1_000011111110_010_0_000111111101;
      patterns[34803] = 29'b1_000011111110_011_0_001111111010;
      patterns[34804] = 29'b1_000011111110_100_0_100001111111;
      patterns[34805] = 29'b1_000011111110_101_1_010000111111;
      patterns[34806] = 29'b1_000011111110_110_1_000011111110;
      patterns[34807] = 29'b1_000011111110_111_1_000011111110;
      patterns[34808] = 29'b1_000011111111_000_1_000011111111;
      patterns[34809] = 29'b1_000011111111_001_1_111111000011;
      patterns[34810] = 29'b1_000011111111_010_0_000111111111;
      patterns[34811] = 29'b1_000011111111_011_0_001111111110;
      patterns[34812] = 29'b1_000011111111_100_1_100001111111;
      patterns[34813] = 29'b1_000011111111_101_1_110000111111;
      patterns[34814] = 29'b1_000011111111_110_1_000011111111;
      patterns[34815] = 29'b1_000011111111_111_1_000011111111;
      patterns[34816] = 29'b1_000100000000_000_1_000100000000;
      patterns[34817] = 29'b1_000100000000_001_1_000000000100;
      patterns[34818] = 29'b1_000100000000_010_0_001000000001;
      patterns[34819] = 29'b1_000100000000_011_0_010000000010;
      patterns[34820] = 29'b1_000100000000_100_0_100010000000;
      patterns[34821] = 29'b1_000100000000_101_0_010001000000;
      patterns[34822] = 29'b1_000100000000_110_1_000100000000;
      patterns[34823] = 29'b1_000100000000_111_1_000100000000;
      patterns[34824] = 29'b1_000100000001_000_1_000100000001;
      patterns[34825] = 29'b1_000100000001_001_1_000001000100;
      patterns[34826] = 29'b1_000100000001_010_0_001000000011;
      patterns[34827] = 29'b1_000100000001_011_0_010000000110;
      patterns[34828] = 29'b1_000100000001_100_1_100010000000;
      patterns[34829] = 29'b1_000100000001_101_0_110001000000;
      patterns[34830] = 29'b1_000100000001_110_1_000100000001;
      patterns[34831] = 29'b1_000100000001_111_1_000100000001;
      patterns[34832] = 29'b1_000100000010_000_1_000100000010;
      patterns[34833] = 29'b1_000100000010_001_1_000010000100;
      patterns[34834] = 29'b1_000100000010_010_0_001000000101;
      patterns[34835] = 29'b1_000100000010_011_0_010000001010;
      patterns[34836] = 29'b1_000100000010_100_0_100010000001;
      patterns[34837] = 29'b1_000100000010_101_1_010001000000;
      patterns[34838] = 29'b1_000100000010_110_1_000100000010;
      patterns[34839] = 29'b1_000100000010_111_1_000100000010;
      patterns[34840] = 29'b1_000100000011_000_1_000100000011;
      patterns[34841] = 29'b1_000100000011_001_1_000011000100;
      patterns[34842] = 29'b1_000100000011_010_0_001000000111;
      patterns[34843] = 29'b1_000100000011_011_0_010000001110;
      patterns[34844] = 29'b1_000100000011_100_1_100010000001;
      patterns[34845] = 29'b1_000100000011_101_1_110001000000;
      patterns[34846] = 29'b1_000100000011_110_1_000100000011;
      patterns[34847] = 29'b1_000100000011_111_1_000100000011;
      patterns[34848] = 29'b1_000100000100_000_1_000100000100;
      patterns[34849] = 29'b1_000100000100_001_1_000100000100;
      patterns[34850] = 29'b1_000100000100_010_0_001000001001;
      patterns[34851] = 29'b1_000100000100_011_0_010000010010;
      patterns[34852] = 29'b1_000100000100_100_0_100010000010;
      patterns[34853] = 29'b1_000100000100_101_0_010001000001;
      patterns[34854] = 29'b1_000100000100_110_1_000100000100;
      patterns[34855] = 29'b1_000100000100_111_1_000100000100;
      patterns[34856] = 29'b1_000100000101_000_1_000100000101;
      patterns[34857] = 29'b1_000100000101_001_1_000101000100;
      patterns[34858] = 29'b1_000100000101_010_0_001000001011;
      patterns[34859] = 29'b1_000100000101_011_0_010000010110;
      patterns[34860] = 29'b1_000100000101_100_1_100010000010;
      patterns[34861] = 29'b1_000100000101_101_0_110001000001;
      patterns[34862] = 29'b1_000100000101_110_1_000100000101;
      patterns[34863] = 29'b1_000100000101_111_1_000100000101;
      patterns[34864] = 29'b1_000100000110_000_1_000100000110;
      patterns[34865] = 29'b1_000100000110_001_1_000110000100;
      patterns[34866] = 29'b1_000100000110_010_0_001000001101;
      patterns[34867] = 29'b1_000100000110_011_0_010000011010;
      patterns[34868] = 29'b1_000100000110_100_0_100010000011;
      patterns[34869] = 29'b1_000100000110_101_1_010001000001;
      patterns[34870] = 29'b1_000100000110_110_1_000100000110;
      patterns[34871] = 29'b1_000100000110_111_1_000100000110;
      patterns[34872] = 29'b1_000100000111_000_1_000100000111;
      patterns[34873] = 29'b1_000100000111_001_1_000111000100;
      patterns[34874] = 29'b1_000100000111_010_0_001000001111;
      patterns[34875] = 29'b1_000100000111_011_0_010000011110;
      patterns[34876] = 29'b1_000100000111_100_1_100010000011;
      patterns[34877] = 29'b1_000100000111_101_1_110001000001;
      patterns[34878] = 29'b1_000100000111_110_1_000100000111;
      patterns[34879] = 29'b1_000100000111_111_1_000100000111;
      patterns[34880] = 29'b1_000100001000_000_1_000100001000;
      patterns[34881] = 29'b1_000100001000_001_1_001000000100;
      patterns[34882] = 29'b1_000100001000_010_0_001000010001;
      patterns[34883] = 29'b1_000100001000_011_0_010000100010;
      patterns[34884] = 29'b1_000100001000_100_0_100010000100;
      patterns[34885] = 29'b1_000100001000_101_0_010001000010;
      patterns[34886] = 29'b1_000100001000_110_1_000100001000;
      patterns[34887] = 29'b1_000100001000_111_1_000100001000;
      patterns[34888] = 29'b1_000100001001_000_1_000100001001;
      patterns[34889] = 29'b1_000100001001_001_1_001001000100;
      patterns[34890] = 29'b1_000100001001_010_0_001000010011;
      patterns[34891] = 29'b1_000100001001_011_0_010000100110;
      patterns[34892] = 29'b1_000100001001_100_1_100010000100;
      patterns[34893] = 29'b1_000100001001_101_0_110001000010;
      patterns[34894] = 29'b1_000100001001_110_1_000100001001;
      patterns[34895] = 29'b1_000100001001_111_1_000100001001;
      patterns[34896] = 29'b1_000100001010_000_1_000100001010;
      patterns[34897] = 29'b1_000100001010_001_1_001010000100;
      patterns[34898] = 29'b1_000100001010_010_0_001000010101;
      patterns[34899] = 29'b1_000100001010_011_0_010000101010;
      patterns[34900] = 29'b1_000100001010_100_0_100010000101;
      patterns[34901] = 29'b1_000100001010_101_1_010001000010;
      patterns[34902] = 29'b1_000100001010_110_1_000100001010;
      patterns[34903] = 29'b1_000100001010_111_1_000100001010;
      patterns[34904] = 29'b1_000100001011_000_1_000100001011;
      patterns[34905] = 29'b1_000100001011_001_1_001011000100;
      patterns[34906] = 29'b1_000100001011_010_0_001000010111;
      patterns[34907] = 29'b1_000100001011_011_0_010000101110;
      patterns[34908] = 29'b1_000100001011_100_1_100010000101;
      patterns[34909] = 29'b1_000100001011_101_1_110001000010;
      patterns[34910] = 29'b1_000100001011_110_1_000100001011;
      patterns[34911] = 29'b1_000100001011_111_1_000100001011;
      patterns[34912] = 29'b1_000100001100_000_1_000100001100;
      patterns[34913] = 29'b1_000100001100_001_1_001100000100;
      patterns[34914] = 29'b1_000100001100_010_0_001000011001;
      patterns[34915] = 29'b1_000100001100_011_0_010000110010;
      patterns[34916] = 29'b1_000100001100_100_0_100010000110;
      patterns[34917] = 29'b1_000100001100_101_0_010001000011;
      patterns[34918] = 29'b1_000100001100_110_1_000100001100;
      patterns[34919] = 29'b1_000100001100_111_1_000100001100;
      patterns[34920] = 29'b1_000100001101_000_1_000100001101;
      patterns[34921] = 29'b1_000100001101_001_1_001101000100;
      patterns[34922] = 29'b1_000100001101_010_0_001000011011;
      patterns[34923] = 29'b1_000100001101_011_0_010000110110;
      patterns[34924] = 29'b1_000100001101_100_1_100010000110;
      patterns[34925] = 29'b1_000100001101_101_0_110001000011;
      patterns[34926] = 29'b1_000100001101_110_1_000100001101;
      patterns[34927] = 29'b1_000100001101_111_1_000100001101;
      patterns[34928] = 29'b1_000100001110_000_1_000100001110;
      patterns[34929] = 29'b1_000100001110_001_1_001110000100;
      patterns[34930] = 29'b1_000100001110_010_0_001000011101;
      patterns[34931] = 29'b1_000100001110_011_0_010000111010;
      patterns[34932] = 29'b1_000100001110_100_0_100010000111;
      patterns[34933] = 29'b1_000100001110_101_1_010001000011;
      patterns[34934] = 29'b1_000100001110_110_1_000100001110;
      patterns[34935] = 29'b1_000100001110_111_1_000100001110;
      patterns[34936] = 29'b1_000100001111_000_1_000100001111;
      patterns[34937] = 29'b1_000100001111_001_1_001111000100;
      patterns[34938] = 29'b1_000100001111_010_0_001000011111;
      patterns[34939] = 29'b1_000100001111_011_0_010000111110;
      patterns[34940] = 29'b1_000100001111_100_1_100010000111;
      patterns[34941] = 29'b1_000100001111_101_1_110001000011;
      patterns[34942] = 29'b1_000100001111_110_1_000100001111;
      patterns[34943] = 29'b1_000100001111_111_1_000100001111;
      patterns[34944] = 29'b1_000100010000_000_1_000100010000;
      patterns[34945] = 29'b1_000100010000_001_1_010000000100;
      patterns[34946] = 29'b1_000100010000_010_0_001000100001;
      patterns[34947] = 29'b1_000100010000_011_0_010001000010;
      patterns[34948] = 29'b1_000100010000_100_0_100010001000;
      patterns[34949] = 29'b1_000100010000_101_0_010001000100;
      patterns[34950] = 29'b1_000100010000_110_1_000100010000;
      patterns[34951] = 29'b1_000100010000_111_1_000100010000;
      patterns[34952] = 29'b1_000100010001_000_1_000100010001;
      patterns[34953] = 29'b1_000100010001_001_1_010001000100;
      patterns[34954] = 29'b1_000100010001_010_0_001000100011;
      patterns[34955] = 29'b1_000100010001_011_0_010001000110;
      patterns[34956] = 29'b1_000100010001_100_1_100010001000;
      patterns[34957] = 29'b1_000100010001_101_0_110001000100;
      patterns[34958] = 29'b1_000100010001_110_1_000100010001;
      patterns[34959] = 29'b1_000100010001_111_1_000100010001;
      patterns[34960] = 29'b1_000100010010_000_1_000100010010;
      patterns[34961] = 29'b1_000100010010_001_1_010010000100;
      patterns[34962] = 29'b1_000100010010_010_0_001000100101;
      patterns[34963] = 29'b1_000100010010_011_0_010001001010;
      patterns[34964] = 29'b1_000100010010_100_0_100010001001;
      patterns[34965] = 29'b1_000100010010_101_1_010001000100;
      patterns[34966] = 29'b1_000100010010_110_1_000100010010;
      patterns[34967] = 29'b1_000100010010_111_1_000100010010;
      patterns[34968] = 29'b1_000100010011_000_1_000100010011;
      patterns[34969] = 29'b1_000100010011_001_1_010011000100;
      patterns[34970] = 29'b1_000100010011_010_0_001000100111;
      patterns[34971] = 29'b1_000100010011_011_0_010001001110;
      patterns[34972] = 29'b1_000100010011_100_1_100010001001;
      patterns[34973] = 29'b1_000100010011_101_1_110001000100;
      patterns[34974] = 29'b1_000100010011_110_1_000100010011;
      patterns[34975] = 29'b1_000100010011_111_1_000100010011;
      patterns[34976] = 29'b1_000100010100_000_1_000100010100;
      patterns[34977] = 29'b1_000100010100_001_1_010100000100;
      patterns[34978] = 29'b1_000100010100_010_0_001000101001;
      patterns[34979] = 29'b1_000100010100_011_0_010001010010;
      patterns[34980] = 29'b1_000100010100_100_0_100010001010;
      patterns[34981] = 29'b1_000100010100_101_0_010001000101;
      patterns[34982] = 29'b1_000100010100_110_1_000100010100;
      patterns[34983] = 29'b1_000100010100_111_1_000100010100;
      patterns[34984] = 29'b1_000100010101_000_1_000100010101;
      patterns[34985] = 29'b1_000100010101_001_1_010101000100;
      patterns[34986] = 29'b1_000100010101_010_0_001000101011;
      patterns[34987] = 29'b1_000100010101_011_0_010001010110;
      patterns[34988] = 29'b1_000100010101_100_1_100010001010;
      patterns[34989] = 29'b1_000100010101_101_0_110001000101;
      patterns[34990] = 29'b1_000100010101_110_1_000100010101;
      patterns[34991] = 29'b1_000100010101_111_1_000100010101;
      patterns[34992] = 29'b1_000100010110_000_1_000100010110;
      patterns[34993] = 29'b1_000100010110_001_1_010110000100;
      patterns[34994] = 29'b1_000100010110_010_0_001000101101;
      patterns[34995] = 29'b1_000100010110_011_0_010001011010;
      patterns[34996] = 29'b1_000100010110_100_0_100010001011;
      patterns[34997] = 29'b1_000100010110_101_1_010001000101;
      patterns[34998] = 29'b1_000100010110_110_1_000100010110;
      patterns[34999] = 29'b1_000100010110_111_1_000100010110;
      patterns[35000] = 29'b1_000100010111_000_1_000100010111;
      patterns[35001] = 29'b1_000100010111_001_1_010111000100;
      patterns[35002] = 29'b1_000100010111_010_0_001000101111;
      patterns[35003] = 29'b1_000100010111_011_0_010001011110;
      patterns[35004] = 29'b1_000100010111_100_1_100010001011;
      patterns[35005] = 29'b1_000100010111_101_1_110001000101;
      patterns[35006] = 29'b1_000100010111_110_1_000100010111;
      patterns[35007] = 29'b1_000100010111_111_1_000100010111;
      patterns[35008] = 29'b1_000100011000_000_1_000100011000;
      patterns[35009] = 29'b1_000100011000_001_1_011000000100;
      patterns[35010] = 29'b1_000100011000_010_0_001000110001;
      patterns[35011] = 29'b1_000100011000_011_0_010001100010;
      patterns[35012] = 29'b1_000100011000_100_0_100010001100;
      patterns[35013] = 29'b1_000100011000_101_0_010001000110;
      patterns[35014] = 29'b1_000100011000_110_1_000100011000;
      patterns[35015] = 29'b1_000100011000_111_1_000100011000;
      patterns[35016] = 29'b1_000100011001_000_1_000100011001;
      patterns[35017] = 29'b1_000100011001_001_1_011001000100;
      patterns[35018] = 29'b1_000100011001_010_0_001000110011;
      patterns[35019] = 29'b1_000100011001_011_0_010001100110;
      patterns[35020] = 29'b1_000100011001_100_1_100010001100;
      patterns[35021] = 29'b1_000100011001_101_0_110001000110;
      patterns[35022] = 29'b1_000100011001_110_1_000100011001;
      patterns[35023] = 29'b1_000100011001_111_1_000100011001;
      patterns[35024] = 29'b1_000100011010_000_1_000100011010;
      patterns[35025] = 29'b1_000100011010_001_1_011010000100;
      patterns[35026] = 29'b1_000100011010_010_0_001000110101;
      patterns[35027] = 29'b1_000100011010_011_0_010001101010;
      patterns[35028] = 29'b1_000100011010_100_0_100010001101;
      patterns[35029] = 29'b1_000100011010_101_1_010001000110;
      patterns[35030] = 29'b1_000100011010_110_1_000100011010;
      patterns[35031] = 29'b1_000100011010_111_1_000100011010;
      patterns[35032] = 29'b1_000100011011_000_1_000100011011;
      patterns[35033] = 29'b1_000100011011_001_1_011011000100;
      patterns[35034] = 29'b1_000100011011_010_0_001000110111;
      patterns[35035] = 29'b1_000100011011_011_0_010001101110;
      patterns[35036] = 29'b1_000100011011_100_1_100010001101;
      patterns[35037] = 29'b1_000100011011_101_1_110001000110;
      patterns[35038] = 29'b1_000100011011_110_1_000100011011;
      patterns[35039] = 29'b1_000100011011_111_1_000100011011;
      patterns[35040] = 29'b1_000100011100_000_1_000100011100;
      patterns[35041] = 29'b1_000100011100_001_1_011100000100;
      patterns[35042] = 29'b1_000100011100_010_0_001000111001;
      patterns[35043] = 29'b1_000100011100_011_0_010001110010;
      patterns[35044] = 29'b1_000100011100_100_0_100010001110;
      patterns[35045] = 29'b1_000100011100_101_0_010001000111;
      patterns[35046] = 29'b1_000100011100_110_1_000100011100;
      patterns[35047] = 29'b1_000100011100_111_1_000100011100;
      patterns[35048] = 29'b1_000100011101_000_1_000100011101;
      patterns[35049] = 29'b1_000100011101_001_1_011101000100;
      patterns[35050] = 29'b1_000100011101_010_0_001000111011;
      patterns[35051] = 29'b1_000100011101_011_0_010001110110;
      patterns[35052] = 29'b1_000100011101_100_1_100010001110;
      patterns[35053] = 29'b1_000100011101_101_0_110001000111;
      patterns[35054] = 29'b1_000100011101_110_1_000100011101;
      patterns[35055] = 29'b1_000100011101_111_1_000100011101;
      patterns[35056] = 29'b1_000100011110_000_1_000100011110;
      patterns[35057] = 29'b1_000100011110_001_1_011110000100;
      patterns[35058] = 29'b1_000100011110_010_0_001000111101;
      patterns[35059] = 29'b1_000100011110_011_0_010001111010;
      patterns[35060] = 29'b1_000100011110_100_0_100010001111;
      patterns[35061] = 29'b1_000100011110_101_1_010001000111;
      patterns[35062] = 29'b1_000100011110_110_1_000100011110;
      patterns[35063] = 29'b1_000100011110_111_1_000100011110;
      patterns[35064] = 29'b1_000100011111_000_1_000100011111;
      patterns[35065] = 29'b1_000100011111_001_1_011111000100;
      patterns[35066] = 29'b1_000100011111_010_0_001000111111;
      patterns[35067] = 29'b1_000100011111_011_0_010001111110;
      patterns[35068] = 29'b1_000100011111_100_1_100010001111;
      patterns[35069] = 29'b1_000100011111_101_1_110001000111;
      patterns[35070] = 29'b1_000100011111_110_1_000100011111;
      patterns[35071] = 29'b1_000100011111_111_1_000100011111;
      patterns[35072] = 29'b1_000100100000_000_1_000100100000;
      patterns[35073] = 29'b1_000100100000_001_1_100000000100;
      patterns[35074] = 29'b1_000100100000_010_0_001001000001;
      patterns[35075] = 29'b1_000100100000_011_0_010010000010;
      patterns[35076] = 29'b1_000100100000_100_0_100010010000;
      patterns[35077] = 29'b1_000100100000_101_0_010001001000;
      patterns[35078] = 29'b1_000100100000_110_1_000100100000;
      patterns[35079] = 29'b1_000100100000_111_1_000100100000;
      patterns[35080] = 29'b1_000100100001_000_1_000100100001;
      patterns[35081] = 29'b1_000100100001_001_1_100001000100;
      patterns[35082] = 29'b1_000100100001_010_0_001001000011;
      patterns[35083] = 29'b1_000100100001_011_0_010010000110;
      patterns[35084] = 29'b1_000100100001_100_1_100010010000;
      patterns[35085] = 29'b1_000100100001_101_0_110001001000;
      patterns[35086] = 29'b1_000100100001_110_1_000100100001;
      patterns[35087] = 29'b1_000100100001_111_1_000100100001;
      patterns[35088] = 29'b1_000100100010_000_1_000100100010;
      patterns[35089] = 29'b1_000100100010_001_1_100010000100;
      patterns[35090] = 29'b1_000100100010_010_0_001001000101;
      patterns[35091] = 29'b1_000100100010_011_0_010010001010;
      patterns[35092] = 29'b1_000100100010_100_0_100010010001;
      patterns[35093] = 29'b1_000100100010_101_1_010001001000;
      patterns[35094] = 29'b1_000100100010_110_1_000100100010;
      patterns[35095] = 29'b1_000100100010_111_1_000100100010;
      patterns[35096] = 29'b1_000100100011_000_1_000100100011;
      patterns[35097] = 29'b1_000100100011_001_1_100011000100;
      patterns[35098] = 29'b1_000100100011_010_0_001001000111;
      patterns[35099] = 29'b1_000100100011_011_0_010010001110;
      patterns[35100] = 29'b1_000100100011_100_1_100010010001;
      patterns[35101] = 29'b1_000100100011_101_1_110001001000;
      patterns[35102] = 29'b1_000100100011_110_1_000100100011;
      patterns[35103] = 29'b1_000100100011_111_1_000100100011;
      patterns[35104] = 29'b1_000100100100_000_1_000100100100;
      patterns[35105] = 29'b1_000100100100_001_1_100100000100;
      patterns[35106] = 29'b1_000100100100_010_0_001001001001;
      patterns[35107] = 29'b1_000100100100_011_0_010010010010;
      patterns[35108] = 29'b1_000100100100_100_0_100010010010;
      patterns[35109] = 29'b1_000100100100_101_0_010001001001;
      patterns[35110] = 29'b1_000100100100_110_1_000100100100;
      patterns[35111] = 29'b1_000100100100_111_1_000100100100;
      patterns[35112] = 29'b1_000100100101_000_1_000100100101;
      patterns[35113] = 29'b1_000100100101_001_1_100101000100;
      patterns[35114] = 29'b1_000100100101_010_0_001001001011;
      patterns[35115] = 29'b1_000100100101_011_0_010010010110;
      patterns[35116] = 29'b1_000100100101_100_1_100010010010;
      patterns[35117] = 29'b1_000100100101_101_0_110001001001;
      patterns[35118] = 29'b1_000100100101_110_1_000100100101;
      patterns[35119] = 29'b1_000100100101_111_1_000100100101;
      patterns[35120] = 29'b1_000100100110_000_1_000100100110;
      patterns[35121] = 29'b1_000100100110_001_1_100110000100;
      patterns[35122] = 29'b1_000100100110_010_0_001001001101;
      patterns[35123] = 29'b1_000100100110_011_0_010010011010;
      patterns[35124] = 29'b1_000100100110_100_0_100010010011;
      patterns[35125] = 29'b1_000100100110_101_1_010001001001;
      patterns[35126] = 29'b1_000100100110_110_1_000100100110;
      patterns[35127] = 29'b1_000100100110_111_1_000100100110;
      patterns[35128] = 29'b1_000100100111_000_1_000100100111;
      patterns[35129] = 29'b1_000100100111_001_1_100111000100;
      patterns[35130] = 29'b1_000100100111_010_0_001001001111;
      patterns[35131] = 29'b1_000100100111_011_0_010010011110;
      patterns[35132] = 29'b1_000100100111_100_1_100010010011;
      patterns[35133] = 29'b1_000100100111_101_1_110001001001;
      patterns[35134] = 29'b1_000100100111_110_1_000100100111;
      patterns[35135] = 29'b1_000100100111_111_1_000100100111;
      patterns[35136] = 29'b1_000100101000_000_1_000100101000;
      patterns[35137] = 29'b1_000100101000_001_1_101000000100;
      patterns[35138] = 29'b1_000100101000_010_0_001001010001;
      patterns[35139] = 29'b1_000100101000_011_0_010010100010;
      patterns[35140] = 29'b1_000100101000_100_0_100010010100;
      patterns[35141] = 29'b1_000100101000_101_0_010001001010;
      patterns[35142] = 29'b1_000100101000_110_1_000100101000;
      patterns[35143] = 29'b1_000100101000_111_1_000100101000;
      patterns[35144] = 29'b1_000100101001_000_1_000100101001;
      patterns[35145] = 29'b1_000100101001_001_1_101001000100;
      patterns[35146] = 29'b1_000100101001_010_0_001001010011;
      patterns[35147] = 29'b1_000100101001_011_0_010010100110;
      patterns[35148] = 29'b1_000100101001_100_1_100010010100;
      patterns[35149] = 29'b1_000100101001_101_0_110001001010;
      patterns[35150] = 29'b1_000100101001_110_1_000100101001;
      patterns[35151] = 29'b1_000100101001_111_1_000100101001;
      patterns[35152] = 29'b1_000100101010_000_1_000100101010;
      patterns[35153] = 29'b1_000100101010_001_1_101010000100;
      patterns[35154] = 29'b1_000100101010_010_0_001001010101;
      patterns[35155] = 29'b1_000100101010_011_0_010010101010;
      patterns[35156] = 29'b1_000100101010_100_0_100010010101;
      patterns[35157] = 29'b1_000100101010_101_1_010001001010;
      patterns[35158] = 29'b1_000100101010_110_1_000100101010;
      patterns[35159] = 29'b1_000100101010_111_1_000100101010;
      patterns[35160] = 29'b1_000100101011_000_1_000100101011;
      patterns[35161] = 29'b1_000100101011_001_1_101011000100;
      patterns[35162] = 29'b1_000100101011_010_0_001001010111;
      patterns[35163] = 29'b1_000100101011_011_0_010010101110;
      patterns[35164] = 29'b1_000100101011_100_1_100010010101;
      patterns[35165] = 29'b1_000100101011_101_1_110001001010;
      patterns[35166] = 29'b1_000100101011_110_1_000100101011;
      patterns[35167] = 29'b1_000100101011_111_1_000100101011;
      patterns[35168] = 29'b1_000100101100_000_1_000100101100;
      patterns[35169] = 29'b1_000100101100_001_1_101100000100;
      patterns[35170] = 29'b1_000100101100_010_0_001001011001;
      patterns[35171] = 29'b1_000100101100_011_0_010010110010;
      patterns[35172] = 29'b1_000100101100_100_0_100010010110;
      patterns[35173] = 29'b1_000100101100_101_0_010001001011;
      patterns[35174] = 29'b1_000100101100_110_1_000100101100;
      patterns[35175] = 29'b1_000100101100_111_1_000100101100;
      patterns[35176] = 29'b1_000100101101_000_1_000100101101;
      patterns[35177] = 29'b1_000100101101_001_1_101101000100;
      patterns[35178] = 29'b1_000100101101_010_0_001001011011;
      patterns[35179] = 29'b1_000100101101_011_0_010010110110;
      patterns[35180] = 29'b1_000100101101_100_1_100010010110;
      patterns[35181] = 29'b1_000100101101_101_0_110001001011;
      patterns[35182] = 29'b1_000100101101_110_1_000100101101;
      patterns[35183] = 29'b1_000100101101_111_1_000100101101;
      patterns[35184] = 29'b1_000100101110_000_1_000100101110;
      patterns[35185] = 29'b1_000100101110_001_1_101110000100;
      patterns[35186] = 29'b1_000100101110_010_0_001001011101;
      patterns[35187] = 29'b1_000100101110_011_0_010010111010;
      patterns[35188] = 29'b1_000100101110_100_0_100010010111;
      patterns[35189] = 29'b1_000100101110_101_1_010001001011;
      patterns[35190] = 29'b1_000100101110_110_1_000100101110;
      patterns[35191] = 29'b1_000100101110_111_1_000100101110;
      patterns[35192] = 29'b1_000100101111_000_1_000100101111;
      patterns[35193] = 29'b1_000100101111_001_1_101111000100;
      patterns[35194] = 29'b1_000100101111_010_0_001001011111;
      patterns[35195] = 29'b1_000100101111_011_0_010010111110;
      patterns[35196] = 29'b1_000100101111_100_1_100010010111;
      patterns[35197] = 29'b1_000100101111_101_1_110001001011;
      patterns[35198] = 29'b1_000100101111_110_1_000100101111;
      patterns[35199] = 29'b1_000100101111_111_1_000100101111;
      patterns[35200] = 29'b1_000100110000_000_1_000100110000;
      patterns[35201] = 29'b1_000100110000_001_1_110000000100;
      patterns[35202] = 29'b1_000100110000_010_0_001001100001;
      patterns[35203] = 29'b1_000100110000_011_0_010011000010;
      patterns[35204] = 29'b1_000100110000_100_0_100010011000;
      patterns[35205] = 29'b1_000100110000_101_0_010001001100;
      patterns[35206] = 29'b1_000100110000_110_1_000100110000;
      patterns[35207] = 29'b1_000100110000_111_1_000100110000;
      patterns[35208] = 29'b1_000100110001_000_1_000100110001;
      patterns[35209] = 29'b1_000100110001_001_1_110001000100;
      patterns[35210] = 29'b1_000100110001_010_0_001001100011;
      patterns[35211] = 29'b1_000100110001_011_0_010011000110;
      patterns[35212] = 29'b1_000100110001_100_1_100010011000;
      patterns[35213] = 29'b1_000100110001_101_0_110001001100;
      patterns[35214] = 29'b1_000100110001_110_1_000100110001;
      patterns[35215] = 29'b1_000100110001_111_1_000100110001;
      patterns[35216] = 29'b1_000100110010_000_1_000100110010;
      patterns[35217] = 29'b1_000100110010_001_1_110010000100;
      patterns[35218] = 29'b1_000100110010_010_0_001001100101;
      patterns[35219] = 29'b1_000100110010_011_0_010011001010;
      patterns[35220] = 29'b1_000100110010_100_0_100010011001;
      patterns[35221] = 29'b1_000100110010_101_1_010001001100;
      patterns[35222] = 29'b1_000100110010_110_1_000100110010;
      patterns[35223] = 29'b1_000100110010_111_1_000100110010;
      patterns[35224] = 29'b1_000100110011_000_1_000100110011;
      patterns[35225] = 29'b1_000100110011_001_1_110011000100;
      patterns[35226] = 29'b1_000100110011_010_0_001001100111;
      patterns[35227] = 29'b1_000100110011_011_0_010011001110;
      patterns[35228] = 29'b1_000100110011_100_1_100010011001;
      patterns[35229] = 29'b1_000100110011_101_1_110001001100;
      patterns[35230] = 29'b1_000100110011_110_1_000100110011;
      patterns[35231] = 29'b1_000100110011_111_1_000100110011;
      patterns[35232] = 29'b1_000100110100_000_1_000100110100;
      patterns[35233] = 29'b1_000100110100_001_1_110100000100;
      patterns[35234] = 29'b1_000100110100_010_0_001001101001;
      patterns[35235] = 29'b1_000100110100_011_0_010011010010;
      patterns[35236] = 29'b1_000100110100_100_0_100010011010;
      patterns[35237] = 29'b1_000100110100_101_0_010001001101;
      patterns[35238] = 29'b1_000100110100_110_1_000100110100;
      patterns[35239] = 29'b1_000100110100_111_1_000100110100;
      patterns[35240] = 29'b1_000100110101_000_1_000100110101;
      patterns[35241] = 29'b1_000100110101_001_1_110101000100;
      patterns[35242] = 29'b1_000100110101_010_0_001001101011;
      patterns[35243] = 29'b1_000100110101_011_0_010011010110;
      patterns[35244] = 29'b1_000100110101_100_1_100010011010;
      patterns[35245] = 29'b1_000100110101_101_0_110001001101;
      patterns[35246] = 29'b1_000100110101_110_1_000100110101;
      patterns[35247] = 29'b1_000100110101_111_1_000100110101;
      patterns[35248] = 29'b1_000100110110_000_1_000100110110;
      patterns[35249] = 29'b1_000100110110_001_1_110110000100;
      patterns[35250] = 29'b1_000100110110_010_0_001001101101;
      patterns[35251] = 29'b1_000100110110_011_0_010011011010;
      patterns[35252] = 29'b1_000100110110_100_0_100010011011;
      patterns[35253] = 29'b1_000100110110_101_1_010001001101;
      patterns[35254] = 29'b1_000100110110_110_1_000100110110;
      patterns[35255] = 29'b1_000100110110_111_1_000100110110;
      patterns[35256] = 29'b1_000100110111_000_1_000100110111;
      patterns[35257] = 29'b1_000100110111_001_1_110111000100;
      patterns[35258] = 29'b1_000100110111_010_0_001001101111;
      patterns[35259] = 29'b1_000100110111_011_0_010011011110;
      patterns[35260] = 29'b1_000100110111_100_1_100010011011;
      patterns[35261] = 29'b1_000100110111_101_1_110001001101;
      patterns[35262] = 29'b1_000100110111_110_1_000100110111;
      patterns[35263] = 29'b1_000100110111_111_1_000100110111;
      patterns[35264] = 29'b1_000100111000_000_1_000100111000;
      patterns[35265] = 29'b1_000100111000_001_1_111000000100;
      patterns[35266] = 29'b1_000100111000_010_0_001001110001;
      patterns[35267] = 29'b1_000100111000_011_0_010011100010;
      patterns[35268] = 29'b1_000100111000_100_0_100010011100;
      patterns[35269] = 29'b1_000100111000_101_0_010001001110;
      patterns[35270] = 29'b1_000100111000_110_1_000100111000;
      patterns[35271] = 29'b1_000100111000_111_1_000100111000;
      patterns[35272] = 29'b1_000100111001_000_1_000100111001;
      patterns[35273] = 29'b1_000100111001_001_1_111001000100;
      patterns[35274] = 29'b1_000100111001_010_0_001001110011;
      patterns[35275] = 29'b1_000100111001_011_0_010011100110;
      patterns[35276] = 29'b1_000100111001_100_1_100010011100;
      patterns[35277] = 29'b1_000100111001_101_0_110001001110;
      patterns[35278] = 29'b1_000100111001_110_1_000100111001;
      patterns[35279] = 29'b1_000100111001_111_1_000100111001;
      patterns[35280] = 29'b1_000100111010_000_1_000100111010;
      patterns[35281] = 29'b1_000100111010_001_1_111010000100;
      patterns[35282] = 29'b1_000100111010_010_0_001001110101;
      patterns[35283] = 29'b1_000100111010_011_0_010011101010;
      patterns[35284] = 29'b1_000100111010_100_0_100010011101;
      patterns[35285] = 29'b1_000100111010_101_1_010001001110;
      patterns[35286] = 29'b1_000100111010_110_1_000100111010;
      patterns[35287] = 29'b1_000100111010_111_1_000100111010;
      patterns[35288] = 29'b1_000100111011_000_1_000100111011;
      patterns[35289] = 29'b1_000100111011_001_1_111011000100;
      patterns[35290] = 29'b1_000100111011_010_0_001001110111;
      patterns[35291] = 29'b1_000100111011_011_0_010011101110;
      patterns[35292] = 29'b1_000100111011_100_1_100010011101;
      patterns[35293] = 29'b1_000100111011_101_1_110001001110;
      patterns[35294] = 29'b1_000100111011_110_1_000100111011;
      patterns[35295] = 29'b1_000100111011_111_1_000100111011;
      patterns[35296] = 29'b1_000100111100_000_1_000100111100;
      patterns[35297] = 29'b1_000100111100_001_1_111100000100;
      patterns[35298] = 29'b1_000100111100_010_0_001001111001;
      patterns[35299] = 29'b1_000100111100_011_0_010011110010;
      patterns[35300] = 29'b1_000100111100_100_0_100010011110;
      patterns[35301] = 29'b1_000100111100_101_0_010001001111;
      patterns[35302] = 29'b1_000100111100_110_1_000100111100;
      patterns[35303] = 29'b1_000100111100_111_1_000100111100;
      patterns[35304] = 29'b1_000100111101_000_1_000100111101;
      patterns[35305] = 29'b1_000100111101_001_1_111101000100;
      patterns[35306] = 29'b1_000100111101_010_0_001001111011;
      patterns[35307] = 29'b1_000100111101_011_0_010011110110;
      patterns[35308] = 29'b1_000100111101_100_1_100010011110;
      patterns[35309] = 29'b1_000100111101_101_0_110001001111;
      patterns[35310] = 29'b1_000100111101_110_1_000100111101;
      patterns[35311] = 29'b1_000100111101_111_1_000100111101;
      patterns[35312] = 29'b1_000100111110_000_1_000100111110;
      patterns[35313] = 29'b1_000100111110_001_1_111110000100;
      patterns[35314] = 29'b1_000100111110_010_0_001001111101;
      patterns[35315] = 29'b1_000100111110_011_0_010011111010;
      patterns[35316] = 29'b1_000100111110_100_0_100010011111;
      patterns[35317] = 29'b1_000100111110_101_1_010001001111;
      patterns[35318] = 29'b1_000100111110_110_1_000100111110;
      patterns[35319] = 29'b1_000100111110_111_1_000100111110;
      patterns[35320] = 29'b1_000100111111_000_1_000100111111;
      patterns[35321] = 29'b1_000100111111_001_1_111111000100;
      patterns[35322] = 29'b1_000100111111_010_0_001001111111;
      patterns[35323] = 29'b1_000100111111_011_0_010011111110;
      patterns[35324] = 29'b1_000100111111_100_1_100010011111;
      patterns[35325] = 29'b1_000100111111_101_1_110001001111;
      patterns[35326] = 29'b1_000100111111_110_1_000100111111;
      patterns[35327] = 29'b1_000100111111_111_1_000100111111;
      patterns[35328] = 29'b1_000101000000_000_1_000101000000;
      patterns[35329] = 29'b1_000101000000_001_1_000000000101;
      patterns[35330] = 29'b1_000101000000_010_0_001010000001;
      patterns[35331] = 29'b1_000101000000_011_0_010100000010;
      patterns[35332] = 29'b1_000101000000_100_0_100010100000;
      patterns[35333] = 29'b1_000101000000_101_0_010001010000;
      patterns[35334] = 29'b1_000101000000_110_1_000101000000;
      patterns[35335] = 29'b1_000101000000_111_1_000101000000;
      patterns[35336] = 29'b1_000101000001_000_1_000101000001;
      patterns[35337] = 29'b1_000101000001_001_1_000001000101;
      patterns[35338] = 29'b1_000101000001_010_0_001010000011;
      patterns[35339] = 29'b1_000101000001_011_0_010100000110;
      patterns[35340] = 29'b1_000101000001_100_1_100010100000;
      patterns[35341] = 29'b1_000101000001_101_0_110001010000;
      patterns[35342] = 29'b1_000101000001_110_1_000101000001;
      patterns[35343] = 29'b1_000101000001_111_1_000101000001;
      patterns[35344] = 29'b1_000101000010_000_1_000101000010;
      patterns[35345] = 29'b1_000101000010_001_1_000010000101;
      patterns[35346] = 29'b1_000101000010_010_0_001010000101;
      patterns[35347] = 29'b1_000101000010_011_0_010100001010;
      patterns[35348] = 29'b1_000101000010_100_0_100010100001;
      patterns[35349] = 29'b1_000101000010_101_1_010001010000;
      patterns[35350] = 29'b1_000101000010_110_1_000101000010;
      patterns[35351] = 29'b1_000101000010_111_1_000101000010;
      patterns[35352] = 29'b1_000101000011_000_1_000101000011;
      patterns[35353] = 29'b1_000101000011_001_1_000011000101;
      patterns[35354] = 29'b1_000101000011_010_0_001010000111;
      patterns[35355] = 29'b1_000101000011_011_0_010100001110;
      patterns[35356] = 29'b1_000101000011_100_1_100010100001;
      patterns[35357] = 29'b1_000101000011_101_1_110001010000;
      patterns[35358] = 29'b1_000101000011_110_1_000101000011;
      patterns[35359] = 29'b1_000101000011_111_1_000101000011;
      patterns[35360] = 29'b1_000101000100_000_1_000101000100;
      patterns[35361] = 29'b1_000101000100_001_1_000100000101;
      patterns[35362] = 29'b1_000101000100_010_0_001010001001;
      patterns[35363] = 29'b1_000101000100_011_0_010100010010;
      patterns[35364] = 29'b1_000101000100_100_0_100010100010;
      patterns[35365] = 29'b1_000101000100_101_0_010001010001;
      patterns[35366] = 29'b1_000101000100_110_1_000101000100;
      patterns[35367] = 29'b1_000101000100_111_1_000101000100;
      patterns[35368] = 29'b1_000101000101_000_1_000101000101;
      patterns[35369] = 29'b1_000101000101_001_1_000101000101;
      patterns[35370] = 29'b1_000101000101_010_0_001010001011;
      patterns[35371] = 29'b1_000101000101_011_0_010100010110;
      patterns[35372] = 29'b1_000101000101_100_1_100010100010;
      patterns[35373] = 29'b1_000101000101_101_0_110001010001;
      patterns[35374] = 29'b1_000101000101_110_1_000101000101;
      patterns[35375] = 29'b1_000101000101_111_1_000101000101;
      patterns[35376] = 29'b1_000101000110_000_1_000101000110;
      patterns[35377] = 29'b1_000101000110_001_1_000110000101;
      patterns[35378] = 29'b1_000101000110_010_0_001010001101;
      patterns[35379] = 29'b1_000101000110_011_0_010100011010;
      patterns[35380] = 29'b1_000101000110_100_0_100010100011;
      patterns[35381] = 29'b1_000101000110_101_1_010001010001;
      patterns[35382] = 29'b1_000101000110_110_1_000101000110;
      patterns[35383] = 29'b1_000101000110_111_1_000101000110;
      patterns[35384] = 29'b1_000101000111_000_1_000101000111;
      patterns[35385] = 29'b1_000101000111_001_1_000111000101;
      patterns[35386] = 29'b1_000101000111_010_0_001010001111;
      patterns[35387] = 29'b1_000101000111_011_0_010100011110;
      patterns[35388] = 29'b1_000101000111_100_1_100010100011;
      patterns[35389] = 29'b1_000101000111_101_1_110001010001;
      patterns[35390] = 29'b1_000101000111_110_1_000101000111;
      patterns[35391] = 29'b1_000101000111_111_1_000101000111;
      patterns[35392] = 29'b1_000101001000_000_1_000101001000;
      patterns[35393] = 29'b1_000101001000_001_1_001000000101;
      patterns[35394] = 29'b1_000101001000_010_0_001010010001;
      patterns[35395] = 29'b1_000101001000_011_0_010100100010;
      patterns[35396] = 29'b1_000101001000_100_0_100010100100;
      patterns[35397] = 29'b1_000101001000_101_0_010001010010;
      patterns[35398] = 29'b1_000101001000_110_1_000101001000;
      patterns[35399] = 29'b1_000101001000_111_1_000101001000;
      patterns[35400] = 29'b1_000101001001_000_1_000101001001;
      patterns[35401] = 29'b1_000101001001_001_1_001001000101;
      patterns[35402] = 29'b1_000101001001_010_0_001010010011;
      patterns[35403] = 29'b1_000101001001_011_0_010100100110;
      patterns[35404] = 29'b1_000101001001_100_1_100010100100;
      patterns[35405] = 29'b1_000101001001_101_0_110001010010;
      patterns[35406] = 29'b1_000101001001_110_1_000101001001;
      patterns[35407] = 29'b1_000101001001_111_1_000101001001;
      patterns[35408] = 29'b1_000101001010_000_1_000101001010;
      patterns[35409] = 29'b1_000101001010_001_1_001010000101;
      patterns[35410] = 29'b1_000101001010_010_0_001010010101;
      patterns[35411] = 29'b1_000101001010_011_0_010100101010;
      patterns[35412] = 29'b1_000101001010_100_0_100010100101;
      patterns[35413] = 29'b1_000101001010_101_1_010001010010;
      patterns[35414] = 29'b1_000101001010_110_1_000101001010;
      patterns[35415] = 29'b1_000101001010_111_1_000101001010;
      patterns[35416] = 29'b1_000101001011_000_1_000101001011;
      patterns[35417] = 29'b1_000101001011_001_1_001011000101;
      patterns[35418] = 29'b1_000101001011_010_0_001010010111;
      patterns[35419] = 29'b1_000101001011_011_0_010100101110;
      patterns[35420] = 29'b1_000101001011_100_1_100010100101;
      patterns[35421] = 29'b1_000101001011_101_1_110001010010;
      patterns[35422] = 29'b1_000101001011_110_1_000101001011;
      patterns[35423] = 29'b1_000101001011_111_1_000101001011;
      patterns[35424] = 29'b1_000101001100_000_1_000101001100;
      patterns[35425] = 29'b1_000101001100_001_1_001100000101;
      patterns[35426] = 29'b1_000101001100_010_0_001010011001;
      patterns[35427] = 29'b1_000101001100_011_0_010100110010;
      patterns[35428] = 29'b1_000101001100_100_0_100010100110;
      patterns[35429] = 29'b1_000101001100_101_0_010001010011;
      patterns[35430] = 29'b1_000101001100_110_1_000101001100;
      patterns[35431] = 29'b1_000101001100_111_1_000101001100;
      patterns[35432] = 29'b1_000101001101_000_1_000101001101;
      patterns[35433] = 29'b1_000101001101_001_1_001101000101;
      patterns[35434] = 29'b1_000101001101_010_0_001010011011;
      patterns[35435] = 29'b1_000101001101_011_0_010100110110;
      patterns[35436] = 29'b1_000101001101_100_1_100010100110;
      patterns[35437] = 29'b1_000101001101_101_0_110001010011;
      patterns[35438] = 29'b1_000101001101_110_1_000101001101;
      patterns[35439] = 29'b1_000101001101_111_1_000101001101;
      patterns[35440] = 29'b1_000101001110_000_1_000101001110;
      patterns[35441] = 29'b1_000101001110_001_1_001110000101;
      patterns[35442] = 29'b1_000101001110_010_0_001010011101;
      patterns[35443] = 29'b1_000101001110_011_0_010100111010;
      patterns[35444] = 29'b1_000101001110_100_0_100010100111;
      patterns[35445] = 29'b1_000101001110_101_1_010001010011;
      patterns[35446] = 29'b1_000101001110_110_1_000101001110;
      patterns[35447] = 29'b1_000101001110_111_1_000101001110;
      patterns[35448] = 29'b1_000101001111_000_1_000101001111;
      patterns[35449] = 29'b1_000101001111_001_1_001111000101;
      patterns[35450] = 29'b1_000101001111_010_0_001010011111;
      patterns[35451] = 29'b1_000101001111_011_0_010100111110;
      patterns[35452] = 29'b1_000101001111_100_1_100010100111;
      patterns[35453] = 29'b1_000101001111_101_1_110001010011;
      patterns[35454] = 29'b1_000101001111_110_1_000101001111;
      patterns[35455] = 29'b1_000101001111_111_1_000101001111;
      patterns[35456] = 29'b1_000101010000_000_1_000101010000;
      patterns[35457] = 29'b1_000101010000_001_1_010000000101;
      patterns[35458] = 29'b1_000101010000_010_0_001010100001;
      patterns[35459] = 29'b1_000101010000_011_0_010101000010;
      patterns[35460] = 29'b1_000101010000_100_0_100010101000;
      patterns[35461] = 29'b1_000101010000_101_0_010001010100;
      patterns[35462] = 29'b1_000101010000_110_1_000101010000;
      patterns[35463] = 29'b1_000101010000_111_1_000101010000;
      patterns[35464] = 29'b1_000101010001_000_1_000101010001;
      patterns[35465] = 29'b1_000101010001_001_1_010001000101;
      patterns[35466] = 29'b1_000101010001_010_0_001010100011;
      patterns[35467] = 29'b1_000101010001_011_0_010101000110;
      patterns[35468] = 29'b1_000101010001_100_1_100010101000;
      patterns[35469] = 29'b1_000101010001_101_0_110001010100;
      patterns[35470] = 29'b1_000101010001_110_1_000101010001;
      patterns[35471] = 29'b1_000101010001_111_1_000101010001;
      patterns[35472] = 29'b1_000101010010_000_1_000101010010;
      patterns[35473] = 29'b1_000101010010_001_1_010010000101;
      patterns[35474] = 29'b1_000101010010_010_0_001010100101;
      patterns[35475] = 29'b1_000101010010_011_0_010101001010;
      patterns[35476] = 29'b1_000101010010_100_0_100010101001;
      patterns[35477] = 29'b1_000101010010_101_1_010001010100;
      patterns[35478] = 29'b1_000101010010_110_1_000101010010;
      patterns[35479] = 29'b1_000101010010_111_1_000101010010;
      patterns[35480] = 29'b1_000101010011_000_1_000101010011;
      patterns[35481] = 29'b1_000101010011_001_1_010011000101;
      patterns[35482] = 29'b1_000101010011_010_0_001010100111;
      patterns[35483] = 29'b1_000101010011_011_0_010101001110;
      patterns[35484] = 29'b1_000101010011_100_1_100010101001;
      patterns[35485] = 29'b1_000101010011_101_1_110001010100;
      patterns[35486] = 29'b1_000101010011_110_1_000101010011;
      patterns[35487] = 29'b1_000101010011_111_1_000101010011;
      patterns[35488] = 29'b1_000101010100_000_1_000101010100;
      patterns[35489] = 29'b1_000101010100_001_1_010100000101;
      patterns[35490] = 29'b1_000101010100_010_0_001010101001;
      patterns[35491] = 29'b1_000101010100_011_0_010101010010;
      patterns[35492] = 29'b1_000101010100_100_0_100010101010;
      patterns[35493] = 29'b1_000101010100_101_0_010001010101;
      patterns[35494] = 29'b1_000101010100_110_1_000101010100;
      patterns[35495] = 29'b1_000101010100_111_1_000101010100;
      patterns[35496] = 29'b1_000101010101_000_1_000101010101;
      patterns[35497] = 29'b1_000101010101_001_1_010101000101;
      patterns[35498] = 29'b1_000101010101_010_0_001010101011;
      patterns[35499] = 29'b1_000101010101_011_0_010101010110;
      patterns[35500] = 29'b1_000101010101_100_1_100010101010;
      patterns[35501] = 29'b1_000101010101_101_0_110001010101;
      patterns[35502] = 29'b1_000101010101_110_1_000101010101;
      patterns[35503] = 29'b1_000101010101_111_1_000101010101;
      patterns[35504] = 29'b1_000101010110_000_1_000101010110;
      patterns[35505] = 29'b1_000101010110_001_1_010110000101;
      patterns[35506] = 29'b1_000101010110_010_0_001010101101;
      patterns[35507] = 29'b1_000101010110_011_0_010101011010;
      patterns[35508] = 29'b1_000101010110_100_0_100010101011;
      patterns[35509] = 29'b1_000101010110_101_1_010001010101;
      patterns[35510] = 29'b1_000101010110_110_1_000101010110;
      patterns[35511] = 29'b1_000101010110_111_1_000101010110;
      patterns[35512] = 29'b1_000101010111_000_1_000101010111;
      patterns[35513] = 29'b1_000101010111_001_1_010111000101;
      patterns[35514] = 29'b1_000101010111_010_0_001010101111;
      patterns[35515] = 29'b1_000101010111_011_0_010101011110;
      patterns[35516] = 29'b1_000101010111_100_1_100010101011;
      patterns[35517] = 29'b1_000101010111_101_1_110001010101;
      patterns[35518] = 29'b1_000101010111_110_1_000101010111;
      patterns[35519] = 29'b1_000101010111_111_1_000101010111;
      patterns[35520] = 29'b1_000101011000_000_1_000101011000;
      patterns[35521] = 29'b1_000101011000_001_1_011000000101;
      patterns[35522] = 29'b1_000101011000_010_0_001010110001;
      patterns[35523] = 29'b1_000101011000_011_0_010101100010;
      patterns[35524] = 29'b1_000101011000_100_0_100010101100;
      patterns[35525] = 29'b1_000101011000_101_0_010001010110;
      patterns[35526] = 29'b1_000101011000_110_1_000101011000;
      patterns[35527] = 29'b1_000101011000_111_1_000101011000;
      patterns[35528] = 29'b1_000101011001_000_1_000101011001;
      patterns[35529] = 29'b1_000101011001_001_1_011001000101;
      patterns[35530] = 29'b1_000101011001_010_0_001010110011;
      patterns[35531] = 29'b1_000101011001_011_0_010101100110;
      patterns[35532] = 29'b1_000101011001_100_1_100010101100;
      patterns[35533] = 29'b1_000101011001_101_0_110001010110;
      patterns[35534] = 29'b1_000101011001_110_1_000101011001;
      patterns[35535] = 29'b1_000101011001_111_1_000101011001;
      patterns[35536] = 29'b1_000101011010_000_1_000101011010;
      patterns[35537] = 29'b1_000101011010_001_1_011010000101;
      patterns[35538] = 29'b1_000101011010_010_0_001010110101;
      patterns[35539] = 29'b1_000101011010_011_0_010101101010;
      patterns[35540] = 29'b1_000101011010_100_0_100010101101;
      patterns[35541] = 29'b1_000101011010_101_1_010001010110;
      patterns[35542] = 29'b1_000101011010_110_1_000101011010;
      patterns[35543] = 29'b1_000101011010_111_1_000101011010;
      patterns[35544] = 29'b1_000101011011_000_1_000101011011;
      patterns[35545] = 29'b1_000101011011_001_1_011011000101;
      patterns[35546] = 29'b1_000101011011_010_0_001010110111;
      patterns[35547] = 29'b1_000101011011_011_0_010101101110;
      patterns[35548] = 29'b1_000101011011_100_1_100010101101;
      patterns[35549] = 29'b1_000101011011_101_1_110001010110;
      patterns[35550] = 29'b1_000101011011_110_1_000101011011;
      patterns[35551] = 29'b1_000101011011_111_1_000101011011;
      patterns[35552] = 29'b1_000101011100_000_1_000101011100;
      patterns[35553] = 29'b1_000101011100_001_1_011100000101;
      patterns[35554] = 29'b1_000101011100_010_0_001010111001;
      patterns[35555] = 29'b1_000101011100_011_0_010101110010;
      patterns[35556] = 29'b1_000101011100_100_0_100010101110;
      patterns[35557] = 29'b1_000101011100_101_0_010001010111;
      patterns[35558] = 29'b1_000101011100_110_1_000101011100;
      patterns[35559] = 29'b1_000101011100_111_1_000101011100;
      patterns[35560] = 29'b1_000101011101_000_1_000101011101;
      patterns[35561] = 29'b1_000101011101_001_1_011101000101;
      patterns[35562] = 29'b1_000101011101_010_0_001010111011;
      patterns[35563] = 29'b1_000101011101_011_0_010101110110;
      patterns[35564] = 29'b1_000101011101_100_1_100010101110;
      patterns[35565] = 29'b1_000101011101_101_0_110001010111;
      patterns[35566] = 29'b1_000101011101_110_1_000101011101;
      patterns[35567] = 29'b1_000101011101_111_1_000101011101;
      patterns[35568] = 29'b1_000101011110_000_1_000101011110;
      patterns[35569] = 29'b1_000101011110_001_1_011110000101;
      patterns[35570] = 29'b1_000101011110_010_0_001010111101;
      patterns[35571] = 29'b1_000101011110_011_0_010101111010;
      patterns[35572] = 29'b1_000101011110_100_0_100010101111;
      patterns[35573] = 29'b1_000101011110_101_1_010001010111;
      patterns[35574] = 29'b1_000101011110_110_1_000101011110;
      patterns[35575] = 29'b1_000101011110_111_1_000101011110;
      patterns[35576] = 29'b1_000101011111_000_1_000101011111;
      patterns[35577] = 29'b1_000101011111_001_1_011111000101;
      patterns[35578] = 29'b1_000101011111_010_0_001010111111;
      patterns[35579] = 29'b1_000101011111_011_0_010101111110;
      patterns[35580] = 29'b1_000101011111_100_1_100010101111;
      patterns[35581] = 29'b1_000101011111_101_1_110001010111;
      patterns[35582] = 29'b1_000101011111_110_1_000101011111;
      patterns[35583] = 29'b1_000101011111_111_1_000101011111;
      patterns[35584] = 29'b1_000101100000_000_1_000101100000;
      patterns[35585] = 29'b1_000101100000_001_1_100000000101;
      patterns[35586] = 29'b1_000101100000_010_0_001011000001;
      patterns[35587] = 29'b1_000101100000_011_0_010110000010;
      patterns[35588] = 29'b1_000101100000_100_0_100010110000;
      patterns[35589] = 29'b1_000101100000_101_0_010001011000;
      patterns[35590] = 29'b1_000101100000_110_1_000101100000;
      patterns[35591] = 29'b1_000101100000_111_1_000101100000;
      patterns[35592] = 29'b1_000101100001_000_1_000101100001;
      patterns[35593] = 29'b1_000101100001_001_1_100001000101;
      patterns[35594] = 29'b1_000101100001_010_0_001011000011;
      patterns[35595] = 29'b1_000101100001_011_0_010110000110;
      patterns[35596] = 29'b1_000101100001_100_1_100010110000;
      patterns[35597] = 29'b1_000101100001_101_0_110001011000;
      patterns[35598] = 29'b1_000101100001_110_1_000101100001;
      patterns[35599] = 29'b1_000101100001_111_1_000101100001;
      patterns[35600] = 29'b1_000101100010_000_1_000101100010;
      patterns[35601] = 29'b1_000101100010_001_1_100010000101;
      patterns[35602] = 29'b1_000101100010_010_0_001011000101;
      patterns[35603] = 29'b1_000101100010_011_0_010110001010;
      patterns[35604] = 29'b1_000101100010_100_0_100010110001;
      patterns[35605] = 29'b1_000101100010_101_1_010001011000;
      patterns[35606] = 29'b1_000101100010_110_1_000101100010;
      patterns[35607] = 29'b1_000101100010_111_1_000101100010;
      patterns[35608] = 29'b1_000101100011_000_1_000101100011;
      patterns[35609] = 29'b1_000101100011_001_1_100011000101;
      patterns[35610] = 29'b1_000101100011_010_0_001011000111;
      patterns[35611] = 29'b1_000101100011_011_0_010110001110;
      patterns[35612] = 29'b1_000101100011_100_1_100010110001;
      patterns[35613] = 29'b1_000101100011_101_1_110001011000;
      patterns[35614] = 29'b1_000101100011_110_1_000101100011;
      patterns[35615] = 29'b1_000101100011_111_1_000101100011;
      patterns[35616] = 29'b1_000101100100_000_1_000101100100;
      patterns[35617] = 29'b1_000101100100_001_1_100100000101;
      patterns[35618] = 29'b1_000101100100_010_0_001011001001;
      patterns[35619] = 29'b1_000101100100_011_0_010110010010;
      patterns[35620] = 29'b1_000101100100_100_0_100010110010;
      patterns[35621] = 29'b1_000101100100_101_0_010001011001;
      patterns[35622] = 29'b1_000101100100_110_1_000101100100;
      patterns[35623] = 29'b1_000101100100_111_1_000101100100;
      patterns[35624] = 29'b1_000101100101_000_1_000101100101;
      patterns[35625] = 29'b1_000101100101_001_1_100101000101;
      patterns[35626] = 29'b1_000101100101_010_0_001011001011;
      patterns[35627] = 29'b1_000101100101_011_0_010110010110;
      patterns[35628] = 29'b1_000101100101_100_1_100010110010;
      patterns[35629] = 29'b1_000101100101_101_0_110001011001;
      patterns[35630] = 29'b1_000101100101_110_1_000101100101;
      patterns[35631] = 29'b1_000101100101_111_1_000101100101;
      patterns[35632] = 29'b1_000101100110_000_1_000101100110;
      patterns[35633] = 29'b1_000101100110_001_1_100110000101;
      patterns[35634] = 29'b1_000101100110_010_0_001011001101;
      patterns[35635] = 29'b1_000101100110_011_0_010110011010;
      patterns[35636] = 29'b1_000101100110_100_0_100010110011;
      patterns[35637] = 29'b1_000101100110_101_1_010001011001;
      patterns[35638] = 29'b1_000101100110_110_1_000101100110;
      patterns[35639] = 29'b1_000101100110_111_1_000101100110;
      patterns[35640] = 29'b1_000101100111_000_1_000101100111;
      patterns[35641] = 29'b1_000101100111_001_1_100111000101;
      patterns[35642] = 29'b1_000101100111_010_0_001011001111;
      patterns[35643] = 29'b1_000101100111_011_0_010110011110;
      patterns[35644] = 29'b1_000101100111_100_1_100010110011;
      patterns[35645] = 29'b1_000101100111_101_1_110001011001;
      patterns[35646] = 29'b1_000101100111_110_1_000101100111;
      patterns[35647] = 29'b1_000101100111_111_1_000101100111;
      patterns[35648] = 29'b1_000101101000_000_1_000101101000;
      patterns[35649] = 29'b1_000101101000_001_1_101000000101;
      patterns[35650] = 29'b1_000101101000_010_0_001011010001;
      patterns[35651] = 29'b1_000101101000_011_0_010110100010;
      patterns[35652] = 29'b1_000101101000_100_0_100010110100;
      patterns[35653] = 29'b1_000101101000_101_0_010001011010;
      patterns[35654] = 29'b1_000101101000_110_1_000101101000;
      patterns[35655] = 29'b1_000101101000_111_1_000101101000;
      patterns[35656] = 29'b1_000101101001_000_1_000101101001;
      patterns[35657] = 29'b1_000101101001_001_1_101001000101;
      patterns[35658] = 29'b1_000101101001_010_0_001011010011;
      patterns[35659] = 29'b1_000101101001_011_0_010110100110;
      patterns[35660] = 29'b1_000101101001_100_1_100010110100;
      patterns[35661] = 29'b1_000101101001_101_0_110001011010;
      patterns[35662] = 29'b1_000101101001_110_1_000101101001;
      patterns[35663] = 29'b1_000101101001_111_1_000101101001;
      patterns[35664] = 29'b1_000101101010_000_1_000101101010;
      patterns[35665] = 29'b1_000101101010_001_1_101010000101;
      patterns[35666] = 29'b1_000101101010_010_0_001011010101;
      patterns[35667] = 29'b1_000101101010_011_0_010110101010;
      patterns[35668] = 29'b1_000101101010_100_0_100010110101;
      patterns[35669] = 29'b1_000101101010_101_1_010001011010;
      patterns[35670] = 29'b1_000101101010_110_1_000101101010;
      patterns[35671] = 29'b1_000101101010_111_1_000101101010;
      patterns[35672] = 29'b1_000101101011_000_1_000101101011;
      patterns[35673] = 29'b1_000101101011_001_1_101011000101;
      patterns[35674] = 29'b1_000101101011_010_0_001011010111;
      patterns[35675] = 29'b1_000101101011_011_0_010110101110;
      patterns[35676] = 29'b1_000101101011_100_1_100010110101;
      patterns[35677] = 29'b1_000101101011_101_1_110001011010;
      patterns[35678] = 29'b1_000101101011_110_1_000101101011;
      patterns[35679] = 29'b1_000101101011_111_1_000101101011;
      patterns[35680] = 29'b1_000101101100_000_1_000101101100;
      patterns[35681] = 29'b1_000101101100_001_1_101100000101;
      patterns[35682] = 29'b1_000101101100_010_0_001011011001;
      patterns[35683] = 29'b1_000101101100_011_0_010110110010;
      patterns[35684] = 29'b1_000101101100_100_0_100010110110;
      patterns[35685] = 29'b1_000101101100_101_0_010001011011;
      patterns[35686] = 29'b1_000101101100_110_1_000101101100;
      patterns[35687] = 29'b1_000101101100_111_1_000101101100;
      patterns[35688] = 29'b1_000101101101_000_1_000101101101;
      patterns[35689] = 29'b1_000101101101_001_1_101101000101;
      patterns[35690] = 29'b1_000101101101_010_0_001011011011;
      patterns[35691] = 29'b1_000101101101_011_0_010110110110;
      patterns[35692] = 29'b1_000101101101_100_1_100010110110;
      patterns[35693] = 29'b1_000101101101_101_0_110001011011;
      patterns[35694] = 29'b1_000101101101_110_1_000101101101;
      patterns[35695] = 29'b1_000101101101_111_1_000101101101;
      patterns[35696] = 29'b1_000101101110_000_1_000101101110;
      patterns[35697] = 29'b1_000101101110_001_1_101110000101;
      patterns[35698] = 29'b1_000101101110_010_0_001011011101;
      patterns[35699] = 29'b1_000101101110_011_0_010110111010;
      patterns[35700] = 29'b1_000101101110_100_0_100010110111;
      patterns[35701] = 29'b1_000101101110_101_1_010001011011;
      patterns[35702] = 29'b1_000101101110_110_1_000101101110;
      patterns[35703] = 29'b1_000101101110_111_1_000101101110;
      patterns[35704] = 29'b1_000101101111_000_1_000101101111;
      patterns[35705] = 29'b1_000101101111_001_1_101111000101;
      patterns[35706] = 29'b1_000101101111_010_0_001011011111;
      patterns[35707] = 29'b1_000101101111_011_0_010110111110;
      patterns[35708] = 29'b1_000101101111_100_1_100010110111;
      patterns[35709] = 29'b1_000101101111_101_1_110001011011;
      patterns[35710] = 29'b1_000101101111_110_1_000101101111;
      patterns[35711] = 29'b1_000101101111_111_1_000101101111;
      patterns[35712] = 29'b1_000101110000_000_1_000101110000;
      patterns[35713] = 29'b1_000101110000_001_1_110000000101;
      patterns[35714] = 29'b1_000101110000_010_0_001011100001;
      patterns[35715] = 29'b1_000101110000_011_0_010111000010;
      patterns[35716] = 29'b1_000101110000_100_0_100010111000;
      patterns[35717] = 29'b1_000101110000_101_0_010001011100;
      patterns[35718] = 29'b1_000101110000_110_1_000101110000;
      patterns[35719] = 29'b1_000101110000_111_1_000101110000;
      patterns[35720] = 29'b1_000101110001_000_1_000101110001;
      patterns[35721] = 29'b1_000101110001_001_1_110001000101;
      patterns[35722] = 29'b1_000101110001_010_0_001011100011;
      patterns[35723] = 29'b1_000101110001_011_0_010111000110;
      patterns[35724] = 29'b1_000101110001_100_1_100010111000;
      patterns[35725] = 29'b1_000101110001_101_0_110001011100;
      patterns[35726] = 29'b1_000101110001_110_1_000101110001;
      patterns[35727] = 29'b1_000101110001_111_1_000101110001;
      patterns[35728] = 29'b1_000101110010_000_1_000101110010;
      patterns[35729] = 29'b1_000101110010_001_1_110010000101;
      patterns[35730] = 29'b1_000101110010_010_0_001011100101;
      patterns[35731] = 29'b1_000101110010_011_0_010111001010;
      patterns[35732] = 29'b1_000101110010_100_0_100010111001;
      patterns[35733] = 29'b1_000101110010_101_1_010001011100;
      patterns[35734] = 29'b1_000101110010_110_1_000101110010;
      patterns[35735] = 29'b1_000101110010_111_1_000101110010;
      patterns[35736] = 29'b1_000101110011_000_1_000101110011;
      patterns[35737] = 29'b1_000101110011_001_1_110011000101;
      patterns[35738] = 29'b1_000101110011_010_0_001011100111;
      patterns[35739] = 29'b1_000101110011_011_0_010111001110;
      patterns[35740] = 29'b1_000101110011_100_1_100010111001;
      patterns[35741] = 29'b1_000101110011_101_1_110001011100;
      patterns[35742] = 29'b1_000101110011_110_1_000101110011;
      patterns[35743] = 29'b1_000101110011_111_1_000101110011;
      patterns[35744] = 29'b1_000101110100_000_1_000101110100;
      patterns[35745] = 29'b1_000101110100_001_1_110100000101;
      patterns[35746] = 29'b1_000101110100_010_0_001011101001;
      patterns[35747] = 29'b1_000101110100_011_0_010111010010;
      patterns[35748] = 29'b1_000101110100_100_0_100010111010;
      patterns[35749] = 29'b1_000101110100_101_0_010001011101;
      patterns[35750] = 29'b1_000101110100_110_1_000101110100;
      patterns[35751] = 29'b1_000101110100_111_1_000101110100;
      patterns[35752] = 29'b1_000101110101_000_1_000101110101;
      patterns[35753] = 29'b1_000101110101_001_1_110101000101;
      patterns[35754] = 29'b1_000101110101_010_0_001011101011;
      patterns[35755] = 29'b1_000101110101_011_0_010111010110;
      patterns[35756] = 29'b1_000101110101_100_1_100010111010;
      patterns[35757] = 29'b1_000101110101_101_0_110001011101;
      patterns[35758] = 29'b1_000101110101_110_1_000101110101;
      patterns[35759] = 29'b1_000101110101_111_1_000101110101;
      patterns[35760] = 29'b1_000101110110_000_1_000101110110;
      patterns[35761] = 29'b1_000101110110_001_1_110110000101;
      patterns[35762] = 29'b1_000101110110_010_0_001011101101;
      patterns[35763] = 29'b1_000101110110_011_0_010111011010;
      patterns[35764] = 29'b1_000101110110_100_0_100010111011;
      patterns[35765] = 29'b1_000101110110_101_1_010001011101;
      patterns[35766] = 29'b1_000101110110_110_1_000101110110;
      patterns[35767] = 29'b1_000101110110_111_1_000101110110;
      patterns[35768] = 29'b1_000101110111_000_1_000101110111;
      patterns[35769] = 29'b1_000101110111_001_1_110111000101;
      patterns[35770] = 29'b1_000101110111_010_0_001011101111;
      patterns[35771] = 29'b1_000101110111_011_0_010111011110;
      patterns[35772] = 29'b1_000101110111_100_1_100010111011;
      patterns[35773] = 29'b1_000101110111_101_1_110001011101;
      patterns[35774] = 29'b1_000101110111_110_1_000101110111;
      patterns[35775] = 29'b1_000101110111_111_1_000101110111;
      patterns[35776] = 29'b1_000101111000_000_1_000101111000;
      patterns[35777] = 29'b1_000101111000_001_1_111000000101;
      patterns[35778] = 29'b1_000101111000_010_0_001011110001;
      patterns[35779] = 29'b1_000101111000_011_0_010111100010;
      patterns[35780] = 29'b1_000101111000_100_0_100010111100;
      patterns[35781] = 29'b1_000101111000_101_0_010001011110;
      patterns[35782] = 29'b1_000101111000_110_1_000101111000;
      patterns[35783] = 29'b1_000101111000_111_1_000101111000;
      patterns[35784] = 29'b1_000101111001_000_1_000101111001;
      patterns[35785] = 29'b1_000101111001_001_1_111001000101;
      patterns[35786] = 29'b1_000101111001_010_0_001011110011;
      patterns[35787] = 29'b1_000101111001_011_0_010111100110;
      patterns[35788] = 29'b1_000101111001_100_1_100010111100;
      patterns[35789] = 29'b1_000101111001_101_0_110001011110;
      patterns[35790] = 29'b1_000101111001_110_1_000101111001;
      patterns[35791] = 29'b1_000101111001_111_1_000101111001;
      patterns[35792] = 29'b1_000101111010_000_1_000101111010;
      patterns[35793] = 29'b1_000101111010_001_1_111010000101;
      patterns[35794] = 29'b1_000101111010_010_0_001011110101;
      patterns[35795] = 29'b1_000101111010_011_0_010111101010;
      patterns[35796] = 29'b1_000101111010_100_0_100010111101;
      patterns[35797] = 29'b1_000101111010_101_1_010001011110;
      patterns[35798] = 29'b1_000101111010_110_1_000101111010;
      patterns[35799] = 29'b1_000101111010_111_1_000101111010;
      patterns[35800] = 29'b1_000101111011_000_1_000101111011;
      patterns[35801] = 29'b1_000101111011_001_1_111011000101;
      patterns[35802] = 29'b1_000101111011_010_0_001011110111;
      patterns[35803] = 29'b1_000101111011_011_0_010111101110;
      patterns[35804] = 29'b1_000101111011_100_1_100010111101;
      patterns[35805] = 29'b1_000101111011_101_1_110001011110;
      patterns[35806] = 29'b1_000101111011_110_1_000101111011;
      patterns[35807] = 29'b1_000101111011_111_1_000101111011;
      patterns[35808] = 29'b1_000101111100_000_1_000101111100;
      patterns[35809] = 29'b1_000101111100_001_1_111100000101;
      patterns[35810] = 29'b1_000101111100_010_0_001011111001;
      patterns[35811] = 29'b1_000101111100_011_0_010111110010;
      patterns[35812] = 29'b1_000101111100_100_0_100010111110;
      patterns[35813] = 29'b1_000101111100_101_0_010001011111;
      patterns[35814] = 29'b1_000101111100_110_1_000101111100;
      patterns[35815] = 29'b1_000101111100_111_1_000101111100;
      patterns[35816] = 29'b1_000101111101_000_1_000101111101;
      patterns[35817] = 29'b1_000101111101_001_1_111101000101;
      patterns[35818] = 29'b1_000101111101_010_0_001011111011;
      patterns[35819] = 29'b1_000101111101_011_0_010111110110;
      patterns[35820] = 29'b1_000101111101_100_1_100010111110;
      patterns[35821] = 29'b1_000101111101_101_0_110001011111;
      patterns[35822] = 29'b1_000101111101_110_1_000101111101;
      patterns[35823] = 29'b1_000101111101_111_1_000101111101;
      patterns[35824] = 29'b1_000101111110_000_1_000101111110;
      patterns[35825] = 29'b1_000101111110_001_1_111110000101;
      patterns[35826] = 29'b1_000101111110_010_0_001011111101;
      patterns[35827] = 29'b1_000101111110_011_0_010111111010;
      patterns[35828] = 29'b1_000101111110_100_0_100010111111;
      patterns[35829] = 29'b1_000101111110_101_1_010001011111;
      patterns[35830] = 29'b1_000101111110_110_1_000101111110;
      patterns[35831] = 29'b1_000101111110_111_1_000101111110;
      patterns[35832] = 29'b1_000101111111_000_1_000101111111;
      patterns[35833] = 29'b1_000101111111_001_1_111111000101;
      patterns[35834] = 29'b1_000101111111_010_0_001011111111;
      patterns[35835] = 29'b1_000101111111_011_0_010111111110;
      patterns[35836] = 29'b1_000101111111_100_1_100010111111;
      patterns[35837] = 29'b1_000101111111_101_1_110001011111;
      patterns[35838] = 29'b1_000101111111_110_1_000101111111;
      patterns[35839] = 29'b1_000101111111_111_1_000101111111;
      patterns[35840] = 29'b1_000110000000_000_1_000110000000;
      patterns[35841] = 29'b1_000110000000_001_1_000000000110;
      patterns[35842] = 29'b1_000110000000_010_0_001100000001;
      patterns[35843] = 29'b1_000110000000_011_0_011000000010;
      patterns[35844] = 29'b1_000110000000_100_0_100011000000;
      patterns[35845] = 29'b1_000110000000_101_0_010001100000;
      patterns[35846] = 29'b1_000110000000_110_1_000110000000;
      patterns[35847] = 29'b1_000110000000_111_1_000110000000;
      patterns[35848] = 29'b1_000110000001_000_1_000110000001;
      patterns[35849] = 29'b1_000110000001_001_1_000001000110;
      patterns[35850] = 29'b1_000110000001_010_0_001100000011;
      patterns[35851] = 29'b1_000110000001_011_0_011000000110;
      patterns[35852] = 29'b1_000110000001_100_1_100011000000;
      patterns[35853] = 29'b1_000110000001_101_0_110001100000;
      patterns[35854] = 29'b1_000110000001_110_1_000110000001;
      patterns[35855] = 29'b1_000110000001_111_1_000110000001;
      patterns[35856] = 29'b1_000110000010_000_1_000110000010;
      patterns[35857] = 29'b1_000110000010_001_1_000010000110;
      patterns[35858] = 29'b1_000110000010_010_0_001100000101;
      patterns[35859] = 29'b1_000110000010_011_0_011000001010;
      patterns[35860] = 29'b1_000110000010_100_0_100011000001;
      patterns[35861] = 29'b1_000110000010_101_1_010001100000;
      patterns[35862] = 29'b1_000110000010_110_1_000110000010;
      patterns[35863] = 29'b1_000110000010_111_1_000110000010;
      patterns[35864] = 29'b1_000110000011_000_1_000110000011;
      patterns[35865] = 29'b1_000110000011_001_1_000011000110;
      patterns[35866] = 29'b1_000110000011_010_0_001100000111;
      patterns[35867] = 29'b1_000110000011_011_0_011000001110;
      patterns[35868] = 29'b1_000110000011_100_1_100011000001;
      patterns[35869] = 29'b1_000110000011_101_1_110001100000;
      patterns[35870] = 29'b1_000110000011_110_1_000110000011;
      patterns[35871] = 29'b1_000110000011_111_1_000110000011;
      patterns[35872] = 29'b1_000110000100_000_1_000110000100;
      patterns[35873] = 29'b1_000110000100_001_1_000100000110;
      patterns[35874] = 29'b1_000110000100_010_0_001100001001;
      patterns[35875] = 29'b1_000110000100_011_0_011000010010;
      patterns[35876] = 29'b1_000110000100_100_0_100011000010;
      patterns[35877] = 29'b1_000110000100_101_0_010001100001;
      patterns[35878] = 29'b1_000110000100_110_1_000110000100;
      patterns[35879] = 29'b1_000110000100_111_1_000110000100;
      patterns[35880] = 29'b1_000110000101_000_1_000110000101;
      patterns[35881] = 29'b1_000110000101_001_1_000101000110;
      patterns[35882] = 29'b1_000110000101_010_0_001100001011;
      patterns[35883] = 29'b1_000110000101_011_0_011000010110;
      patterns[35884] = 29'b1_000110000101_100_1_100011000010;
      patterns[35885] = 29'b1_000110000101_101_0_110001100001;
      patterns[35886] = 29'b1_000110000101_110_1_000110000101;
      patterns[35887] = 29'b1_000110000101_111_1_000110000101;
      patterns[35888] = 29'b1_000110000110_000_1_000110000110;
      patterns[35889] = 29'b1_000110000110_001_1_000110000110;
      patterns[35890] = 29'b1_000110000110_010_0_001100001101;
      patterns[35891] = 29'b1_000110000110_011_0_011000011010;
      patterns[35892] = 29'b1_000110000110_100_0_100011000011;
      patterns[35893] = 29'b1_000110000110_101_1_010001100001;
      patterns[35894] = 29'b1_000110000110_110_1_000110000110;
      patterns[35895] = 29'b1_000110000110_111_1_000110000110;
      patterns[35896] = 29'b1_000110000111_000_1_000110000111;
      patterns[35897] = 29'b1_000110000111_001_1_000111000110;
      patterns[35898] = 29'b1_000110000111_010_0_001100001111;
      patterns[35899] = 29'b1_000110000111_011_0_011000011110;
      patterns[35900] = 29'b1_000110000111_100_1_100011000011;
      patterns[35901] = 29'b1_000110000111_101_1_110001100001;
      patterns[35902] = 29'b1_000110000111_110_1_000110000111;
      patterns[35903] = 29'b1_000110000111_111_1_000110000111;
      patterns[35904] = 29'b1_000110001000_000_1_000110001000;
      patterns[35905] = 29'b1_000110001000_001_1_001000000110;
      patterns[35906] = 29'b1_000110001000_010_0_001100010001;
      patterns[35907] = 29'b1_000110001000_011_0_011000100010;
      patterns[35908] = 29'b1_000110001000_100_0_100011000100;
      patterns[35909] = 29'b1_000110001000_101_0_010001100010;
      patterns[35910] = 29'b1_000110001000_110_1_000110001000;
      patterns[35911] = 29'b1_000110001000_111_1_000110001000;
      patterns[35912] = 29'b1_000110001001_000_1_000110001001;
      patterns[35913] = 29'b1_000110001001_001_1_001001000110;
      patterns[35914] = 29'b1_000110001001_010_0_001100010011;
      patterns[35915] = 29'b1_000110001001_011_0_011000100110;
      patterns[35916] = 29'b1_000110001001_100_1_100011000100;
      patterns[35917] = 29'b1_000110001001_101_0_110001100010;
      patterns[35918] = 29'b1_000110001001_110_1_000110001001;
      patterns[35919] = 29'b1_000110001001_111_1_000110001001;
      patterns[35920] = 29'b1_000110001010_000_1_000110001010;
      patterns[35921] = 29'b1_000110001010_001_1_001010000110;
      patterns[35922] = 29'b1_000110001010_010_0_001100010101;
      patterns[35923] = 29'b1_000110001010_011_0_011000101010;
      patterns[35924] = 29'b1_000110001010_100_0_100011000101;
      patterns[35925] = 29'b1_000110001010_101_1_010001100010;
      patterns[35926] = 29'b1_000110001010_110_1_000110001010;
      patterns[35927] = 29'b1_000110001010_111_1_000110001010;
      patterns[35928] = 29'b1_000110001011_000_1_000110001011;
      patterns[35929] = 29'b1_000110001011_001_1_001011000110;
      patterns[35930] = 29'b1_000110001011_010_0_001100010111;
      patterns[35931] = 29'b1_000110001011_011_0_011000101110;
      patterns[35932] = 29'b1_000110001011_100_1_100011000101;
      patterns[35933] = 29'b1_000110001011_101_1_110001100010;
      patterns[35934] = 29'b1_000110001011_110_1_000110001011;
      patterns[35935] = 29'b1_000110001011_111_1_000110001011;
      patterns[35936] = 29'b1_000110001100_000_1_000110001100;
      patterns[35937] = 29'b1_000110001100_001_1_001100000110;
      patterns[35938] = 29'b1_000110001100_010_0_001100011001;
      patterns[35939] = 29'b1_000110001100_011_0_011000110010;
      patterns[35940] = 29'b1_000110001100_100_0_100011000110;
      patterns[35941] = 29'b1_000110001100_101_0_010001100011;
      patterns[35942] = 29'b1_000110001100_110_1_000110001100;
      patterns[35943] = 29'b1_000110001100_111_1_000110001100;
      patterns[35944] = 29'b1_000110001101_000_1_000110001101;
      patterns[35945] = 29'b1_000110001101_001_1_001101000110;
      patterns[35946] = 29'b1_000110001101_010_0_001100011011;
      patterns[35947] = 29'b1_000110001101_011_0_011000110110;
      patterns[35948] = 29'b1_000110001101_100_1_100011000110;
      patterns[35949] = 29'b1_000110001101_101_0_110001100011;
      patterns[35950] = 29'b1_000110001101_110_1_000110001101;
      patterns[35951] = 29'b1_000110001101_111_1_000110001101;
      patterns[35952] = 29'b1_000110001110_000_1_000110001110;
      patterns[35953] = 29'b1_000110001110_001_1_001110000110;
      patterns[35954] = 29'b1_000110001110_010_0_001100011101;
      patterns[35955] = 29'b1_000110001110_011_0_011000111010;
      patterns[35956] = 29'b1_000110001110_100_0_100011000111;
      patterns[35957] = 29'b1_000110001110_101_1_010001100011;
      patterns[35958] = 29'b1_000110001110_110_1_000110001110;
      patterns[35959] = 29'b1_000110001110_111_1_000110001110;
      patterns[35960] = 29'b1_000110001111_000_1_000110001111;
      patterns[35961] = 29'b1_000110001111_001_1_001111000110;
      patterns[35962] = 29'b1_000110001111_010_0_001100011111;
      patterns[35963] = 29'b1_000110001111_011_0_011000111110;
      patterns[35964] = 29'b1_000110001111_100_1_100011000111;
      patterns[35965] = 29'b1_000110001111_101_1_110001100011;
      patterns[35966] = 29'b1_000110001111_110_1_000110001111;
      patterns[35967] = 29'b1_000110001111_111_1_000110001111;
      patterns[35968] = 29'b1_000110010000_000_1_000110010000;
      patterns[35969] = 29'b1_000110010000_001_1_010000000110;
      patterns[35970] = 29'b1_000110010000_010_0_001100100001;
      patterns[35971] = 29'b1_000110010000_011_0_011001000010;
      patterns[35972] = 29'b1_000110010000_100_0_100011001000;
      patterns[35973] = 29'b1_000110010000_101_0_010001100100;
      patterns[35974] = 29'b1_000110010000_110_1_000110010000;
      patterns[35975] = 29'b1_000110010000_111_1_000110010000;
      patterns[35976] = 29'b1_000110010001_000_1_000110010001;
      patterns[35977] = 29'b1_000110010001_001_1_010001000110;
      patterns[35978] = 29'b1_000110010001_010_0_001100100011;
      patterns[35979] = 29'b1_000110010001_011_0_011001000110;
      patterns[35980] = 29'b1_000110010001_100_1_100011001000;
      patterns[35981] = 29'b1_000110010001_101_0_110001100100;
      patterns[35982] = 29'b1_000110010001_110_1_000110010001;
      patterns[35983] = 29'b1_000110010001_111_1_000110010001;
      patterns[35984] = 29'b1_000110010010_000_1_000110010010;
      patterns[35985] = 29'b1_000110010010_001_1_010010000110;
      patterns[35986] = 29'b1_000110010010_010_0_001100100101;
      patterns[35987] = 29'b1_000110010010_011_0_011001001010;
      patterns[35988] = 29'b1_000110010010_100_0_100011001001;
      patterns[35989] = 29'b1_000110010010_101_1_010001100100;
      patterns[35990] = 29'b1_000110010010_110_1_000110010010;
      patterns[35991] = 29'b1_000110010010_111_1_000110010010;
      patterns[35992] = 29'b1_000110010011_000_1_000110010011;
      patterns[35993] = 29'b1_000110010011_001_1_010011000110;
      patterns[35994] = 29'b1_000110010011_010_0_001100100111;
      patterns[35995] = 29'b1_000110010011_011_0_011001001110;
      patterns[35996] = 29'b1_000110010011_100_1_100011001001;
      patterns[35997] = 29'b1_000110010011_101_1_110001100100;
      patterns[35998] = 29'b1_000110010011_110_1_000110010011;
      patterns[35999] = 29'b1_000110010011_111_1_000110010011;
      patterns[36000] = 29'b1_000110010100_000_1_000110010100;
      patterns[36001] = 29'b1_000110010100_001_1_010100000110;
      patterns[36002] = 29'b1_000110010100_010_0_001100101001;
      patterns[36003] = 29'b1_000110010100_011_0_011001010010;
      patterns[36004] = 29'b1_000110010100_100_0_100011001010;
      patterns[36005] = 29'b1_000110010100_101_0_010001100101;
      patterns[36006] = 29'b1_000110010100_110_1_000110010100;
      patterns[36007] = 29'b1_000110010100_111_1_000110010100;
      patterns[36008] = 29'b1_000110010101_000_1_000110010101;
      patterns[36009] = 29'b1_000110010101_001_1_010101000110;
      patterns[36010] = 29'b1_000110010101_010_0_001100101011;
      patterns[36011] = 29'b1_000110010101_011_0_011001010110;
      patterns[36012] = 29'b1_000110010101_100_1_100011001010;
      patterns[36013] = 29'b1_000110010101_101_0_110001100101;
      patterns[36014] = 29'b1_000110010101_110_1_000110010101;
      patterns[36015] = 29'b1_000110010101_111_1_000110010101;
      patterns[36016] = 29'b1_000110010110_000_1_000110010110;
      patterns[36017] = 29'b1_000110010110_001_1_010110000110;
      patterns[36018] = 29'b1_000110010110_010_0_001100101101;
      patterns[36019] = 29'b1_000110010110_011_0_011001011010;
      patterns[36020] = 29'b1_000110010110_100_0_100011001011;
      patterns[36021] = 29'b1_000110010110_101_1_010001100101;
      patterns[36022] = 29'b1_000110010110_110_1_000110010110;
      patterns[36023] = 29'b1_000110010110_111_1_000110010110;
      patterns[36024] = 29'b1_000110010111_000_1_000110010111;
      patterns[36025] = 29'b1_000110010111_001_1_010111000110;
      patterns[36026] = 29'b1_000110010111_010_0_001100101111;
      patterns[36027] = 29'b1_000110010111_011_0_011001011110;
      patterns[36028] = 29'b1_000110010111_100_1_100011001011;
      patterns[36029] = 29'b1_000110010111_101_1_110001100101;
      patterns[36030] = 29'b1_000110010111_110_1_000110010111;
      patterns[36031] = 29'b1_000110010111_111_1_000110010111;
      patterns[36032] = 29'b1_000110011000_000_1_000110011000;
      patterns[36033] = 29'b1_000110011000_001_1_011000000110;
      patterns[36034] = 29'b1_000110011000_010_0_001100110001;
      patterns[36035] = 29'b1_000110011000_011_0_011001100010;
      patterns[36036] = 29'b1_000110011000_100_0_100011001100;
      patterns[36037] = 29'b1_000110011000_101_0_010001100110;
      patterns[36038] = 29'b1_000110011000_110_1_000110011000;
      patterns[36039] = 29'b1_000110011000_111_1_000110011000;
      patterns[36040] = 29'b1_000110011001_000_1_000110011001;
      patterns[36041] = 29'b1_000110011001_001_1_011001000110;
      patterns[36042] = 29'b1_000110011001_010_0_001100110011;
      patterns[36043] = 29'b1_000110011001_011_0_011001100110;
      patterns[36044] = 29'b1_000110011001_100_1_100011001100;
      patterns[36045] = 29'b1_000110011001_101_0_110001100110;
      patterns[36046] = 29'b1_000110011001_110_1_000110011001;
      patterns[36047] = 29'b1_000110011001_111_1_000110011001;
      patterns[36048] = 29'b1_000110011010_000_1_000110011010;
      patterns[36049] = 29'b1_000110011010_001_1_011010000110;
      patterns[36050] = 29'b1_000110011010_010_0_001100110101;
      patterns[36051] = 29'b1_000110011010_011_0_011001101010;
      patterns[36052] = 29'b1_000110011010_100_0_100011001101;
      patterns[36053] = 29'b1_000110011010_101_1_010001100110;
      patterns[36054] = 29'b1_000110011010_110_1_000110011010;
      patterns[36055] = 29'b1_000110011010_111_1_000110011010;
      patterns[36056] = 29'b1_000110011011_000_1_000110011011;
      patterns[36057] = 29'b1_000110011011_001_1_011011000110;
      patterns[36058] = 29'b1_000110011011_010_0_001100110111;
      patterns[36059] = 29'b1_000110011011_011_0_011001101110;
      patterns[36060] = 29'b1_000110011011_100_1_100011001101;
      patterns[36061] = 29'b1_000110011011_101_1_110001100110;
      patterns[36062] = 29'b1_000110011011_110_1_000110011011;
      patterns[36063] = 29'b1_000110011011_111_1_000110011011;
      patterns[36064] = 29'b1_000110011100_000_1_000110011100;
      patterns[36065] = 29'b1_000110011100_001_1_011100000110;
      patterns[36066] = 29'b1_000110011100_010_0_001100111001;
      patterns[36067] = 29'b1_000110011100_011_0_011001110010;
      patterns[36068] = 29'b1_000110011100_100_0_100011001110;
      patterns[36069] = 29'b1_000110011100_101_0_010001100111;
      patterns[36070] = 29'b1_000110011100_110_1_000110011100;
      patterns[36071] = 29'b1_000110011100_111_1_000110011100;
      patterns[36072] = 29'b1_000110011101_000_1_000110011101;
      patterns[36073] = 29'b1_000110011101_001_1_011101000110;
      patterns[36074] = 29'b1_000110011101_010_0_001100111011;
      patterns[36075] = 29'b1_000110011101_011_0_011001110110;
      patterns[36076] = 29'b1_000110011101_100_1_100011001110;
      patterns[36077] = 29'b1_000110011101_101_0_110001100111;
      patterns[36078] = 29'b1_000110011101_110_1_000110011101;
      patterns[36079] = 29'b1_000110011101_111_1_000110011101;
      patterns[36080] = 29'b1_000110011110_000_1_000110011110;
      patterns[36081] = 29'b1_000110011110_001_1_011110000110;
      patterns[36082] = 29'b1_000110011110_010_0_001100111101;
      patterns[36083] = 29'b1_000110011110_011_0_011001111010;
      patterns[36084] = 29'b1_000110011110_100_0_100011001111;
      patterns[36085] = 29'b1_000110011110_101_1_010001100111;
      patterns[36086] = 29'b1_000110011110_110_1_000110011110;
      patterns[36087] = 29'b1_000110011110_111_1_000110011110;
      patterns[36088] = 29'b1_000110011111_000_1_000110011111;
      patterns[36089] = 29'b1_000110011111_001_1_011111000110;
      patterns[36090] = 29'b1_000110011111_010_0_001100111111;
      patterns[36091] = 29'b1_000110011111_011_0_011001111110;
      patterns[36092] = 29'b1_000110011111_100_1_100011001111;
      patterns[36093] = 29'b1_000110011111_101_1_110001100111;
      patterns[36094] = 29'b1_000110011111_110_1_000110011111;
      patterns[36095] = 29'b1_000110011111_111_1_000110011111;
      patterns[36096] = 29'b1_000110100000_000_1_000110100000;
      patterns[36097] = 29'b1_000110100000_001_1_100000000110;
      patterns[36098] = 29'b1_000110100000_010_0_001101000001;
      patterns[36099] = 29'b1_000110100000_011_0_011010000010;
      patterns[36100] = 29'b1_000110100000_100_0_100011010000;
      patterns[36101] = 29'b1_000110100000_101_0_010001101000;
      patterns[36102] = 29'b1_000110100000_110_1_000110100000;
      patterns[36103] = 29'b1_000110100000_111_1_000110100000;
      patterns[36104] = 29'b1_000110100001_000_1_000110100001;
      patterns[36105] = 29'b1_000110100001_001_1_100001000110;
      patterns[36106] = 29'b1_000110100001_010_0_001101000011;
      patterns[36107] = 29'b1_000110100001_011_0_011010000110;
      patterns[36108] = 29'b1_000110100001_100_1_100011010000;
      patterns[36109] = 29'b1_000110100001_101_0_110001101000;
      patterns[36110] = 29'b1_000110100001_110_1_000110100001;
      patterns[36111] = 29'b1_000110100001_111_1_000110100001;
      patterns[36112] = 29'b1_000110100010_000_1_000110100010;
      patterns[36113] = 29'b1_000110100010_001_1_100010000110;
      patterns[36114] = 29'b1_000110100010_010_0_001101000101;
      patterns[36115] = 29'b1_000110100010_011_0_011010001010;
      patterns[36116] = 29'b1_000110100010_100_0_100011010001;
      patterns[36117] = 29'b1_000110100010_101_1_010001101000;
      patterns[36118] = 29'b1_000110100010_110_1_000110100010;
      patterns[36119] = 29'b1_000110100010_111_1_000110100010;
      patterns[36120] = 29'b1_000110100011_000_1_000110100011;
      patterns[36121] = 29'b1_000110100011_001_1_100011000110;
      patterns[36122] = 29'b1_000110100011_010_0_001101000111;
      patterns[36123] = 29'b1_000110100011_011_0_011010001110;
      patterns[36124] = 29'b1_000110100011_100_1_100011010001;
      patterns[36125] = 29'b1_000110100011_101_1_110001101000;
      patterns[36126] = 29'b1_000110100011_110_1_000110100011;
      patterns[36127] = 29'b1_000110100011_111_1_000110100011;
      patterns[36128] = 29'b1_000110100100_000_1_000110100100;
      patterns[36129] = 29'b1_000110100100_001_1_100100000110;
      patterns[36130] = 29'b1_000110100100_010_0_001101001001;
      patterns[36131] = 29'b1_000110100100_011_0_011010010010;
      patterns[36132] = 29'b1_000110100100_100_0_100011010010;
      patterns[36133] = 29'b1_000110100100_101_0_010001101001;
      patterns[36134] = 29'b1_000110100100_110_1_000110100100;
      patterns[36135] = 29'b1_000110100100_111_1_000110100100;
      patterns[36136] = 29'b1_000110100101_000_1_000110100101;
      patterns[36137] = 29'b1_000110100101_001_1_100101000110;
      patterns[36138] = 29'b1_000110100101_010_0_001101001011;
      patterns[36139] = 29'b1_000110100101_011_0_011010010110;
      patterns[36140] = 29'b1_000110100101_100_1_100011010010;
      patterns[36141] = 29'b1_000110100101_101_0_110001101001;
      patterns[36142] = 29'b1_000110100101_110_1_000110100101;
      patterns[36143] = 29'b1_000110100101_111_1_000110100101;
      patterns[36144] = 29'b1_000110100110_000_1_000110100110;
      patterns[36145] = 29'b1_000110100110_001_1_100110000110;
      patterns[36146] = 29'b1_000110100110_010_0_001101001101;
      patterns[36147] = 29'b1_000110100110_011_0_011010011010;
      patterns[36148] = 29'b1_000110100110_100_0_100011010011;
      patterns[36149] = 29'b1_000110100110_101_1_010001101001;
      patterns[36150] = 29'b1_000110100110_110_1_000110100110;
      patterns[36151] = 29'b1_000110100110_111_1_000110100110;
      patterns[36152] = 29'b1_000110100111_000_1_000110100111;
      patterns[36153] = 29'b1_000110100111_001_1_100111000110;
      patterns[36154] = 29'b1_000110100111_010_0_001101001111;
      patterns[36155] = 29'b1_000110100111_011_0_011010011110;
      patterns[36156] = 29'b1_000110100111_100_1_100011010011;
      patterns[36157] = 29'b1_000110100111_101_1_110001101001;
      patterns[36158] = 29'b1_000110100111_110_1_000110100111;
      patterns[36159] = 29'b1_000110100111_111_1_000110100111;
      patterns[36160] = 29'b1_000110101000_000_1_000110101000;
      patterns[36161] = 29'b1_000110101000_001_1_101000000110;
      patterns[36162] = 29'b1_000110101000_010_0_001101010001;
      patterns[36163] = 29'b1_000110101000_011_0_011010100010;
      patterns[36164] = 29'b1_000110101000_100_0_100011010100;
      patterns[36165] = 29'b1_000110101000_101_0_010001101010;
      patterns[36166] = 29'b1_000110101000_110_1_000110101000;
      patterns[36167] = 29'b1_000110101000_111_1_000110101000;
      patterns[36168] = 29'b1_000110101001_000_1_000110101001;
      patterns[36169] = 29'b1_000110101001_001_1_101001000110;
      patterns[36170] = 29'b1_000110101001_010_0_001101010011;
      patterns[36171] = 29'b1_000110101001_011_0_011010100110;
      patterns[36172] = 29'b1_000110101001_100_1_100011010100;
      patterns[36173] = 29'b1_000110101001_101_0_110001101010;
      patterns[36174] = 29'b1_000110101001_110_1_000110101001;
      patterns[36175] = 29'b1_000110101001_111_1_000110101001;
      patterns[36176] = 29'b1_000110101010_000_1_000110101010;
      patterns[36177] = 29'b1_000110101010_001_1_101010000110;
      patterns[36178] = 29'b1_000110101010_010_0_001101010101;
      patterns[36179] = 29'b1_000110101010_011_0_011010101010;
      patterns[36180] = 29'b1_000110101010_100_0_100011010101;
      patterns[36181] = 29'b1_000110101010_101_1_010001101010;
      patterns[36182] = 29'b1_000110101010_110_1_000110101010;
      patterns[36183] = 29'b1_000110101010_111_1_000110101010;
      patterns[36184] = 29'b1_000110101011_000_1_000110101011;
      patterns[36185] = 29'b1_000110101011_001_1_101011000110;
      patterns[36186] = 29'b1_000110101011_010_0_001101010111;
      patterns[36187] = 29'b1_000110101011_011_0_011010101110;
      patterns[36188] = 29'b1_000110101011_100_1_100011010101;
      patterns[36189] = 29'b1_000110101011_101_1_110001101010;
      patterns[36190] = 29'b1_000110101011_110_1_000110101011;
      patterns[36191] = 29'b1_000110101011_111_1_000110101011;
      patterns[36192] = 29'b1_000110101100_000_1_000110101100;
      patterns[36193] = 29'b1_000110101100_001_1_101100000110;
      patterns[36194] = 29'b1_000110101100_010_0_001101011001;
      patterns[36195] = 29'b1_000110101100_011_0_011010110010;
      patterns[36196] = 29'b1_000110101100_100_0_100011010110;
      patterns[36197] = 29'b1_000110101100_101_0_010001101011;
      patterns[36198] = 29'b1_000110101100_110_1_000110101100;
      patterns[36199] = 29'b1_000110101100_111_1_000110101100;
      patterns[36200] = 29'b1_000110101101_000_1_000110101101;
      patterns[36201] = 29'b1_000110101101_001_1_101101000110;
      patterns[36202] = 29'b1_000110101101_010_0_001101011011;
      patterns[36203] = 29'b1_000110101101_011_0_011010110110;
      patterns[36204] = 29'b1_000110101101_100_1_100011010110;
      patterns[36205] = 29'b1_000110101101_101_0_110001101011;
      patterns[36206] = 29'b1_000110101101_110_1_000110101101;
      patterns[36207] = 29'b1_000110101101_111_1_000110101101;
      patterns[36208] = 29'b1_000110101110_000_1_000110101110;
      patterns[36209] = 29'b1_000110101110_001_1_101110000110;
      patterns[36210] = 29'b1_000110101110_010_0_001101011101;
      patterns[36211] = 29'b1_000110101110_011_0_011010111010;
      patterns[36212] = 29'b1_000110101110_100_0_100011010111;
      patterns[36213] = 29'b1_000110101110_101_1_010001101011;
      patterns[36214] = 29'b1_000110101110_110_1_000110101110;
      patterns[36215] = 29'b1_000110101110_111_1_000110101110;
      patterns[36216] = 29'b1_000110101111_000_1_000110101111;
      patterns[36217] = 29'b1_000110101111_001_1_101111000110;
      patterns[36218] = 29'b1_000110101111_010_0_001101011111;
      patterns[36219] = 29'b1_000110101111_011_0_011010111110;
      patterns[36220] = 29'b1_000110101111_100_1_100011010111;
      patterns[36221] = 29'b1_000110101111_101_1_110001101011;
      patterns[36222] = 29'b1_000110101111_110_1_000110101111;
      patterns[36223] = 29'b1_000110101111_111_1_000110101111;
      patterns[36224] = 29'b1_000110110000_000_1_000110110000;
      patterns[36225] = 29'b1_000110110000_001_1_110000000110;
      patterns[36226] = 29'b1_000110110000_010_0_001101100001;
      patterns[36227] = 29'b1_000110110000_011_0_011011000010;
      patterns[36228] = 29'b1_000110110000_100_0_100011011000;
      patterns[36229] = 29'b1_000110110000_101_0_010001101100;
      patterns[36230] = 29'b1_000110110000_110_1_000110110000;
      patterns[36231] = 29'b1_000110110000_111_1_000110110000;
      patterns[36232] = 29'b1_000110110001_000_1_000110110001;
      patterns[36233] = 29'b1_000110110001_001_1_110001000110;
      patterns[36234] = 29'b1_000110110001_010_0_001101100011;
      patterns[36235] = 29'b1_000110110001_011_0_011011000110;
      patterns[36236] = 29'b1_000110110001_100_1_100011011000;
      patterns[36237] = 29'b1_000110110001_101_0_110001101100;
      patterns[36238] = 29'b1_000110110001_110_1_000110110001;
      patterns[36239] = 29'b1_000110110001_111_1_000110110001;
      patterns[36240] = 29'b1_000110110010_000_1_000110110010;
      patterns[36241] = 29'b1_000110110010_001_1_110010000110;
      patterns[36242] = 29'b1_000110110010_010_0_001101100101;
      patterns[36243] = 29'b1_000110110010_011_0_011011001010;
      patterns[36244] = 29'b1_000110110010_100_0_100011011001;
      patterns[36245] = 29'b1_000110110010_101_1_010001101100;
      patterns[36246] = 29'b1_000110110010_110_1_000110110010;
      patterns[36247] = 29'b1_000110110010_111_1_000110110010;
      patterns[36248] = 29'b1_000110110011_000_1_000110110011;
      patterns[36249] = 29'b1_000110110011_001_1_110011000110;
      patterns[36250] = 29'b1_000110110011_010_0_001101100111;
      patterns[36251] = 29'b1_000110110011_011_0_011011001110;
      patterns[36252] = 29'b1_000110110011_100_1_100011011001;
      patterns[36253] = 29'b1_000110110011_101_1_110001101100;
      patterns[36254] = 29'b1_000110110011_110_1_000110110011;
      patterns[36255] = 29'b1_000110110011_111_1_000110110011;
      patterns[36256] = 29'b1_000110110100_000_1_000110110100;
      patterns[36257] = 29'b1_000110110100_001_1_110100000110;
      patterns[36258] = 29'b1_000110110100_010_0_001101101001;
      patterns[36259] = 29'b1_000110110100_011_0_011011010010;
      patterns[36260] = 29'b1_000110110100_100_0_100011011010;
      patterns[36261] = 29'b1_000110110100_101_0_010001101101;
      patterns[36262] = 29'b1_000110110100_110_1_000110110100;
      patterns[36263] = 29'b1_000110110100_111_1_000110110100;
      patterns[36264] = 29'b1_000110110101_000_1_000110110101;
      patterns[36265] = 29'b1_000110110101_001_1_110101000110;
      patterns[36266] = 29'b1_000110110101_010_0_001101101011;
      patterns[36267] = 29'b1_000110110101_011_0_011011010110;
      patterns[36268] = 29'b1_000110110101_100_1_100011011010;
      patterns[36269] = 29'b1_000110110101_101_0_110001101101;
      patterns[36270] = 29'b1_000110110101_110_1_000110110101;
      patterns[36271] = 29'b1_000110110101_111_1_000110110101;
      patterns[36272] = 29'b1_000110110110_000_1_000110110110;
      patterns[36273] = 29'b1_000110110110_001_1_110110000110;
      patterns[36274] = 29'b1_000110110110_010_0_001101101101;
      patterns[36275] = 29'b1_000110110110_011_0_011011011010;
      patterns[36276] = 29'b1_000110110110_100_0_100011011011;
      patterns[36277] = 29'b1_000110110110_101_1_010001101101;
      patterns[36278] = 29'b1_000110110110_110_1_000110110110;
      patterns[36279] = 29'b1_000110110110_111_1_000110110110;
      patterns[36280] = 29'b1_000110110111_000_1_000110110111;
      patterns[36281] = 29'b1_000110110111_001_1_110111000110;
      patterns[36282] = 29'b1_000110110111_010_0_001101101111;
      patterns[36283] = 29'b1_000110110111_011_0_011011011110;
      patterns[36284] = 29'b1_000110110111_100_1_100011011011;
      patterns[36285] = 29'b1_000110110111_101_1_110001101101;
      patterns[36286] = 29'b1_000110110111_110_1_000110110111;
      patterns[36287] = 29'b1_000110110111_111_1_000110110111;
      patterns[36288] = 29'b1_000110111000_000_1_000110111000;
      patterns[36289] = 29'b1_000110111000_001_1_111000000110;
      patterns[36290] = 29'b1_000110111000_010_0_001101110001;
      patterns[36291] = 29'b1_000110111000_011_0_011011100010;
      patterns[36292] = 29'b1_000110111000_100_0_100011011100;
      patterns[36293] = 29'b1_000110111000_101_0_010001101110;
      patterns[36294] = 29'b1_000110111000_110_1_000110111000;
      patterns[36295] = 29'b1_000110111000_111_1_000110111000;
      patterns[36296] = 29'b1_000110111001_000_1_000110111001;
      patterns[36297] = 29'b1_000110111001_001_1_111001000110;
      patterns[36298] = 29'b1_000110111001_010_0_001101110011;
      patterns[36299] = 29'b1_000110111001_011_0_011011100110;
      patterns[36300] = 29'b1_000110111001_100_1_100011011100;
      patterns[36301] = 29'b1_000110111001_101_0_110001101110;
      patterns[36302] = 29'b1_000110111001_110_1_000110111001;
      patterns[36303] = 29'b1_000110111001_111_1_000110111001;
      patterns[36304] = 29'b1_000110111010_000_1_000110111010;
      patterns[36305] = 29'b1_000110111010_001_1_111010000110;
      patterns[36306] = 29'b1_000110111010_010_0_001101110101;
      patterns[36307] = 29'b1_000110111010_011_0_011011101010;
      patterns[36308] = 29'b1_000110111010_100_0_100011011101;
      patterns[36309] = 29'b1_000110111010_101_1_010001101110;
      patterns[36310] = 29'b1_000110111010_110_1_000110111010;
      patterns[36311] = 29'b1_000110111010_111_1_000110111010;
      patterns[36312] = 29'b1_000110111011_000_1_000110111011;
      patterns[36313] = 29'b1_000110111011_001_1_111011000110;
      patterns[36314] = 29'b1_000110111011_010_0_001101110111;
      patterns[36315] = 29'b1_000110111011_011_0_011011101110;
      patterns[36316] = 29'b1_000110111011_100_1_100011011101;
      patterns[36317] = 29'b1_000110111011_101_1_110001101110;
      patterns[36318] = 29'b1_000110111011_110_1_000110111011;
      patterns[36319] = 29'b1_000110111011_111_1_000110111011;
      patterns[36320] = 29'b1_000110111100_000_1_000110111100;
      patterns[36321] = 29'b1_000110111100_001_1_111100000110;
      patterns[36322] = 29'b1_000110111100_010_0_001101111001;
      patterns[36323] = 29'b1_000110111100_011_0_011011110010;
      patterns[36324] = 29'b1_000110111100_100_0_100011011110;
      patterns[36325] = 29'b1_000110111100_101_0_010001101111;
      patterns[36326] = 29'b1_000110111100_110_1_000110111100;
      patterns[36327] = 29'b1_000110111100_111_1_000110111100;
      patterns[36328] = 29'b1_000110111101_000_1_000110111101;
      patterns[36329] = 29'b1_000110111101_001_1_111101000110;
      patterns[36330] = 29'b1_000110111101_010_0_001101111011;
      patterns[36331] = 29'b1_000110111101_011_0_011011110110;
      patterns[36332] = 29'b1_000110111101_100_1_100011011110;
      patterns[36333] = 29'b1_000110111101_101_0_110001101111;
      patterns[36334] = 29'b1_000110111101_110_1_000110111101;
      patterns[36335] = 29'b1_000110111101_111_1_000110111101;
      patterns[36336] = 29'b1_000110111110_000_1_000110111110;
      patterns[36337] = 29'b1_000110111110_001_1_111110000110;
      patterns[36338] = 29'b1_000110111110_010_0_001101111101;
      patterns[36339] = 29'b1_000110111110_011_0_011011111010;
      patterns[36340] = 29'b1_000110111110_100_0_100011011111;
      patterns[36341] = 29'b1_000110111110_101_1_010001101111;
      patterns[36342] = 29'b1_000110111110_110_1_000110111110;
      patterns[36343] = 29'b1_000110111110_111_1_000110111110;
      patterns[36344] = 29'b1_000110111111_000_1_000110111111;
      patterns[36345] = 29'b1_000110111111_001_1_111111000110;
      patterns[36346] = 29'b1_000110111111_010_0_001101111111;
      patterns[36347] = 29'b1_000110111111_011_0_011011111110;
      patterns[36348] = 29'b1_000110111111_100_1_100011011111;
      patterns[36349] = 29'b1_000110111111_101_1_110001101111;
      patterns[36350] = 29'b1_000110111111_110_1_000110111111;
      patterns[36351] = 29'b1_000110111111_111_1_000110111111;
      patterns[36352] = 29'b1_000111000000_000_1_000111000000;
      patterns[36353] = 29'b1_000111000000_001_1_000000000111;
      patterns[36354] = 29'b1_000111000000_010_0_001110000001;
      patterns[36355] = 29'b1_000111000000_011_0_011100000010;
      patterns[36356] = 29'b1_000111000000_100_0_100011100000;
      patterns[36357] = 29'b1_000111000000_101_0_010001110000;
      patterns[36358] = 29'b1_000111000000_110_1_000111000000;
      patterns[36359] = 29'b1_000111000000_111_1_000111000000;
      patterns[36360] = 29'b1_000111000001_000_1_000111000001;
      patterns[36361] = 29'b1_000111000001_001_1_000001000111;
      patterns[36362] = 29'b1_000111000001_010_0_001110000011;
      patterns[36363] = 29'b1_000111000001_011_0_011100000110;
      patterns[36364] = 29'b1_000111000001_100_1_100011100000;
      patterns[36365] = 29'b1_000111000001_101_0_110001110000;
      patterns[36366] = 29'b1_000111000001_110_1_000111000001;
      patterns[36367] = 29'b1_000111000001_111_1_000111000001;
      patterns[36368] = 29'b1_000111000010_000_1_000111000010;
      patterns[36369] = 29'b1_000111000010_001_1_000010000111;
      patterns[36370] = 29'b1_000111000010_010_0_001110000101;
      patterns[36371] = 29'b1_000111000010_011_0_011100001010;
      patterns[36372] = 29'b1_000111000010_100_0_100011100001;
      patterns[36373] = 29'b1_000111000010_101_1_010001110000;
      patterns[36374] = 29'b1_000111000010_110_1_000111000010;
      patterns[36375] = 29'b1_000111000010_111_1_000111000010;
      patterns[36376] = 29'b1_000111000011_000_1_000111000011;
      patterns[36377] = 29'b1_000111000011_001_1_000011000111;
      patterns[36378] = 29'b1_000111000011_010_0_001110000111;
      patterns[36379] = 29'b1_000111000011_011_0_011100001110;
      patterns[36380] = 29'b1_000111000011_100_1_100011100001;
      patterns[36381] = 29'b1_000111000011_101_1_110001110000;
      patterns[36382] = 29'b1_000111000011_110_1_000111000011;
      patterns[36383] = 29'b1_000111000011_111_1_000111000011;
      patterns[36384] = 29'b1_000111000100_000_1_000111000100;
      patterns[36385] = 29'b1_000111000100_001_1_000100000111;
      patterns[36386] = 29'b1_000111000100_010_0_001110001001;
      patterns[36387] = 29'b1_000111000100_011_0_011100010010;
      patterns[36388] = 29'b1_000111000100_100_0_100011100010;
      patterns[36389] = 29'b1_000111000100_101_0_010001110001;
      patterns[36390] = 29'b1_000111000100_110_1_000111000100;
      patterns[36391] = 29'b1_000111000100_111_1_000111000100;
      patterns[36392] = 29'b1_000111000101_000_1_000111000101;
      patterns[36393] = 29'b1_000111000101_001_1_000101000111;
      patterns[36394] = 29'b1_000111000101_010_0_001110001011;
      patterns[36395] = 29'b1_000111000101_011_0_011100010110;
      patterns[36396] = 29'b1_000111000101_100_1_100011100010;
      patterns[36397] = 29'b1_000111000101_101_0_110001110001;
      patterns[36398] = 29'b1_000111000101_110_1_000111000101;
      patterns[36399] = 29'b1_000111000101_111_1_000111000101;
      patterns[36400] = 29'b1_000111000110_000_1_000111000110;
      patterns[36401] = 29'b1_000111000110_001_1_000110000111;
      patterns[36402] = 29'b1_000111000110_010_0_001110001101;
      patterns[36403] = 29'b1_000111000110_011_0_011100011010;
      patterns[36404] = 29'b1_000111000110_100_0_100011100011;
      patterns[36405] = 29'b1_000111000110_101_1_010001110001;
      patterns[36406] = 29'b1_000111000110_110_1_000111000110;
      patterns[36407] = 29'b1_000111000110_111_1_000111000110;
      patterns[36408] = 29'b1_000111000111_000_1_000111000111;
      patterns[36409] = 29'b1_000111000111_001_1_000111000111;
      patterns[36410] = 29'b1_000111000111_010_0_001110001111;
      patterns[36411] = 29'b1_000111000111_011_0_011100011110;
      patterns[36412] = 29'b1_000111000111_100_1_100011100011;
      patterns[36413] = 29'b1_000111000111_101_1_110001110001;
      patterns[36414] = 29'b1_000111000111_110_1_000111000111;
      patterns[36415] = 29'b1_000111000111_111_1_000111000111;
      patterns[36416] = 29'b1_000111001000_000_1_000111001000;
      patterns[36417] = 29'b1_000111001000_001_1_001000000111;
      patterns[36418] = 29'b1_000111001000_010_0_001110010001;
      patterns[36419] = 29'b1_000111001000_011_0_011100100010;
      patterns[36420] = 29'b1_000111001000_100_0_100011100100;
      patterns[36421] = 29'b1_000111001000_101_0_010001110010;
      patterns[36422] = 29'b1_000111001000_110_1_000111001000;
      patterns[36423] = 29'b1_000111001000_111_1_000111001000;
      patterns[36424] = 29'b1_000111001001_000_1_000111001001;
      patterns[36425] = 29'b1_000111001001_001_1_001001000111;
      patterns[36426] = 29'b1_000111001001_010_0_001110010011;
      patterns[36427] = 29'b1_000111001001_011_0_011100100110;
      patterns[36428] = 29'b1_000111001001_100_1_100011100100;
      patterns[36429] = 29'b1_000111001001_101_0_110001110010;
      patterns[36430] = 29'b1_000111001001_110_1_000111001001;
      patterns[36431] = 29'b1_000111001001_111_1_000111001001;
      patterns[36432] = 29'b1_000111001010_000_1_000111001010;
      patterns[36433] = 29'b1_000111001010_001_1_001010000111;
      patterns[36434] = 29'b1_000111001010_010_0_001110010101;
      patterns[36435] = 29'b1_000111001010_011_0_011100101010;
      patterns[36436] = 29'b1_000111001010_100_0_100011100101;
      patterns[36437] = 29'b1_000111001010_101_1_010001110010;
      patterns[36438] = 29'b1_000111001010_110_1_000111001010;
      patterns[36439] = 29'b1_000111001010_111_1_000111001010;
      patterns[36440] = 29'b1_000111001011_000_1_000111001011;
      patterns[36441] = 29'b1_000111001011_001_1_001011000111;
      patterns[36442] = 29'b1_000111001011_010_0_001110010111;
      patterns[36443] = 29'b1_000111001011_011_0_011100101110;
      patterns[36444] = 29'b1_000111001011_100_1_100011100101;
      patterns[36445] = 29'b1_000111001011_101_1_110001110010;
      patterns[36446] = 29'b1_000111001011_110_1_000111001011;
      patterns[36447] = 29'b1_000111001011_111_1_000111001011;
      patterns[36448] = 29'b1_000111001100_000_1_000111001100;
      patterns[36449] = 29'b1_000111001100_001_1_001100000111;
      patterns[36450] = 29'b1_000111001100_010_0_001110011001;
      patterns[36451] = 29'b1_000111001100_011_0_011100110010;
      patterns[36452] = 29'b1_000111001100_100_0_100011100110;
      patterns[36453] = 29'b1_000111001100_101_0_010001110011;
      patterns[36454] = 29'b1_000111001100_110_1_000111001100;
      patterns[36455] = 29'b1_000111001100_111_1_000111001100;
      patterns[36456] = 29'b1_000111001101_000_1_000111001101;
      patterns[36457] = 29'b1_000111001101_001_1_001101000111;
      patterns[36458] = 29'b1_000111001101_010_0_001110011011;
      patterns[36459] = 29'b1_000111001101_011_0_011100110110;
      patterns[36460] = 29'b1_000111001101_100_1_100011100110;
      patterns[36461] = 29'b1_000111001101_101_0_110001110011;
      patterns[36462] = 29'b1_000111001101_110_1_000111001101;
      patterns[36463] = 29'b1_000111001101_111_1_000111001101;
      patterns[36464] = 29'b1_000111001110_000_1_000111001110;
      patterns[36465] = 29'b1_000111001110_001_1_001110000111;
      patterns[36466] = 29'b1_000111001110_010_0_001110011101;
      patterns[36467] = 29'b1_000111001110_011_0_011100111010;
      patterns[36468] = 29'b1_000111001110_100_0_100011100111;
      patterns[36469] = 29'b1_000111001110_101_1_010001110011;
      patterns[36470] = 29'b1_000111001110_110_1_000111001110;
      patterns[36471] = 29'b1_000111001110_111_1_000111001110;
      patterns[36472] = 29'b1_000111001111_000_1_000111001111;
      patterns[36473] = 29'b1_000111001111_001_1_001111000111;
      patterns[36474] = 29'b1_000111001111_010_0_001110011111;
      patterns[36475] = 29'b1_000111001111_011_0_011100111110;
      patterns[36476] = 29'b1_000111001111_100_1_100011100111;
      patterns[36477] = 29'b1_000111001111_101_1_110001110011;
      patterns[36478] = 29'b1_000111001111_110_1_000111001111;
      patterns[36479] = 29'b1_000111001111_111_1_000111001111;
      patterns[36480] = 29'b1_000111010000_000_1_000111010000;
      patterns[36481] = 29'b1_000111010000_001_1_010000000111;
      patterns[36482] = 29'b1_000111010000_010_0_001110100001;
      patterns[36483] = 29'b1_000111010000_011_0_011101000010;
      patterns[36484] = 29'b1_000111010000_100_0_100011101000;
      patterns[36485] = 29'b1_000111010000_101_0_010001110100;
      patterns[36486] = 29'b1_000111010000_110_1_000111010000;
      patterns[36487] = 29'b1_000111010000_111_1_000111010000;
      patterns[36488] = 29'b1_000111010001_000_1_000111010001;
      patterns[36489] = 29'b1_000111010001_001_1_010001000111;
      patterns[36490] = 29'b1_000111010001_010_0_001110100011;
      patterns[36491] = 29'b1_000111010001_011_0_011101000110;
      patterns[36492] = 29'b1_000111010001_100_1_100011101000;
      patterns[36493] = 29'b1_000111010001_101_0_110001110100;
      patterns[36494] = 29'b1_000111010001_110_1_000111010001;
      patterns[36495] = 29'b1_000111010001_111_1_000111010001;
      patterns[36496] = 29'b1_000111010010_000_1_000111010010;
      patterns[36497] = 29'b1_000111010010_001_1_010010000111;
      patterns[36498] = 29'b1_000111010010_010_0_001110100101;
      patterns[36499] = 29'b1_000111010010_011_0_011101001010;
      patterns[36500] = 29'b1_000111010010_100_0_100011101001;
      patterns[36501] = 29'b1_000111010010_101_1_010001110100;
      patterns[36502] = 29'b1_000111010010_110_1_000111010010;
      patterns[36503] = 29'b1_000111010010_111_1_000111010010;
      patterns[36504] = 29'b1_000111010011_000_1_000111010011;
      patterns[36505] = 29'b1_000111010011_001_1_010011000111;
      patterns[36506] = 29'b1_000111010011_010_0_001110100111;
      patterns[36507] = 29'b1_000111010011_011_0_011101001110;
      patterns[36508] = 29'b1_000111010011_100_1_100011101001;
      patterns[36509] = 29'b1_000111010011_101_1_110001110100;
      patterns[36510] = 29'b1_000111010011_110_1_000111010011;
      patterns[36511] = 29'b1_000111010011_111_1_000111010011;
      patterns[36512] = 29'b1_000111010100_000_1_000111010100;
      patterns[36513] = 29'b1_000111010100_001_1_010100000111;
      patterns[36514] = 29'b1_000111010100_010_0_001110101001;
      patterns[36515] = 29'b1_000111010100_011_0_011101010010;
      patterns[36516] = 29'b1_000111010100_100_0_100011101010;
      patterns[36517] = 29'b1_000111010100_101_0_010001110101;
      patterns[36518] = 29'b1_000111010100_110_1_000111010100;
      patterns[36519] = 29'b1_000111010100_111_1_000111010100;
      patterns[36520] = 29'b1_000111010101_000_1_000111010101;
      patterns[36521] = 29'b1_000111010101_001_1_010101000111;
      patterns[36522] = 29'b1_000111010101_010_0_001110101011;
      patterns[36523] = 29'b1_000111010101_011_0_011101010110;
      patterns[36524] = 29'b1_000111010101_100_1_100011101010;
      patterns[36525] = 29'b1_000111010101_101_0_110001110101;
      patterns[36526] = 29'b1_000111010101_110_1_000111010101;
      patterns[36527] = 29'b1_000111010101_111_1_000111010101;
      patterns[36528] = 29'b1_000111010110_000_1_000111010110;
      patterns[36529] = 29'b1_000111010110_001_1_010110000111;
      patterns[36530] = 29'b1_000111010110_010_0_001110101101;
      patterns[36531] = 29'b1_000111010110_011_0_011101011010;
      patterns[36532] = 29'b1_000111010110_100_0_100011101011;
      patterns[36533] = 29'b1_000111010110_101_1_010001110101;
      patterns[36534] = 29'b1_000111010110_110_1_000111010110;
      patterns[36535] = 29'b1_000111010110_111_1_000111010110;
      patterns[36536] = 29'b1_000111010111_000_1_000111010111;
      patterns[36537] = 29'b1_000111010111_001_1_010111000111;
      patterns[36538] = 29'b1_000111010111_010_0_001110101111;
      patterns[36539] = 29'b1_000111010111_011_0_011101011110;
      patterns[36540] = 29'b1_000111010111_100_1_100011101011;
      patterns[36541] = 29'b1_000111010111_101_1_110001110101;
      patterns[36542] = 29'b1_000111010111_110_1_000111010111;
      patterns[36543] = 29'b1_000111010111_111_1_000111010111;
      patterns[36544] = 29'b1_000111011000_000_1_000111011000;
      patterns[36545] = 29'b1_000111011000_001_1_011000000111;
      patterns[36546] = 29'b1_000111011000_010_0_001110110001;
      patterns[36547] = 29'b1_000111011000_011_0_011101100010;
      patterns[36548] = 29'b1_000111011000_100_0_100011101100;
      patterns[36549] = 29'b1_000111011000_101_0_010001110110;
      patterns[36550] = 29'b1_000111011000_110_1_000111011000;
      patterns[36551] = 29'b1_000111011000_111_1_000111011000;
      patterns[36552] = 29'b1_000111011001_000_1_000111011001;
      patterns[36553] = 29'b1_000111011001_001_1_011001000111;
      patterns[36554] = 29'b1_000111011001_010_0_001110110011;
      patterns[36555] = 29'b1_000111011001_011_0_011101100110;
      patterns[36556] = 29'b1_000111011001_100_1_100011101100;
      patterns[36557] = 29'b1_000111011001_101_0_110001110110;
      patterns[36558] = 29'b1_000111011001_110_1_000111011001;
      patterns[36559] = 29'b1_000111011001_111_1_000111011001;
      patterns[36560] = 29'b1_000111011010_000_1_000111011010;
      patterns[36561] = 29'b1_000111011010_001_1_011010000111;
      patterns[36562] = 29'b1_000111011010_010_0_001110110101;
      patterns[36563] = 29'b1_000111011010_011_0_011101101010;
      patterns[36564] = 29'b1_000111011010_100_0_100011101101;
      patterns[36565] = 29'b1_000111011010_101_1_010001110110;
      patterns[36566] = 29'b1_000111011010_110_1_000111011010;
      patterns[36567] = 29'b1_000111011010_111_1_000111011010;
      patterns[36568] = 29'b1_000111011011_000_1_000111011011;
      patterns[36569] = 29'b1_000111011011_001_1_011011000111;
      patterns[36570] = 29'b1_000111011011_010_0_001110110111;
      patterns[36571] = 29'b1_000111011011_011_0_011101101110;
      patterns[36572] = 29'b1_000111011011_100_1_100011101101;
      patterns[36573] = 29'b1_000111011011_101_1_110001110110;
      patterns[36574] = 29'b1_000111011011_110_1_000111011011;
      patterns[36575] = 29'b1_000111011011_111_1_000111011011;
      patterns[36576] = 29'b1_000111011100_000_1_000111011100;
      patterns[36577] = 29'b1_000111011100_001_1_011100000111;
      patterns[36578] = 29'b1_000111011100_010_0_001110111001;
      patterns[36579] = 29'b1_000111011100_011_0_011101110010;
      patterns[36580] = 29'b1_000111011100_100_0_100011101110;
      patterns[36581] = 29'b1_000111011100_101_0_010001110111;
      patterns[36582] = 29'b1_000111011100_110_1_000111011100;
      patterns[36583] = 29'b1_000111011100_111_1_000111011100;
      patterns[36584] = 29'b1_000111011101_000_1_000111011101;
      patterns[36585] = 29'b1_000111011101_001_1_011101000111;
      patterns[36586] = 29'b1_000111011101_010_0_001110111011;
      patterns[36587] = 29'b1_000111011101_011_0_011101110110;
      patterns[36588] = 29'b1_000111011101_100_1_100011101110;
      patterns[36589] = 29'b1_000111011101_101_0_110001110111;
      patterns[36590] = 29'b1_000111011101_110_1_000111011101;
      patterns[36591] = 29'b1_000111011101_111_1_000111011101;
      patterns[36592] = 29'b1_000111011110_000_1_000111011110;
      patterns[36593] = 29'b1_000111011110_001_1_011110000111;
      patterns[36594] = 29'b1_000111011110_010_0_001110111101;
      patterns[36595] = 29'b1_000111011110_011_0_011101111010;
      patterns[36596] = 29'b1_000111011110_100_0_100011101111;
      patterns[36597] = 29'b1_000111011110_101_1_010001110111;
      patterns[36598] = 29'b1_000111011110_110_1_000111011110;
      patterns[36599] = 29'b1_000111011110_111_1_000111011110;
      patterns[36600] = 29'b1_000111011111_000_1_000111011111;
      patterns[36601] = 29'b1_000111011111_001_1_011111000111;
      patterns[36602] = 29'b1_000111011111_010_0_001110111111;
      patterns[36603] = 29'b1_000111011111_011_0_011101111110;
      patterns[36604] = 29'b1_000111011111_100_1_100011101111;
      patterns[36605] = 29'b1_000111011111_101_1_110001110111;
      patterns[36606] = 29'b1_000111011111_110_1_000111011111;
      patterns[36607] = 29'b1_000111011111_111_1_000111011111;
      patterns[36608] = 29'b1_000111100000_000_1_000111100000;
      patterns[36609] = 29'b1_000111100000_001_1_100000000111;
      patterns[36610] = 29'b1_000111100000_010_0_001111000001;
      patterns[36611] = 29'b1_000111100000_011_0_011110000010;
      patterns[36612] = 29'b1_000111100000_100_0_100011110000;
      patterns[36613] = 29'b1_000111100000_101_0_010001111000;
      patterns[36614] = 29'b1_000111100000_110_1_000111100000;
      patterns[36615] = 29'b1_000111100000_111_1_000111100000;
      patterns[36616] = 29'b1_000111100001_000_1_000111100001;
      patterns[36617] = 29'b1_000111100001_001_1_100001000111;
      patterns[36618] = 29'b1_000111100001_010_0_001111000011;
      patterns[36619] = 29'b1_000111100001_011_0_011110000110;
      patterns[36620] = 29'b1_000111100001_100_1_100011110000;
      patterns[36621] = 29'b1_000111100001_101_0_110001111000;
      patterns[36622] = 29'b1_000111100001_110_1_000111100001;
      patterns[36623] = 29'b1_000111100001_111_1_000111100001;
      patterns[36624] = 29'b1_000111100010_000_1_000111100010;
      patterns[36625] = 29'b1_000111100010_001_1_100010000111;
      patterns[36626] = 29'b1_000111100010_010_0_001111000101;
      patterns[36627] = 29'b1_000111100010_011_0_011110001010;
      patterns[36628] = 29'b1_000111100010_100_0_100011110001;
      patterns[36629] = 29'b1_000111100010_101_1_010001111000;
      patterns[36630] = 29'b1_000111100010_110_1_000111100010;
      patterns[36631] = 29'b1_000111100010_111_1_000111100010;
      patterns[36632] = 29'b1_000111100011_000_1_000111100011;
      patterns[36633] = 29'b1_000111100011_001_1_100011000111;
      patterns[36634] = 29'b1_000111100011_010_0_001111000111;
      patterns[36635] = 29'b1_000111100011_011_0_011110001110;
      patterns[36636] = 29'b1_000111100011_100_1_100011110001;
      patterns[36637] = 29'b1_000111100011_101_1_110001111000;
      patterns[36638] = 29'b1_000111100011_110_1_000111100011;
      patterns[36639] = 29'b1_000111100011_111_1_000111100011;
      patterns[36640] = 29'b1_000111100100_000_1_000111100100;
      patterns[36641] = 29'b1_000111100100_001_1_100100000111;
      patterns[36642] = 29'b1_000111100100_010_0_001111001001;
      patterns[36643] = 29'b1_000111100100_011_0_011110010010;
      patterns[36644] = 29'b1_000111100100_100_0_100011110010;
      patterns[36645] = 29'b1_000111100100_101_0_010001111001;
      patterns[36646] = 29'b1_000111100100_110_1_000111100100;
      patterns[36647] = 29'b1_000111100100_111_1_000111100100;
      patterns[36648] = 29'b1_000111100101_000_1_000111100101;
      patterns[36649] = 29'b1_000111100101_001_1_100101000111;
      patterns[36650] = 29'b1_000111100101_010_0_001111001011;
      patterns[36651] = 29'b1_000111100101_011_0_011110010110;
      patterns[36652] = 29'b1_000111100101_100_1_100011110010;
      patterns[36653] = 29'b1_000111100101_101_0_110001111001;
      patterns[36654] = 29'b1_000111100101_110_1_000111100101;
      patterns[36655] = 29'b1_000111100101_111_1_000111100101;
      patterns[36656] = 29'b1_000111100110_000_1_000111100110;
      patterns[36657] = 29'b1_000111100110_001_1_100110000111;
      patterns[36658] = 29'b1_000111100110_010_0_001111001101;
      patterns[36659] = 29'b1_000111100110_011_0_011110011010;
      patterns[36660] = 29'b1_000111100110_100_0_100011110011;
      patterns[36661] = 29'b1_000111100110_101_1_010001111001;
      patterns[36662] = 29'b1_000111100110_110_1_000111100110;
      patterns[36663] = 29'b1_000111100110_111_1_000111100110;
      patterns[36664] = 29'b1_000111100111_000_1_000111100111;
      patterns[36665] = 29'b1_000111100111_001_1_100111000111;
      patterns[36666] = 29'b1_000111100111_010_0_001111001111;
      patterns[36667] = 29'b1_000111100111_011_0_011110011110;
      patterns[36668] = 29'b1_000111100111_100_1_100011110011;
      patterns[36669] = 29'b1_000111100111_101_1_110001111001;
      patterns[36670] = 29'b1_000111100111_110_1_000111100111;
      patterns[36671] = 29'b1_000111100111_111_1_000111100111;
      patterns[36672] = 29'b1_000111101000_000_1_000111101000;
      patterns[36673] = 29'b1_000111101000_001_1_101000000111;
      patterns[36674] = 29'b1_000111101000_010_0_001111010001;
      patterns[36675] = 29'b1_000111101000_011_0_011110100010;
      patterns[36676] = 29'b1_000111101000_100_0_100011110100;
      patterns[36677] = 29'b1_000111101000_101_0_010001111010;
      patterns[36678] = 29'b1_000111101000_110_1_000111101000;
      patterns[36679] = 29'b1_000111101000_111_1_000111101000;
      patterns[36680] = 29'b1_000111101001_000_1_000111101001;
      patterns[36681] = 29'b1_000111101001_001_1_101001000111;
      patterns[36682] = 29'b1_000111101001_010_0_001111010011;
      patterns[36683] = 29'b1_000111101001_011_0_011110100110;
      patterns[36684] = 29'b1_000111101001_100_1_100011110100;
      patterns[36685] = 29'b1_000111101001_101_0_110001111010;
      patterns[36686] = 29'b1_000111101001_110_1_000111101001;
      patterns[36687] = 29'b1_000111101001_111_1_000111101001;
      patterns[36688] = 29'b1_000111101010_000_1_000111101010;
      patterns[36689] = 29'b1_000111101010_001_1_101010000111;
      patterns[36690] = 29'b1_000111101010_010_0_001111010101;
      patterns[36691] = 29'b1_000111101010_011_0_011110101010;
      patterns[36692] = 29'b1_000111101010_100_0_100011110101;
      patterns[36693] = 29'b1_000111101010_101_1_010001111010;
      patterns[36694] = 29'b1_000111101010_110_1_000111101010;
      patterns[36695] = 29'b1_000111101010_111_1_000111101010;
      patterns[36696] = 29'b1_000111101011_000_1_000111101011;
      patterns[36697] = 29'b1_000111101011_001_1_101011000111;
      patterns[36698] = 29'b1_000111101011_010_0_001111010111;
      patterns[36699] = 29'b1_000111101011_011_0_011110101110;
      patterns[36700] = 29'b1_000111101011_100_1_100011110101;
      patterns[36701] = 29'b1_000111101011_101_1_110001111010;
      patterns[36702] = 29'b1_000111101011_110_1_000111101011;
      patterns[36703] = 29'b1_000111101011_111_1_000111101011;
      patterns[36704] = 29'b1_000111101100_000_1_000111101100;
      patterns[36705] = 29'b1_000111101100_001_1_101100000111;
      patterns[36706] = 29'b1_000111101100_010_0_001111011001;
      patterns[36707] = 29'b1_000111101100_011_0_011110110010;
      patterns[36708] = 29'b1_000111101100_100_0_100011110110;
      patterns[36709] = 29'b1_000111101100_101_0_010001111011;
      patterns[36710] = 29'b1_000111101100_110_1_000111101100;
      patterns[36711] = 29'b1_000111101100_111_1_000111101100;
      patterns[36712] = 29'b1_000111101101_000_1_000111101101;
      patterns[36713] = 29'b1_000111101101_001_1_101101000111;
      patterns[36714] = 29'b1_000111101101_010_0_001111011011;
      patterns[36715] = 29'b1_000111101101_011_0_011110110110;
      patterns[36716] = 29'b1_000111101101_100_1_100011110110;
      patterns[36717] = 29'b1_000111101101_101_0_110001111011;
      patterns[36718] = 29'b1_000111101101_110_1_000111101101;
      patterns[36719] = 29'b1_000111101101_111_1_000111101101;
      patterns[36720] = 29'b1_000111101110_000_1_000111101110;
      patterns[36721] = 29'b1_000111101110_001_1_101110000111;
      patterns[36722] = 29'b1_000111101110_010_0_001111011101;
      patterns[36723] = 29'b1_000111101110_011_0_011110111010;
      patterns[36724] = 29'b1_000111101110_100_0_100011110111;
      patterns[36725] = 29'b1_000111101110_101_1_010001111011;
      patterns[36726] = 29'b1_000111101110_110_1_000111101110;
      patterns[36727] = 29'b1_000111101110_111_1_000111101110;
      patterns[36728] = 29'b1_000111101111_000_1_000111101111;
      patterns[36729] = 29'b1_000111101111_001_1_101111000111;
      patterns[36730] = 29'b1_000111101111_010_0_001111011111;
      patterns[36731] = 29'b1_000111101111_011_0_011110111110;
      patterns[36732] = 29'b1_000111101111_100_1_100011110111;
      patterns[36733] = 29'b1_000111101111_101_1_110001111011;
      patterns[36734] = 29'b1_000111101111_110_1_000111101111;
      patterns[36735] = 29'b1_000111101111_111_1_000111101111;
      patterns[36736] = 29'b1_000111110000_000_1_000111110000;
      patterns[36737] = 29'b1_000111110000_001_1_110000000111;
      patterns[36738] = 29'b1_000111110000_010_0_001111100001;
      patterns[36739] = 29'b1_000111110000_011_0_011111000010;
      patterns[36740] = 29'b1_000111110000_100_0_100011111000;
      patterns[36741] = 29'b1_000111110000_101_0_010001111100;
      patterns[36742] = 29'b1_000111110000_110_1_000111110000;
      patterns[36743] = 29'b1_000111110000_111_1_000111110000;
      patterns[36744] = 29'b1_000111110001_000_1_000111110001;
      patterns[36745] = 29'b1_000111110001_001_1_110001000111;
      patterns[36746] = 29'b1_000111110001_010_0_001111100011;
      patterns[36747] = 29'b1_000111110001_011_0_011111000110;
      patterns[36748] = 29'b1_000111110001_100_1_100011111000;
      patterns[36749] = 29'b1_000111110001_101_0_110001111100;
      patterns[36750] = 29'b1_000111110001_110_1_000111110001;
      patterns[36751] = 29'b1_000111110001_111_1_000111110001;
      patterns[36752] = 29'b1_000111110010_000_1_000111110010;
      patterns[36753] = 29'b1_000111110010_001_1_110010000111;
      patterns[36754] = 29'b1_000111110010_010_0_001111100101;
      patterns[36755] = 29'b1_000111110010_011_0_011111001010;
      patterns[36756] = 29'b1_000111110010_100_0_100011111001;
      patterns[36757] = 29'b1_000111110010_101_1_010001111100;
      patterns[36758] = 29'b1_000111110010_110_1_000111110010;
      patterns[36759] = 29'b1_000111110010_111_1_000111110010;
      patterns[36760] = 29'b1_000111110011_000_1_000111110011;
      patterns[36761] = 29'b1_000111110011_001_1_110011000111;
      patterns[36762] = 29'b1_000111110011_010_0_001111100111;
      patterns[36763] = 29'b1_000111110011_011_0_011111001110;
      patterns[36764] = 29'b1_000111110011_100_1_100011111001;
      patterns[36765] = 29'b1_000111110011_101_1_110001111100;
      patterns[36766] = 29'b1_000111110011_110_1_000111110011;
      patterns[36767] = 29'b1_000111110011_111_1_000111110011;
      patterns[36768] = 29'b1_000111110100_000_1_000111110100;
      patterns[36769] = 29'b1_000111110100_001_1_110100000111;
      patterns[36770] = 29'b1_000111110100_010_0_001111101001;
      patterns[36771] = 29'b1_000111110100_011_0_011111010010;
      patterns[36772] = 29'b1_000111110100_100_0_100011111010;
      patterns[36773] = 29'b1_000111110100_101_0_010001111101;
      patterns[36774] = 29'b1_000111110100_110_1_000111110100;
      patterns[36775] = 29'b1_000111110100_111_1_000111110100;
      patterns[36776] = 29'b1_000111110101_000_1_000111110101;
      patterns[36777] = 29'b1_000111110101_001_1_110101000111;
      patterns[36778] = 29'b1_000111110101_010_0_001111101011;
      patterns[36779] = 29'b1_000111110101_011_0_011111010110;
      patterns[36780] = 29'b1_000111110101_100_1_100011111010;
      patterns[36781] = 29'b1_000111110101_101_0_110001111101;
      patterns[36782] = 29'b1_000111110101_110_1_000111110101;
      patterns[36783] = 29'b1_000111110101_111_1_000111110101;
      patterns[36784] = 29'b1_000111110110_000_1_000111110110;
      patterns[36785] = 29'b1_000111110110_001_1_110110000111;
      patterns[36786] = 29'b1_000111110110_010_0_001111101101;
      patterns[36787] = 29'b1_000111110110_011_0_011111011010;
      patterns[36788] = 29'b1_000111110110_100_0_100011111011;
      patterns[36789] = 29'b1_000111110110_101_1_010001111101;
      patterns[36790] = 29'b1_000111110110_110_1_000111110110;
      patterns[36791] = 29'b1_000111110110_111_1_000111110110;
      patterns[36792] = 29'b1_000111110111_000_1_000111110111;
      patterns[36793] = 29'b1_000111110111_001_1_110111000111;
      patterns[36794] = 29'b1_000111110111_010_0_001111101111;
      patterns[36795] = 29'b1_000111110111_011_0_011111011110;
      patterns[36796] = 29'b1_000111110111_100_1_100011111011;
      patterns[36797] = 29'b1_000111110111_101_1_110001111101;
      patterns[36798] = 29'b1_000111110111_110_1_000111110111;
      patterns[36799] = 29'b1_000111110111_111_1_000111110111;
      patterns[36800] = 29'b1_000111111000_000_1_000111111000;
      patterns[36801] = 29'b1_000111111000_001_1_111000000111;
      patterns[36802] = 29'b1_000111111000_010_0_001111110001;
      patterns[36803] = 29'b1_000111111000_011_0_011111100010;
      patterns[36804] = 29'b1_000111111000_100_0_100011111100;
      patterns[36805] = 29'b1_000111111000_101_0_010001111110;
      patterns[36806] = 29'b1_000111111000_110_1_000111111000;
      patterns[36807] = 29'b1_000111111000_111_1_000111111000;
      patterns[36808] = 29'b1_000111111001_000_1_000111111001;
      patterns[36809] = 29'b1_000111111001_001_1_111001000111;
      patterns[36810] = 29'b1_000111111001_010_0_001111110011;
      patterns[36811] = 29'b1_000111111001_011_0_011111100110;
      patterns[36812] = 29'b1_000111111001_100_1_100011111100;
      patterns[36813] = 29'b1_000111111001_101_0_110001111110;
      patterns[36814] = 29'b1_000111111001_110_1_000111111001;
      patterns[36815] = 29'b1_000111111001_111_1_000111111001;
      patterns[36816] = 29'b1_000111111010_000_1_000111111010;
      patterns[36817] = 29'b1_000111111010_001_1_111010000111;
      patterns[36818] = 29'b1_000111111010_010_0_001111110101;
      patterns[36819] = 29'b1_000111111010_011_0_011111101010;
      patterns[36820] = 29'b1_000111111010_100_0_100011111101;
      patterns[36821] = 29'b1_000111111010_101_1_010001111110;
      patterns[36822] = 29'b1_000111111010_110_1_000111111010;
      patterns[36823] = 29'b1_000111111010_111_1_000111111010;
      patterns[36824] = 29'b1_000111111011_000_1_000111111011;
      patterns[36825] = 29'b1_000111111011_001_1_111011000111;
      patterns[36826] = 29'b1_000111111011_010_0_001111110111;
      patterns[36827] = 29'b1_000111111011_011_0_011111101110;
      patterns[36828] = 29'b1_000111111011_100_1_100011111101;
      patterns[36829] = 29'b1_000111111011_101_1_110001111110;
      patterns[36830] = 29'b1_000111111011_110_1_000111111011;
      patterns[36831] = 29'b1_000111111011_111_1_000111111011;
      patterns[36832] = 29'b1_000111111100_000_1_000111111100;
      patterns[36833] = 29'b1_000111111100_001_1_111100000111;
      patterns[36834] = 29'b1_000111111100_010_0_001111111001;
      patterns[36835] = 29'b1_000111111100_011_0_011111110010;
      patterns[36836] = 29'b1_000111111100_100_0_100011111110;
      patterns[36837] = 29'b1_000111111100_101_0_010001111111;
      patterns[36838] = 29'b1_000111111100_110_1_000111111100;
      patterns[36839] = 29'b1_000111111100_111_1_000111111100;
      patterns[36840] = 29'b1_000111111101_000_1_000111111101;
      patterns[36841] = 29'b1_000111111101_001_1_111101000111;
      patterns[36842] = 29'b1_000111111101_010_0_001111111011;
      patterns[36843] = 29'b1_000111111101_011_0_011111110110;
      patterns[36844] = 29'b1_000111111101_100_1_100011111110;
      patterns[36845] = 29'b1_000111111101_101_0_110001111111;
      patterns[36846] = 29'b1_000111111101_110_1_000111111101;
      patterns[36847] = 29'b1_000111111101_111_1_000111111101;
      patterns[36848] = 29'b1_000111111110_000_1_000111111110;
      patterns[36849] = 29'b1_000111111110_001_1_111110000111;
      patterns[36850] = 29'b1_000111111110_010_0_001111111101;
      patterns[36851] = 29'b1_000111111110_011_0_011111111010;
      patterns[36852] = 29'b1_000111111110_100_0_100011111111;
      patterns[36853] = 29'b1_000111111110_101_1_010001111111;
      patterns[36854] = 29'b1_000111111110_110_1_000111111110;
      patterns[36855] = 29'b1_000111111110_111_1_000111111110;
      patterns[36856] = 29'b1_000111111111_000_1_000111111111;
      patterns[36857] = 29'b1_000111111111_001_1_111111000111;
      patterns[36858] = 29'b1_000111111111_010_0_001111111111;
      patterns[36859] = 29'b1_000111111111_011_0_011111111110;
      patterns[36860] = 29'b1_000111111111_100_1_100011111111;
      patterns[36861] = 29'b1_000111111111_101_1_110001111111;
      patterns[36862] = 29'b1_000111111111_110_1_000111111111;
      patterns[36863] = 29'b1_000111111111_111_1_000111111111;
      patterns[36864] = 29'b1_001000000000_000_1_001000000000;
      patterns[36865] = 29'b1_001000000000_001_1_000000001000;
      patterns[36866] = 29'b1_001000000000_010_0_010000000001;
      patterns[36867] = 29'b1_001000000000_011_0_100000000010;
      patterns[36868] = 29'b1_001000000000_100_0_100100000000;
      patterns[36869] = 29'b1_001000000000_101_0_010010000000;
      patterns[36870] = 29'b1_001000000000_110_1_001000000000;
      patterns[36871] = 29'b1_001000000000_111_1_001000000000;
      patterns[36872] = 29'b1_001000000001_000_1_001000000001;
      patterns[36873] = 29'b1_001000000001_001_1_000001001000;
      patterns[36874] = 29'b1_001000000001_010_0_010000000011;
      patterns[36875] = 29'b1_001000000001_011_0_100000000110;
      patterns[36876] = 29'b1_001000000001_100_1_100100000000;
      patterns[36877] = 29'b1_001000000001_101_0_110010000000;
      patterns[36878] = 29'b1_001000000001_110_1_001000000001;
      patterns[36879] = 29'b1_001000000001_111_1_001000000001;
      patterns[36880] = 29'b1_001000000010_000_1_001000000010;
      patterns[36881] = 29'b1_001000000010_001_1_000010001000;
      patterns[36882] = 29'b1_001000000010_010_0_010000000101;
      patterns[36883] = 29'b1_001000000010_011_0_100000001010;
      patterns[36884] = 29'b1_001000000010_100_0_100100000001;
      patterns[36885] = 29'b1_001000000010_101_1_010010000000;
      patterns[36886] = 29'b1_001000000010_110_1_001000000010;
      patterns[36887] = 29'b1_001000000010_111_1_001000000010;
      patterns[36888] = 29'b1_001000000011_000_1_001000000011;
      patterns[36889] = 29'b1_001000000011_001_1_000011001000;
      patterns[36890] = 29'b1_001000000011_010_0_010000000111;
      patterns[36891] = 29'b1_001000000011_011_0_100000001110;
      patterns[36892] = 29'b1_001000000011_100_1_100100000001;
      patterns[36893] = 29'b1_001000000011_101_1_110010000000;
      patterns[36894] = 29'b1_001000000011_110_1_001000000011;
      patterns[36895] = 29'b1_001000000011_111_1_001000000011;
      patterns[36896] = 29'b1_001000000100_000_1_001000000100;
      patterns[36897] = 29'b1_001000000100_001_1_000100001000;
      patterns[36898] = 29'b1_001000000100_010_0_010000001001;
      patterns[36899] = 29'b1_001000000100_011_0_100000010010;
      patterns[36900] = 29'b1_001000000100_100_0_100100000010;
      patterns[36901] = 29'b1_001000000100_101_0_010010000001;
      patterns[36902] = 29'b1_001000000100_110_1_001000000100;
      patterns[36903] = 29'b1_001000000100_111_1_001000000100;
      patterns[36904] = 29'b1_001000000101_000_1_001000000101;
      patterns[36905] = 29'b1_001000000101_001_1_000101001000;
      patterns[36906] = 29'b1_001000000101_010_0_010000001011;
      patterns[36907] = 29'b1_001000000101_011_0_100000010110;
      patterns[36908] = 29'b1_001000000101_100_1_100100000010;
      patterns[36909] = 29'b1_001000000101_101_0_110010000001;
      patterns[36910] = 29'b1_001000000101_110_1_001000000101;
      patterns[36911] = 29'b1_001000000101_111_1_001000000101;
      patterns[36912] = 29'b1_001000000110_000_1_001000000110;
      patterns[36913] = 29'b1_001000000110_001_1_000110001000;
      patterns[36914] = 29'b1_001000000110_010_0_010000001101;
      patterns[36915] = 29'b1_001000000110_011_0_100000011010;
      patterns[36916] = 29'b1_001000000110_100_0_100100000011;
      patterns[36917] = 29'b1_001000000110_101_1_010010000001;
      patterns[36918] = 29'b1_001000000110_110_1_001000000110;
      patterns[36919] = 29'b1_001000000110_111_1_001000000110;
      patterns[36920] = 29'b1_001000000111_000_1_001000000111;
      patterns[36921] = 29'b1_001000000111_001_1_000111001000;
      patterns[36922] = 29'b1_001000000111_010_0_010000001111;
      patterns[36923] = 29'b1_001000000111_011_0_100000011110;
      patterns[36924] = 29'b1_001000000111_100_1_100100000011;
      patterns[36925] = 29'b1_001000000111_101_1_110010000001;
      patterns[36926] = 29'b1_001000000111_110_1_001000000111;
      patterns[36927] = 29'b1_001000000111_111_1_001000000111;
      patterns[36928] = 29'b1_001000001000_000_1_001000001000;
      patterns[36929] = 29'b1_001000001000_001_1_001000001000;
      patterns[36930] = 29'b1_001000001000_010_0_010000010001;
      patterns[36931] = 29'b1_001000001000_011_0_100000100010;
      patterns[36932] = 29'b1_001000001000_100_0_100100000100;
      patterns[36933] = 29'b1_001000001000_101_0_010010000010;
      patterns[36934] = 29'b1_001000001000_110_1_001000001000;
      patterns[36935] = 29'b1_001000001000_111_1_001000001000;
      patterns[36936] = 29'b1_001000001001_000_1_001000001001;
      patterns[36937] = 29'b1_001000001001_001_1_001001001000;
      patterns[36938] = 29'b1_001000001001_010_0_010000010011;
      patterns[36939] = 29'b1_001000001001_011_0_100000100110;
      patterns[36940] = 29'b1_001000001001_100_1_100100000100;
      patterns[36941] = 29'b1_001000001001_101_0_110010000010;
      patterns[36942] = 29'b1_001000001001_110_1_001000001001;
      patterns[36943] = 29'b1_001000001001_111_1_001000001001;
      patterns[36944] = 29'b1_001000001010_000_1_001000001010;
      patterns[36945] = 29'b1_001000001010_001_1_001010001000;
      patterns[36946] = 29'b1_001000001010_010_0_010000010101;
      patterns[36947] = 29'b1_001000001010_011_0_100000101010;
      patterns[36948] = 29'b1_001000001010_100_0_100100000101;
      patterns[36949] = 29'b1_001000001010_101_1_010010000010;
      patterns[36950] = 29'b1_001000001010_110_1_001000001010;
      patterns[36951] = 29'b1_001000001010_111_1_001000001010;
      patterns[36952] = 29'b1_001000001011_000_1_001000001011;
      patterns[36953] = 29'b1_001000001011_001_1_001011001000;
      patterns[36954] = 29'b1_001000001011_010_0_010000010111;
      patterns[36955] = 29'b1_001000001011_011_0_100000101110;
      patterns[36956] = 29'b1_001000001011_100_1_100100000101;
      patterns[36957] = 29'b1_001000001011_101_1_110010000010;
      patterns[36958] = 29'b1_001000001011_110_1_001000001011;
      patterns[36959] = 29'b1_001000001011_111_1_001000001011;
      patterns[36960] = 29'b1_001000001100_000_1_001000001100;
      patterns[36961] = 29'b1_001000001100_001_1_001100001000;
      patterns[36962] = 29'b1_001000001100_010_0_010000011001;
      patterns[36963] = 29'b1_001000001100_011_0_100000110010;
      patterns[36964] = 29'b1_001000001100_100_0_100100000110;
      patterns[36965] = 29'b1_001000001100_101_0_010010000011;
      patterns[36966] = 29'b1_001000001100_110_1_001000001100;
      patterns[36967] = 29'b1_001000001100_111_1_001000001100;
      patterns[36968] = 29'b1_001000001101_000_1_001000001101;
      patterns[36969] = 29'b1_001000001101_001_1_001101001000;
      patterns[36970] = 29'b1_001000001101_010_0_010000011011;
      patterns[36971] = 29'b1_001000001101_011_0_100000110110;
      patterns[36972] = 29'b1_001000001101_100_1_100100000110;
      patterns[36973] = 29'b1_001000001101_101_0_110010000011;
      patterns[36974] = 29'b1_001000001101_110_1_001000001101;
      patterns[36975] = 29'b1_001000001101_111_1_001000001101;
      patterns[36976] = 29'b1_001000001110_000_1_001000001110;
      patterns[36977] = 29'b1_001000001110_001_1_001110001000;
      patterns[36978] = 29'b1_001000001110_010_0_010000011101;
      patterns[36979] = 29'b1_001000001110_011_0_100000111010;
      patterns[36980] = 29'b1_001000001110_100_0_100100000111;
      patterns[36981] = 29'b1_001000001110_101_1_010010000011;
      patterns[36982] = 29'b1_001000001110_110_1_001000001110;
      patterns[36983] = 29'b1_001000001110_111_1_001000001110;
      patterns[36984] = 29'b1_001000001111_000_1_001000001111;
      patterns[36985] = 29'b1_001000001111_001_1_001111001000;
      patterns[36986] = 29'b1_001000001111_010_0_010000011111;
      patterns[36987] = 29'b1_001000001111_011_0_100000111110;
      patterns[36988] = 29'b1_001000001111_100_1_100100000111;
      patterns[36989] = 29'b1_001000001111_101_1_110010000011;
      patterns[36990] = 29'b1_001000001111_110_1_001000001111;
      patterns[36991] = 29'b1_001000001111_111_1_001000001111;
      patterns[36992] = 29'b1_001000010000_000_1_001000010000;
      patterns[36993] = 29'b1_001000010000_001_1_010000001000;
      patterns[36994] = 29'b1_001000010000_010_0_010000100001;
      patterns[36995] = 29'b1_001000010000_011_0_100001000010;
      patterns[36996] = 29'b1_001000010000_100_0_100100001000;
      patterns[36997] = 29'b1_001000010000_101_0_010010000100;
      patterns[36998] = 29'b1_001000010000_110_1_001000010000;
      patterns[36999] = 29'b1_001000010000_111_1_001000010000;
      patterns[37000] = 29'b1_001000010001_000_1_001000010001;
      patterns[37001] = 29'b1_001000010001_001_1_010001001000;
      patterns[37002] = 29'b1_001000010001_010_0_010000100011;
      patterns[37003] = 29'b1_001000010001_011_0_100001000110;
      patterns[37004] = 29'b1_001000010001_100_1_100100001000;
      patterns[37005] = 29'b1_001000010001_101_0_110010000100;
      patterns[37006] = 29'b1_001000010001_110_1_001000010001;
      patterns[37007] = 29'b1_001000010001_111_1_001000010001;
      patterns[37008] = 29'b1_001000010010_000_1_001000010010;
      patterns[37009] = 29'b1_001000010010_001_1_010010001000;
      patterns[37010] = 29'b1_001000010010_010_0_010000100101;
      patterns[37011] = 29'b1_001000010010_011_0_100001001010;
      patterns[37012] = 29'b1_001000010010_100_0_100100001001;
      patterns[37013] = 29'b1_001000010010_101_1_010010000100;
      patterns[37014] = 29'b1_001000010010_110_1_001000010010;
      patterns[37015] = 29'b1_001000010010_111_1_001000010010;
      patterns[37016] = 29'b1_001000010011_000_1_001000010011;
      patterns[37017] = 29'b1_001000010011_001_1_010011001000;
      patterns[37018] = 29'b1_001000010011_010_0_010000100111;
      patterns[37019] = 29'b1_001000010011_011_0_100001001110;
      patterns[37020] = 29'b1_001000010011_100_1_100100001001;
      patterns[37021] = 29'b1_001000010011_101_1_110010000100;
      patterns[37022] = 29'b1_001000010011_110_1_001000010011;
      patterns[37023] = 29'b1_001000010011_111_1_001000010011;
      patterns[37024] = 29'b1_001000010100_000_1_001000010100;
      patterns[37025] = 29'b1_001000010100_001_1_010100001000;
      patterns[37026] = 29'b1_001000010100_010_0_010000101001;
      patterns[37027] = 29'b1_001000010100_011_0_100001010010;
      patterns[37028] = 29'b1_001000010100_100_0_100100001010;
      patterns[37029] = 29'b1_001000010100_101_0_010010000101;
      patterns[37030] = 29'b1_001000010100_110_1_001000010100;
      patterns[37031] = 29'b1_001000010100_111_1_001000010100;
      patterns[37032] = 29'b1_001000010101_000_1_001000010101;
      patterns[37033] = 29'b1_001000010101_001_1_010101001000;
      patterns[37034] = 29'b1_001000010101_010_0_010000101011;
      patterns[37035] = 29'b1_001000010101_011_0_100001010110;
      patterns[37036] = 29'b1_001000010101_100_1_100100001010;
      patterns[37037] = 29'b1_001000010101_101_0_110010000101;
      patterns[37038] = 29'b1_001000010101_110_1_001000010101;
      patterns[37039] = 29'b1_001000010101_111_1_001000010101;
      patterns[37040] = 29'b1_001000010110_000_1_001000010110;
      patterns[37041] = 29'b1_001000010110_001_1_010110001000;
      patterns[37042] = 29'b1_001000010110_010_0_010000101101;
      patterns[37043] = 29'b1_001000010110_011_0_100001011010;
      patterns[37044] = 29'b1_001000010110_100_0_100100001011;
      patterns[37045] = 29'b1_001000010110_101_1_010010000101;
      patterns[37046] = 29'b1_001000010110_110_1_001000010110;
      patterns[37047] = 29'b1_001000010110_111_1_001000010110;
      patterns[37048] = 29'b1_001000010111_000_1_001000010111;
      patterns[37049] = 29'b1_001000010111_001_1_010111001000;
      patterns[37050] = 29'b1_001000010111_010_0_010000101111;
      patterns[37051] = 29'b1_001000010111_011_0_100001011110;
      patterns[37052] = 29'b1_001000010111_100_1_100100001011;
      patterns[37053] = 29'b1_001000010111_101_1_110010000101;
      patterns[37054] = 29'b1_001000010111_110_1_001000010111;
      patterns[37055] = 29'b1_001000010111_111_1_001000010111;
      patterns[37056] = 29'b1_001000011000_000_1_001000011000;
      patterns[37057] = 29'b1_001000011000_001_1_011000001000;
      patterns[37058] = 29'b1_001000011000_010_0_010000110001;
      patterns[37059] = 29'b1_001000011000_011_0_100001100010;
      patterns[37060] = 29'b1_001000011000_100_0_100100001100;
      patterns[37061] = 29'b1_001000011000_101_0_010010000110;
      patterns[37062] = 29'b1_001000011000_110_1_001000011000;
      patterns[37063] = 29'b1_001000011000_111_1_001000011000;
      patterns[37064] = 29'b1_001000011001_000_1_001000011001;
      patterns[37065] = 29'b1_001000011001_001_1_011001001000;
      patterns[37066] = 29'b1_001000011001_010_0_010000110011;
      patterns[37067] = 29'b1_001000011001_011_0_100001100110;
      patterns[37068] = 29'b1_001000011001_100_1_100100001100;
      patterns[37069] = 29'b1_001000011001_101_0_110010000110;
      patterns[37070] = 29'b1_001000011001_110_1_001000011001;
      patterns[37071] = 29'b1_001000011001_111_1_001000011001;
      patterns[37072] = 29'b1_001000011010_000_1_001000011010;
      patterns[37073] = 29'b1_001000011010_001_1_011010001000;
      patterns[37074] = 29'b1_001000011010_010_0_010000110101;
      patterns[37075] = 29'b1_001000011010_011_0_100001101010;
      patterns[37076] = 29'b1_001000011010_100_0_100100001101;
      patterns[37077] = 29'b1_001000011010_101_1_010010000110;
      patterns[37078] = 29'b1_001000011010_110_1_001000011010;
      patterns[37079] = 29'b1_001000011010_111_1_001000011010;
      patterns[37080] = 29'b1_001000011011_000_1_001000011011;
      patterns[37081] = 29'b1_001000011011_001_1_011011001000;
      patterns[37082] = 29'b1_001000011011_010_0_010000110111;
      patterns[37083] = 29'b1_001000011011_011_0_100001101110;
      patterns[37084] = 29'b1_001000011011_100_1_100100001101;
      patterns[37085] = 29'b1_001000011011_101_1_110010000110;
      patterns[37086] = 29'b1_001000011011_110_1_001000011011;
      patterns[37087] = 29'b1_001000011011_111_1_001000011011;
      patterns[37088] = 29'b1_001000011100_000_1_001000011100;
      patterns[37089] = 29'b1_001000011100_001_1_011100001000;
      patterns[37090] = 29'b1_001000011100_010_0_010000111001;
      patterns[37091] = 29'b1_001000011100_011_0_100001110010;
      patterns[37092] = 29'b1_001000011100_100_0_100100001110;
      patterns[37093] = 29'b1_001000011100_101_0_010010000111;
      patterns[37094] = 29'b1_001000011100_110_1_001000011100;
      patterns[37095] = 29'b1_001000011100_111_1_001000011100;
      patterns[37096] = 29'b1_001000011101_000_1_001000011101;
      patterns[37097] = 29'b1_001000011101_001_1_011101001000;
      patterns[37098] = 29'b1_001000011101_010_0_010000111011;
      patterns[37099] = 29'b1_001000011101_011_0_100001110110;
      patterns[37100] = 29'b1_001000011101_100_1_100100001110;
      patterns[37101] = 29'b1_001000011101_101_0_110010000111;
      patterns[37102] = 29'b1_001000011101_110_1_001000011101;
      patterns[37103] = 29'b1_001000011101_111_1_001000011101;
      patterns[37104] = 29'b1_001000011110_000_1_001000011110;
      patterns[37105] = 29'b1_001000011110_001_1_011110001000;
      patterns[37106] = 29'b1_001000011110_010_0_010000111101;
      patterns[37107] = 29'b1_001000011110_011_0_100001111010;
      patterns[37108] = 29'b1_001000011110_100_0_100100001111;
      patterns[37109] = 29'b1_001000011110_101_1_010010000111;
      patterns[37110] = 29'b1_001000011110_110_1_001000011110;
      patterns[37111] = 29'b1_001000011110_111_1_001000011110;
      patterns[37112] = 29'b1_001000011111_000_1_001000011111;
      patterns[37113] = 29'b1_001000011111_001_1_011111001000;
      patterns[37114] = 29'b1_001000011111_010_0_010000111111;
      patterns[37115] = 29'b1_001000011111_011_0_100001111110;
      patterns[37116] = 29'b1_001000011111_100_1_100100001111;
      patterns[37117] = 29'b1_001000011111_101_1_110010000111;
      patterns[37118] = 29'b1_001000011111_110_1_001000011111;
      patterns[37119] = 29'b1_001000011111_111_1_001000011111;
      patterns[37120] = 29'b1_001000100000_000_1_001000100000;
      patterns[37121] = 29'b1_001000100000_001_1_100000001000;
      patterns[37122] = 29'b1_001000100000_010_0_010001000001;
      patterns[37123] = 29'b1_001000100000_011_0_100010000010;
      patterns[37124] = 29'b1_001000100000_100_0_100100010000;
      patterns[37125] = 29'b1_001000100000_101_0_010010001000;
      patterns[37126] = 29'b1_001000100000_110_1_001000100000;
      patterns[37127] = 29'b1_001000100000_111_1_001000100000;
      patterns[37128] = 29'b1_001000100001_000_1_001000100001;
      patterns[37129] = 29'b1_001000100001_001_1_100001001000;
      patterns[37130] = 29'b1_001000100001_010_0_010001000011;
      patterns[37131] = 29'b1_001000100001_011_0_100010000110;
      patterns[37132] = 29'b1_001000100001_100_1_100100010000;
      patterns[37133] = 29'b1_001000100001_101_0_110010001000;
      patterns[37134] = 29'b1_001000100001_110_1_001000100001;
      patterns[37135] = 29'b1_001000100001_111_1_001000100001;
      patterns[37136] = 29'b1_001000100010_000_1_001000100010;
      patterns[37137] = 29'b1_001000100010_001_1_100010001000;
      patterns[37138] = 29'b1_001000100010_010_0_010001000101;
      patterns[37139] = 29'b1_001000100010_011_0_100010001010;
      patterns[37140] = 29'b1_001000100010_100_0_100100010001;
      patterns[37141] = 29'b1_001000100010_101_1_010010001000;
      patterns[37142] = 29'b1_001000100010_110_1_001000100010;
      patterns[37143] = 29'b1_001000100010_111_1_001000100010;
      patterns[37144] = 29'b1_001000100011_000_1_001000100011;
      patterns[37145] = 29'b1_001000100011_001_1_100011001000;
      patterns[37146] = 29'b1_001000100011_010_0_010001000111;
      patterns[37147] = 29'b1_001000100011_011_0_100010001110;
      patterns[37148] = 29'b1_001000100011_100_1_100100010001;
      patterns[37149] = 29'b1_001000100011_101_1_110010001000;
      patterns[37150] = 29'b1_001000100011_110_1_001000100011;
      patterns[37151] = 29'b1_001000100011_111_1_001000100011;
      patterns[37152] = 29'b1_001000100100_000_1_001000100100;
      patterns[37153] = 29'b1_001000100100_001_1_100100001000;
      patterns[37154] = 29'b1_001000100100_010_0_010001001001;
      patterns[37155] = 29'b1_001000100100_011_0_100010010010;
      patterns[37156] = 29'b1_001000100100_100_0_100100010010;
      patterns[37157] = 29'b1_001000100100_101_0_010010001001;
      patterns[37158] = 29'b1_001000100100_110_1_001000100100;
      patterns[37159] = 29'b1_001000100100_111_1_001000100100;
      patterns[37160] = 29'b1_001000100101_000_1_001000100101;
      patterns[37161] = 29'b1_001000100101_001_1_100101001000;
      patterns[37162] = 29'b1_001000100101_010_0_010001001011;
      patterns[37163] = 29'b1_001000100101_011_0_100010010110;
      patterns[37164] = 29'b1_001000100101_100_1_100100010010;
      patterns[37165] = 29'b1_001000100101_101_0_110010001001;
      patterns[37166] = 29'b1_001000100101_110_1_001000100101;
      patterns[37167] = 29'b1_001000100101_111_1_001000100101;
      patterns[37168] = 29'b1_001000100110_000_1_001000100110;
      patterns[37169] = 29'b1_001000100110_001_1_100110001000;
      patterns[37170] = 29'b1_001000100110_010_0_010001001101;
      patterns[37171] = 29'b1_001000100110_011_0_100010011010;
      patterns[37172] = 29'b1_001000100110_100_0_100100010011;
      patterns[37173] = 29'b1_001000100110_101_1_010010001001;
      patterns[37174] = 29'b1_001000100110_110_1_001000100110;
      patterns[37175] = 29'b1_001000100110_111_1_001000100110;
      patterns[37176] = 29'b1_001000100111_000_1_001000100111;
      patterns[37177] = 29'b1_001000100111_001_1_100111001000;
      patterns[37178] = 29'b1_001000100111_010_0_010001001111;
      patterns[37179] = 29'b1_001000100111_011_0_100010011110;
      patterns[37180] = 29'b1_001000100111_100_1_100100010011;
      patterns[37181] = 29'b1_001000100111_101_1_110010001001;
      patterns[37182] = 29'b1_001000100111_110_1_001000100111;
      patterns[37183] = 29'b1_001000100111_111_1_001000100111;
      patterns[37184] = 29'b1_001000101000_000_1_001000101000;
      patterns[37185] = 29'b1_001000101000_001_1_101000001000;
      patterns[37186] = 29'b1_001000101000_010_0_010001010001;
      patterns[37187] = 29'b1_001000101000_011_0_100010100010;
      patterns[37188] = 29'b1_001000101000_100_0_100100010100;
      patterns[37189] = 29'b1_001000101000_101_0_010010001010;
      patterns[37190] = 29'b1_001000101000_110_1_001000101000;
      patterns[37191] = 29'b1_001000101000_111_1_001000101000;
      patterns[37192] = 29'b1_001000101001_000_1_001000101001;
      patterns[37193] = 29'b1_001000101001_001_1_101001001000;
      patterns[37194] = 29'b1_001000101001_010_0_010001010011;
      patterns[37195] = 29'b1_001000101001_011_0_100010100110;
      patterns[37196] = 29'b1_001000101001_100_1_100100010100;
      patterns[37197] = 29'b1_001000101001_101_0_110010001010;
      patterns[37198] = 29'b1_001000101001_110_1_001000101001;
      patterns[37199] = 29'b1_001000101001_111_1_001000101001;
      patterns[37200] = 29'b1_001000101010_000_1_001000101010;
      patterns[37201] = 29'b1_001000101010_001_1_101010001000;
      patterns[37202] = 29'b1_001000101010_010_0_010001010101;
      patterns[37203] = 29'b1_001000101010_011_0_100010101010;
      patterns[37204] = 29'b1_001000101010_100_0_100100010101;
      patterns[37205] = 29'b1_001000101010_101_1_010010001010;
      patterns[37206] = 29'b1_001000101010_110_1_001000101010;
      patterns[37207] = 29'b1_001000101010_111_1_001000101010;
      patterns[37208] = 29'b1_001000101011_000_1_001000101011;
      patterns[37209] = 29'b1_001000101011_001_1_101011001000;
      patterns[37210] = 29'b1_001000101011_010_0_010001010111;
      patterns[37211] = 29'b1_001000101011_011_0_100010101110;
      patterns[37212] = 29'b1_001000101011_100_1_100100010101;
      patterns[37213] = 29'b1_001000101011_101_1_110010001010;
      patterns[37214] = 29'b1_001000101011_110_1_001000101011;
      patterns[37215] = 29'b1_001000101011_111_1_001000101011;
      patterns[37216] = 29'b1_001000101100_000_1_001000101100;
      patterns[37217] = 29'b1_001000101100_001_1_101100001000;
      patterns[37218] = 29'b1_001000101100_010_0_010001011001;
      patterns[37219] = 29'b1_001000101100_011_0_100010110010;
      patterns[37220] = 29'b1_001000101100_100_0_100100010110;
      patterns[37221] = 29'b1_001000101100_101_0_010010001011;
      patterns[37222] = 29'b1_001000101100_110_1_001000101100;
      patterns[37223] = 29'b1_001000101100_111_1_001000101100;
      patterns[37224] = 29'b1_001000101101_000_1_001000101101;
      patterns[37225] = 29'b1_001000101101_001_1_101101001000;
      patterns[37226] = 29'b1_001000101101_010_0_010001011011;
      patterns[37227] = 29'b1_001000101101_011_0_100010110110;
      patterns[37228] = 29'b1_001000101101_100_1_100100010110;
      patterns[37229] = 29'b1_001000101101_101_0_110010001011;
      patterns[37230] = 29'b1_001000101101_110_1_001000101101;
      patterns[37231] = 29'b1_001000101101_111_1_001000101101;
      patterns[37232] = 29'b1_001000101110_000_1_001000101110;
      patterns[37233] = 29'b1_001000101110_001_1_101110001000;
      patterns[37234] = 29'b1_001000101110_010_0_010001011101;
      patterns[37235] = 29'b1_001000101110_011_0_100010111010;
      patterns[37236] = 29'b1_001000101110_100_0_100100010111;
      patterns[37237] = 29'b1_001000101110_101_1_010010001011;
      patterns[37238] = 29'b1_001000101110_110_1_001000101110;
      patterns[37239] = 29'b1_001000101110_111_1_001000101110;
      patterns[37240] = 29'b1_001000101111_000_1_001000101111;
      patterns[37241] = 29'b1_001000101111_001_1_101111001000;
      patterns[37242] = 29'b1_001000101111_010_0_010001011111;
      patterns[37243] = 29'b1_001000101111_011_0_100010111110;
      patterns[37244] = 29'b1_001000101111_100_1_100100010111;
      patterns[37245] = 29'b1_001000101111_101_1_110010001011;
      patterns[37246] = 29'b1_001000101111_110_1_001000101111;
      patterns[37247] = 29'b1_001000101111_111_1_001000101111;
      patterns[37248] = 29'b1_001000110000_000_1_001000110000;
      patterns[37249] = 29'b1_001000110000_001_1_110000001000;
      patterns[37250] = 29'b1_001000110000_010_0_010001100001;
      patterns[37251] = 29'b1_001000110000_011_0_100011000010;
      patterns[37252] = 29'b1_001000110000_100_0_100100011000;
      patterns[37253] = 29'b1_001000110000_101_0_010010001100;
      patterns[37254] = 29'b1_001000110000_110_1_001000110000;
      patterns[37255] = 29'b1_001000110000_111_1_001000110000;
      patterns[37256] = 29'b1_001000110001_000_1_001000110001;
      patterns[37257] = 29'b1_001000110001_001_1_110001001000;
      patterns[37258] = 29'b1_001000110001_010_0_010001100011;
      patterns[37259] = 29'b1_001000110001_011_0_100011000110;
      patterns[37260] = 29'b1_001000110001_100_1_100100011000;
      patterns[37261] = 29'b1_001000110001_101_0_110010001100;
      patterns[37262] = 29'b1_001000110001_110_1_001000110001;
      patterns[37263] = 29'b1_001000110001_111_1_001000110001;
      patterns[37264] = 29'b1_001000110010_000_1_001000110010;
      patterns[37265] = 29'b1_001000110010_001_1_110010001000;
      patterns[37266] = 29'b1_001000110010_010_0_010001100101;
      patterns[37267] = 29'b1_001000110010_011_0_100011001010;
      patterns[37268] = 29'b1_001000110010_100_0_100100011001;
      patterns[37269] = 29'b1_001000110010_101_1_010010001100;
      patterns[37270] = 29'b1_001000110010_110_1_001000110010;
      patterns[37271] = 29'b1_001000110010_111_1_001000110010;
      patterns[37272] = 29'b1_001000110011_000_1_001000110011;
      patterns[37273] = 29'b1_001000110011_001_1_110011001000;
      patterns[37274] = 29'b1_001000110011_010_0_010001100111;
      patterns[37275] = 29'b1_001000110011_011_0_100011001110;
      patterns[37276] = 29'b1_001000110011_100_1_100100011001;
      patterns[37277] = 29'b1_001000110011_101_1_110010001100;
      patterns[37278] = 29'b1_001000110011_110_1_001000110011;
      patterns[37279] = 29'b1_001000110011_111_1_001000110011;
      patterns[37280] = 29'b1_001000110100_000_1_001000110100;
      patterns[37281] = 29'b1_001000110100_001_1_110100001000;
      patterns[37282] = 29'b1_001000110100_010_0_010001101001;
      patterns[37283] = 29'b1_001000110100_011_0_100011010010;
      patterns[37284] = 29'b1_001000110100_100_0_100100011010;
      patterns[37285] = 29'b1_001000110100_101_0_010010001101;
      patterns[37286] = 29'b1_001000110100_110_1_001000110100;
      patterns[37287] = 29'b1_001000110100_111_1_001000110100;
      patterns[37288] = 29'b1_001000110101_000_1_001000110101;
      patterns[37289] = 29'b1_001000110101_001_1_110101001000;
      patterns[37290] = 29'b1_001000110101_010_0_010001101011;
      patterns[37291] = 29'b1_001000110101_011_0_100011010110;
      patterns[37292] = 29'b1_001000110101_100_1_100100011010;
      patterns[37293] = 29'b1_001000110101_101_0_110010001101;
      patterns[37294] = 29'b1_001000110101_110_1_001000110101;
      patterns[37295] = 29'b1_001000110101_111_1_001000110101;
      patterns[37296] = 29'b1_001000110110_000_1_001000110110;
      patterns[37297] = 29'b1_001000110110_001_1_110110001000;
      patterns[37298] = 29'b1_001000110110_010_0_010001101101;
      patterns[37299] = 29'b1_001000110110_011_0_100011011010;
      patterns[37300] = 29'b1_001000110110_100_0_100100011011;
      patterns[37301] = 29'b1_001000110110_101_1_010010001101;
      patterns[37302] = 29'b1_001000110110_110_1_001000110110;
      patterns[37303] = 29'b1_001000110110_111_1_001000110110;
      patterns[37304] = 29'b1_001000110111_000_1_001000110111;
      patterns[37305] = 29'b1_001000110111_001_1_110111001000;
      patterns[37306] = 29'b1_001000110111_010_0_010001101111;
      patterns[37307] = 29'b1_001000110111_011_0_100011011110;
      patterns[37308] = 29'b1_001000110111_100_1_100100011011;
      patterns[37309] = 29'b1_001000110111_101_1_110010001101;
      patterns[37310] = 29'b1_001000110111_110_1_001000110111;
      patterns[37311] = 29'b1_001000110111_111_1_001000110111;
      patterns[37312] = 29'b1_001000111000_000_1_001000111000;
      patterns[37313] = 29'b1_001000111000_001_1_111000001000;
      patterns[37314] = 29'b1_001000111000_010_0_010001110001;
      patterns[37315] = 29'b1_001000111000_011_0_100011100010;
      patterns[37316] = 29'b1_001000111000_100_0_100100011100;
      patterns[37317] = 29'b1_001000111000_101_0_010010001110;
      patterns[37318] = 29'b1_001000111000_110_1_001000111000;
      patterns[37319] = 29'b1_001000111000_111_1_001000111000;
      patterns[37320] = 29'b1_001000111001_000_1_001000111001;
      patterns[37321] = 29'b1_001000111001_001_1_111001001000;
      patterns[37322] = 29'b1_001000111001_010_0_010001110011;
      patterns[37323] = 29'b1_001000111001_011_0_100011100110;
      patterns[37324] = 29'b1_001000111001_100_1_100100011100;
      patterns[37325] = 29'b1_001000111001_101_0_110010001110;
      patterns[37326] = 29'b1_001000111001_110_1_001000111001;
      patterns[37327] = 29'b1_001000111001_111_1_001000111001;
      patterns[37328] = 29'b1_001000111010_000_1_001000111010;
      patterns[37329] = 29'b1_001000111010_001_1_111010001000;
      patterns[37330] = 29'b1_001000111010_010_0_010001110101;
      patterns[37331] = 29'b1_001000111010_011_0_100011101010;
      patterns[37332] = 29'b1_001000111010_100_0_100100011101;
      patterns[37333] = 29'b1_001000111010_101_1_010010001110;
      patterns[37334] = 29'b1_001000111010_110_1_001000111010;
      patterns[37335] = 29'b1_001000111010_111_1_001000111010;
      patterns[37336] = 29'b1_001000111011_000_1_001000111011;
      patterns[37337] = 29'b1_001000111011_001_1_111011001000;
      patterns[37338] = 29'b1_001000111011_010_0_010001110111;
      patterns[37339] = 29'b1_001000111011_011_0_100011101110;
      patterns[37340] = 29'b1_001000111011_100_1_100100011101;
      patterns[37341] = 29'b1_001000111011_101_1_110010001110;
      patterns[37342] = 29'b1_001000111011_110_1_001000111011;
      patterns[37343] = 29'b1_001000111011_111_1_001000111011;
      patterns[37344] = 29'b1_001000111100_000_1_001000111100;
      patterns[37345] = 29'b1_001000111100_001_1_111100001000;
      patterns[37346] = 29'b1_001000111100_010_0_010001111001;
      patterns[37347] = 29'b1_001000111100_011_0_100011110010;
      patterns[37348] = 29'b1_001000111100_100_0_100100011110;
      patterns[37349] = 29'b1_001000111100_101_0_010010001111;
      patterns[37350] = 29'b1_001000111100_110_1_001000111100;
      patterns[37351] = 29'b1_001000111100_111_1_001000111100;
      patterns[37352] = 29'b1_001000111101_000_1_001000111101;
      patterns[37353] = 29'b1_001000111101_001_1_111101001000;
      patterns[37354] = 29'b1_001000111101_010_0_010001111011;
      patterns[37355] = 29'b1_001000111101_011_0_100011110110;
      patterns[37356] = 29'b1_001000111101_100_1_100100011110;
      patterns[37357] = 29'b1_001000111101_101_0_110010001111;
      patterns[37358] = 29'b1_001000111101_110_1_001000111101;
      patterns[37359] = 29'b1_001000111101_111_1_001000111101;
      patterns[37360] = 29'b1_001000111110_000_1_001000111110;
      patterns[37361] = 29'b1_001000111110_001_1_111110001000;
      patterns[37362] = 29'b1_001000111110_010_0_010001111101;
      patterns[37363] = 29'b1_001000111110_011_0_100011111010;
      patterns[37364] = 29'b1_001000111110_100_0_100100011111;
      patterns[37365] = 29'b1_001000111110_101_1_010010001111;
      patterns[37366] = 29'b1_001000111110_110_1_001000111110;
      patterns[37367] = 29'b1_001000111110_111_1_001000111110;
      patterns[37368] = 29'b1_001000111111_000_1_001000111111;
      patterns[37369] = 29'b1_001000111111_001_1_111111001000;
      patterns[37370] = 29'b1_001000111111_010_0_010001111111;
      patterns[37371] = 29'b1_001000111111_011_0_100011111110;
      patterns[37372] = 29'b1_001000111111_100_1_100100011111;
      patterns[37373] = 29'b1_001000111111_101_1_110010001111;
      patterns[37374] = 29'b1_001000111111_110_1_001000111111;
      patterns[37375] = 29'b1_001000111111_111_1_001000111111;
      patterns[37376] = 29'b1_001001000000_000_1_001001000000;
      patterns[37377] = 29'b1_001001000000_001_1_000000001001;
      patterns[37378] = 29'b1_001001000000_010_0_010010000001;
      patterns[37379] = 29'b1_001001000000_011_0_100100000010;
      patterns[37380] = 29'b1_001001000000_100_0_100100100000;
      patterns[37381] = 29'b1_001001000000_101_0_010010010000;
      patterns[37382] = 29'b1_001001000000_110_1_001001000000;
      patterns[37383] = 29'b1_001001000000_111_1_001001000000;
      patterns[37384] = 29'b1_001001000001_000_1_001001000001;
      patterns[37385] = 29'b1_001001000001_001_1_000001001001;
      patterns[37386] = 29'b1_001001000001_010_0_010010000011;
      patterns[37387] = 29'b1_001001000001_011_0_100100000110;
      patterns[37388] = 29'b1_001001000001_100_1_100100100000;
      patterns[37389] = 29'b1_001001000001_101_0_110010010000;
      patterns[37390] = 29'b1_001001000001_110_1_001001000001;
      patterns[37391] = 29'b1_001001000001_111_1_001001000001;
      patterns[37392] = 29'b1_001001000010_000_1_001001000010;
      patterns[37393] = 29'b1_001001000010_001_1_000010001001;
      patterns[37394] = 29'b1_001001000010_010_0_010010000101;
      patterns[37395] = 29'b1_001001000010_011_0_100100001010;
      patterns[37396] = 29'b1_001001000010_100_0_100100100001;
      patterns[37397] = 29'b1_001001000010_101_1_010010010000;
      patterns[37398] = 29'b1_001001000010_110_1_001001000010;
      patterns[37399] = 29'b1_001001000010_111_1_001001000010;
      patterns[37400] = 29'b1_001001000011_000_1_001001000011;
      patterns[37401] = 29'b1_001001000011_001_1_000011001001;
      patterns[37402] = 29'b1_001001000011_010_0_010010000111;
      patterns[37403] = 29'b1_001001000011_011_0_100100001110;
      patterns[37404] = 29'b1_001001000011_100_1_100100100001;
      patterns[37405] = 29'b1_001001000011_101_1_110010010000;
      patterns[37406] = 29'b1_001001000011_110_1_001001000011;
      patterns[37407] = 29'b1_001001000011_111_1_001001000011;
      patterns[37408] = 29'b1_001001000100_000_1_001001000100;
      patterns[37409] = 29'b1_001001000100_001_1_000100001001;
      patterns[37410] = 29'b1_001001000100_010_0_010010001001;
      patterns[37411] = 29'b1_001001000100_011_0_100100010010;
      patterns[37412] = 29'b1_001001000100_100_0_100100100010;
      patterns[37413] = 29'b1_001001000100_101_0_010010010001;
      patterns[37414] = 29'b1_001001000100_110_1_001001000100;
      patterns[37415] = 29'b1_001001000100_111_1_001001000100;
      patterns[37416] = 29'b1_001001000101_000_1_001001000101;
      patterns[37417] = 29'b1_001001000101_001_1_000101001001;
      patterns[37418] = 29'b1_001001000101_010_0_010010001011;
      patterns[37419] = 29'b1_001001000101_011_0_100100010110;
      patterns[37420] = 29'b1_001001000101_100_1_100100100010;
      patterns[37421] = 29'b1_001001000101_101_0_110010010001;
      patterns[37422] = 29'b1_001001000101_110_1_001001000101;
      patterns[37423] = 29'b1_001001000101_111_1_001001000101;
      patterns[37424] = 29'b1_001001000110_000_1_001001000110;
      patterns[37425] = 29'b1_001001000110_001_1_000110001001;
      patterns[37426] = 29'b1_001001000110_010_0_010010001101;
      patterns[37427] = 29'b1_001001000110_011_0_100100011010;
      patterns[37428] = 29'b1_001001000110_100_0_100100100011;
      patterns[37429] = 29'b1_001001000110_101_1_010010010001;
      patterns[37430] = 29'b1_001001000110_110_1_001001000110;
      patterns[37431] = 29'b1_001001000110_111_1_001001000110;
      patterns[37432] = 29'b1_001001000111_000_1_001001000111;
      patterns[37433] = 29'b1_001001000111_001_1_000111001001;
      patterns[37434] = 29'b1_001001000111_010_0_010010001111;
      patterns[37435] = 29'b1_001001000111_011_0_100100011110;
      patterns[37436] = 29'b1_001001000111_100_1_100100100011;
      patterns[37437] = 29'b1_001001000111_101_1_110010010001;
      patterns[37438] = 29'b1_001001000111_110_1_001001000111;
      patterns[37439] = 29'b1_001001000111_111_1_001001000111;
      patterns[37440] = 29'b1_001001001000_000_1_001001001000;
      patterns[37441] = 29'b1_001001001000_001_1_001000001001;
      patterns[37442] = 29'b1_001001001000_010_0_010010010001;
      patterns[37443] = 29'b1_001001001000_011_0_100100100010;
      patterns[37444] = 29'b1_001001001000_100_0_100100100100;
      patterns[37445] = 29'b1_001001001000_101_0_010010010010;
      patterns[37446] = 29'b1_001001001000_110_1_001001001000;
      patterns[37447] = 29'b1_001001001000_111_1_001001001000;
      patterns[37448] = 29'b1_001001001001_000_1_001001001001;
      patterns[37449] = 29'b1_001001001001_001_1_001001001001;
      patterns[37450] = 29'b1_001001001001_010_0_010010010011;
      patterns[37451] = 29'b1_001001001001_011_0_100100100110;
      patterns[37452] = 29'b1_001001001001_100_1_100100100100;
      patterns[37453] = 29'b1_001001001001_101_0_110010010010;
      patterns[37454] = 29'b1_001001001001_110_1_001001001001;
      patterns[37455] = 29'b1_001001001001_111_1_001001001001;
      patterns[37456] = 29'b1_001001001010_000_1_001001001010;
      patterns[37457] = 29'b1_001001001010_001_1_001010001001;
      patterns[37458] = 29'b1_001001001010_010_0_010010010101;
      patterns[37459] = 29'b1_001001001010_011_0_100100101010;
      patterns[37460] = 29'b1_001001001010_100_0_100100100101;
      patterns[37461] = 29'b1_001001001010_101_1_010010010010;
      patterns[37462] = 29'b1_001001001010_110_1_001001001010;
      patterns[37463] = 29'b1_001001001010_111_1_001001001010;
      patterns[37464] = 29'b1_001001001011_000_1_001001001011;
      patterns[37465] = 29'b1_001001001011_001_1_001011001001;
      patterns[37466] = 29'b1_001001001011_010_0_010010010111;
      patterns[37467] = 29'b1_001001001011_011_0_100100101110;
      patterns[37468] = 29'b1_001001001011_100_1_100100100101;
      patterns[37469] = 29'b1_001001001011_101_1_110010010010;
      patterns[37470] = 29'b1_001001001011_110_1_001001001011;
      patterns[37471] = 29'b1_001001001011_111_1_001001001011;
      patterns[37472] = 29'b1_001001001100_000_1_001001001100;
      patterns[37473] = 29'b1_001001001100_001_1_001100001001;
      patterns[37474] = 29'b1_001001001100_010_0_010010011001;
      patterns[37475] = 29'b1_001001001100_011_0_100100110010;
      patterns[37476] = 29'b1_001001001100_100_0_100100100110;
      patterns[37477] = 29'b1_001001001100_101_0_010010010011;
      patterns[37478] = 29'b1_001001001100_110_1_001001001100;
      patterns[37479] = 29'b1_001001001100_111_1_001001001100;
      patterns[37480] = 29'b1_001001001101_000_1_001001001101;
      patterns[37481] = 29'b1_001001001101_001_1_001101001001;
      patterns[37482] = 29'b1_001001001101_010_0_010010011011;
      patterns[37483] = 29'b1_001001001101_011_0_100100110110;
      patterns[37484] = 29'b1_001001001101_100_1_100100100110;
      patterns[37485] = 29'b1_001001001101_101_0_110010010011;
      patterns[37486] = 29'b1_001001001101_110_1_001001001101;
      patterns[37487] = 29'b1_001001001101_111_1_001001001101;
      patterns[37488] = 29'b1_001001001110_000_1_001001001110;
      patterns[37489] = 29'b1_001001001110_001_1_001110001001;
      patterns[37490] = 29'b1_001001001110_010_0_010010011101;
      patterns[37491] = 29'b1_001001001110_011_0_100100111010;
      patterns[37492] = 29'b1_001001001110_100_0_100100100111;
      patterns[37493] = 29'b1_001001001110_101_1_010010010011;
      patterns[37494] = 29'b1_001001001110_110_1_001001001110;
      patterns[37495] = 29'b1_001001001110_111_1_001001001110;
      patterns[37496] = 29'b1_001001001111_000_1_001001001111;
      patterns[37497] = 29'b1_001001001111_001_1_001111001001;
      patterns[37498] = 29'b1_001001001111_010_0_010010011111;
      patterns[37499] = 29'b1_001001001111_011_0_100100111110;
      patterns[37500] = 29'b1_001001001111_100_1_100100100111;
      patterns[37501] = 29'b1_001001001111_101_1_110010010011;
      patterns[37502] = 29'b1_001001001111_110_1_001001001111;
      patterns[37503] = 29'b1_001001001111_111_1_001001001111;
      patterns[37504] = 29'b1_001001010000_000_1_001001010000;
      patterns[37505] = 29'b1_001001010000_001_1_010000001001;
      patterns[37506] = 29'b1_001001010000_010_0_010010100001;
      patterns[37507] = 29'b1_001001010000_011_0_100101000010;
      patterns[37508] = 29'b1_001001010000_100_0_100100101000;
      patterns[37509] = 29'b1_001001010000_101_0_010010010100;
      patterns[37510] = 29'b1_001001010000_110_1_001001010000;
      patterns[37511] = 29'b1_001001010000_111_1_001001010000;
      patterns[37512] = 29'b1_001001010001_000_1_001001010001;
      patterns[37513] = 29'b1_001001010001_001_1_010001001001;
      patterns[37514] = 29'b1_001001010001_010_0_010010100011;
      patterns[37515] = 29'b1_001001010001_011_0_100101000110;
      patterns[37516] = 29'b1_001001010001_100_1_100100101000;
      patterns[37517] = 29'b1_001001010001_101_0_110010010100;
      patterns[37518] = 29'b1_001001010001_110_1_001001010001;
      patterns[37519] = 29'b1_001001010001_111_1_001001010001;
      patterns[37520] = 29'b1_001001010010_000_1_001001010010;
      patterns[37521] = 29'b1_001001010010_001_1_010010001001;
      patterns[37522] = 29'b1_001001010010_010_0_010010100101;
      patterns[37523] = 29'b1_001001010010_011_0_100101001010;
      patterns[37524] = 29'b1_001001010010_100_0_100100101001;
      patterns[37525] = 29'b1_001001010010_101_1_010010010100;
      patterns[37526] = 29'b1_001001010010_110_1_001001010010;
      patterns[37527] = 29'b1_001001010010_111_1_001001010010;
      patterns[37528] = 29'b1_001001010011_000_1_001001010011;
      patterns[37529] = 29'b1_001001010011_001_1_010011001001;
      patterns[37530] = 29'b1_001001010011_010_0_010010100111;
      patterns[37531] = 29'b1_001001010011_011_0_100101001110;
      patterns[37532] = 29'b1_001001010011_100_1_100100101001;
      patterns[37533] = 29'b1_001001010011_101_1_110010010100;
      patterns[37534] = 29'b1_001001010011_110_1_001001010011;
      patterns[37535] = 29'b1_001001010011_111_1_001001010011;
      patterns[37536] = 29'b1_001001010100_000_1_001001010100;
      patterns[37537] = 29'b1_001001010100_001_1_010100001001;
      patterns[37538] = 29'b1_001001010100_010_0_010010101001;
      patterns[37539] = 29'b1_001001010100_011_0_100101010010;
      patterns[37540] = 29'b1_001001010100_100_0_100100101010;
      patterns[37541] = 29'b1_001001010100_101_0_010010010101;
      patterns[37542] = 29'b1_001001010100_110_1_001001010100;
      patterns[37543] = 29'b1_001001010100_111_1_001001010100;
      patterns[37544] = 29'b1_001001010101_000_1_001001010101;
      patterns[37545] = 29'b1_001001010101_001_1_010101001001;
      patterns[37546] = 29'b1_001001010101_010_0_010010101011;
      patterns[37547] = 29'b1_001001010101_011_0_100101010110;
      patterns[37548] = 29'b1_001001010101_100_1_100100101010;
      patterns[37549] = 29'b1_001001010101_101_0_110010010101;
      patterns[37550] = 29'b1_001001010101_110_1_001001010101;
      patterns[37551] = 29'b1_001001010101_111_1_001001010101;
      patterns[37552] = 29'b1_001001010110_000_1_001001010110;
      patterns[37553] = 29'b1_001001010110_001_1_010110001001;
      patterns[37554] = 29'b1_001001010110_010_0_010010101101;
      patterns[37555] = 29'b1_001001010110_011_0_100101011010;
      patterns[37556] = 29'b1_001001010110_100_0_100100101011;
      patterns[37557] = 29'b1_001001010110_101_1_010010010101;
      patterns[37558] = 29'b1_001001010110_110_1_001001010110;
      patterns[37559] = 29'b1_001001010110_111_1_001001010110;
      patterns[37560] = 29'b1_001001010111_000_1_001001010111;
      patterns[37561] = 29'b1_001001010111_001_1_010111001001;
      patterns[37562] = 29'b1_001001010111_010_0_010010101111;
      patterns[37563] = 29'b1_001001010111_011_0_100101011110;
      patterns[37564] = 29'b1_001001010111_100_1_100100101011;
      patterns[37565] = 29'b1_001001010111_101_1_110010010101;
      patterns[37566] = 29'b1_001001010111_110_1_001001010111;
      patterns[37567] = 29'b1_001001010111_111_1_001001010111;
      patterns[37568] = 29'b1_001001011000_000_1_001001011000;
      patterns[37569] = 29'b1_001001011000_001_1_011000001001;
      patterns[37570] = 29'b1_001001011000_010_0_010010110001;
      patterns[37571] = 29'b1_001001011000_011_0_100101100010;
      patterns[37572] = 29'b1_001001011000_100_0_100100101100;
      patterns[37573] = 29'b1_001001011000_101_0_010010010110;
      patterns[37574] = 29'b1_001001011000_110_1_001001011000;
      patterns[37575] = 29'b1_001001011000_111_1_001001011000;
      patterns[37576] = 29'b1_001001011001_000_1_001001011001;
      patterns[37577] = 29'b1_001001011001_001_1_011001001001;
      patterns[37578] = 29'b1_001001011001_010_0_010010110011;
      patterns[37579] = 29'b1_001001011001_011_0_100101100110;
      patterns[37580] = 29'b1_001001011001_100_1_100100101100;
      patterns[37581] = 29'b1_001001011001_101_0_110010010110;
      patterns[37582] = 29'b1_001001011001_110_1_001001011001;
      patterns[37583] = 29'b1_001001011001_111_1_001001011001;
      patterns[37584] = 29'b1_001001011010_000_1_001001011010;
      patterns[37585] = 29'b1_001001011010_001_1_011010001001;
      patterns[37586] = 29'b1_001001011010_010_0_010010110101;
      patterns[37587] = 29'b1_001001011010_011_0_100101101010;
      patterns[37588] = 29'b1_001001011010_100_0_100100101101;
      patterns[37589] = 29'b1_001001011010_101_1_010010010110;
      patterns[37590] = 29'b1_001001011010_110_1_001001011010;
      patterns[37591] = 29'b1_001001011010_111_1_001001011010;
      patterns[37592] = 29'b1_001001011011_000_1_001001011011;
      patterns[37593] = 29'b1_001001011011_001_1_011011001001;
      patterns[37594] = 29'b1_001001011011_010_0_010010110111;
      patterns[37595] = 29'b1_001001011011_011_0_100101101110;
      patterns[37596] = 29'b1_001001011011_100_1_100100101101;
      patterns[37597] = 29'b1_001001011011_101_1_110010010110;
      patterns[37598] = 29'b1_001001011011_110_1_001001011011;
      patterns[37599] = 29'b1_001001011011_111_1_001001011011;
      patterns[37600] = 29'b1_001001011100_000_1_001001011100;
      patterns[37601] = 29'b1_001001011100_001_1_011100001001;
      patterns[37602] = 29'b1_001001011100_010_0_010010111001;
      patterns[37603] = 29'b1_001001011100_011_0_100101110010;
      patterns[37604] = 29'b1_001001011100_100_0_100100101110;
      patterns[37605] = 29'b1_001001011100_101_0_010010010111;
      patterns[37606] = 29'b1_001001011100_110_1_001001011100;
      patterns[37607] = 29'b1_001001011100_111_1_001001011100;
      patterns[37608] = 29'b1_001001011101_000_1_001001011101;
      patterns[37609] = 29'b1_001001011101_001_1_011101001001;
      patterns[37610] = 29'b1_001001011101_010_0_010010111011;
      patterns[37611] = 29'b1_001001011101_011_0_100101110110;
      patterns[37612] = 29'b1_001001011101_100_1_100100101110;
      patterns[37613] = 29'b1_001001011101_101_0_110010010111;
      patterns[37614] = 29'b1_001001011101_110_1_001001011101;
      patterns[37615] = 29'b1_001001011101_111_1_001001011101;
      patterns[37616] = 29'b1_001001011110_000_1_001001011110;
      patterns[37617] = 29'b1_001001011110_001_1_011110001001;
      patterns[37618] = 29'b1_001001011110_010_0_010010111101;
      patterns[37619] = 29'b1_001001011110_011_0_100101111010;
      patterns[37620] = 29'b1_001001011110_100_0_100100101111;
      patterns[37621] = 29'b1_001001011110_101_1_010010010111;
      patterns[37622] = 29'b1_001001011110_110_1_001001011110;
      patterns[37623] = 29'b1_001001011110_111_1_001001011110;
      patterns[37624] = 29'b1_001001011111_000_1_001001011111;
      patterns[37625] = 29'b1_001001011111_001_1_011111001001;
      patterns[37626] = 29'b1_001001011111_010_0_010010111111;
      patterns[37627] = 29'b1_001001011111_011_0_100101111110;
      patterns[37628] = 29'b1_001001011111_100_1_100100101111;
      patterns[37629] = 29'b1_001001011111_101_1_110010010111;
      patterns[37630] = 29'b1_001001011111_110_1_001001011111;
      patterns[37631] = 29'b1_001001011111_111_1_001001011111;
      patterns[37632] = 29'b1_001001100000_000_1_001001100000;
      patterns[37633] = 29'b1_001001100000_001_1_100000001001;
      patterns[37634] = 29'b1_001001100000_010_0_010011000001;
      patterns[37635] = 29'b1_001001100000_011_0_100110000010;
      patterns[37636] = 29'b1_001001100000_100_0_100100110000;
      patterns[37637] = 29'b1_001001100000_101_0_010010011000;
      patterns[37638] = 29'b1_001001100000_110_1_001001100000;
      patterns[37639] = 29'b1_001001100000_111_1_001001100000;
      patterns[37640] = 29'b1_001001100001_000_1_001001100001;
      patterns[37641] = 29'b1_001001100001_001_1_100001001001;
      patterns[37642] = 29'b1_001001100001_010_0_010011000011;
      patterns[37643] = 29'b1_001001100001_011_0_100110000110;
      patterns[37644] = 29'b1_001001100001_100_1_100100110000;
      patterns[37645] = 29'b1_001001100001_101_0_110010011000;
      patterns[37646] = 29'b1_001001100001_110_1_001001100001;
      patterns[37647] = 29'b1_001001100001_111_1_001001100001;
      patterns[37648] = 29'b1_001001100010_000_1_001001100010;
      patterns[37649] = 29'b1_001001100010_001_1_100010001001;
      patterns[37650] = 29'b1_001001100010_010_0_010011000101;
      patterns[37651] = 29'b1_001001100010_011_0_100110001010;
      patterns[37652] = 29'b1_001001100010_100_0_100100110001;
      patterns[37653] = 29'b1_001001100010_101_1_010010011000;
      patterns[37654] = 29'b1_001001100010_110_1_001001100010;
      patterns[37655] = 29'b1_001001100010_111_1_001001100010;
      patterns[37656] = 29'b1_001001100011_000_1_001001100011;
      patterns[37657] = 29'b1_001001100011_001_1_100011001001;
      patterns[37658] = 29'b1_001001100011_010_0_010011000111;
      patterns[37659] = 29'b1_001001100011_011_0_100110001110;
      patterns[37660] = 29'b1_001001100011_100_1_100100110001;
      patterns[37661] = 29'b1_001001100011_101_1_110010011000;
      patterns[37662] = 29'b1_001001100011_110_1_001001100011;
      patterns[37663] = 29'b1_001001100011_111_1_001001100011;
      patterns[37664] = 29'b1_001001100100_000_1_001001100100;
      patterns[37665] = 29'b1_001001100100_001_1_100100001001;
      patterns[37666] = 29'b1_001001100100_010_0_010011001001;
      patterns[37667] = 29'b1_001001100100_011_0_100110010010;
      patterns[37668] = 29'b1_001001100100_100_0_100100110010;
      patterns[37669] = 29'b1_001001100100_101_0_010010011001;
      patterns[37670] = 29'b1_001001100100_110_1_001001100100;
      patterns[37671] = 29'b1_001001100100_111_1_001001100100;
      patterns[37672] = 29'b1_001001100101_000_1_001001100101;
      patterns[37673] = 29'b1_001001100101_001_1_100101001001;
      patterns[37674] = 29'b1_001001100101_010_0_010011001011;
      patterns[37675] = 29'b1_001001100101_011_0_100110010110;
      patterns[37676] = 29'b1_001001100101_100_1_100100110010;
      patterns[37677] = 29'b1_001001100101_101_0_110010011001;
      patterns[37678] = 29'b1_001001100101_110_1_001001100101;
      patterns[37679] = 29'b1_001001100101_111_1_001001100101;
      patterns[37680] = 29'b1_001001100110_000_1_001001100110;
      patterns[37681] = 29'b1_001001100110_001_1_100110001001;
      patterns[37682] = 29'b1_001001100110_010_0_010011001101;
      patterns[37683] = 29'b1_001001100110_011_0_100110011010;
      patterns[37684] = 29'b1_001001100110_100_0_100100110011;
      patterns[37685] = 29'b1_001001100110_101_1_010010011001;
      patterns[37686] = 29'b1_001001100110_110_1_001001100110;
      patterns[37687] = 29'b1_001001100110_111_1_001001100110;
      patterns[37688] = 29'b1_001001100111_000_1_001001100111;
      patterns[37689] = 29'b1_001001100111_001_1_100111001001;
      patterns[37690] = 29'b1_001001100111_010_0_010011001111;
      patterns[37691] = 29'b1_001001100111_011_0_100110011110;
      patterns[37692] = 29'b1_001001100111_100_1_100100110011;
      patterns[37693] = 29'b1_001001100111_101_1_110010011001;
      patterns[37694] = 29'b1_001001100111_110_1_001001100111;
      patterns[37695] = 29'b1_001001100111_111_1_001001100111;
      patterns[37696] = 29'b1_001001101000_000_1_001001101000;
      patterns[37697] = 29'b1_001001101000_001_1_101000001001;
      patterns[37698] = 29'b1_001001101000_010_0_010011010001;
      patterns[37699] = 29'b1_001001101000_011_0_100110100010;
      patterns[37700] = 29'b1_001001101000_100_0_100100110100;
      patterns[37701] = 29'b1_001001101000_101_0_010010011010;
      patterns[37702] = 29'b1_001001101000_110_1_001001101000;
      patterns[37703] = 29'b1_001001101000_111_1_001001101000;
      patterns[37704] = 29'b1_001001101001_000_1_001001101001;
      patterns[37705] = 29'b1_001001101001_001_1_101001001001;
      patterns[37706] = 29'b1_001001101001_010_0_010011010011;
      patterns[37707] = 29'b1_001001101001_011_0_100110100110;
      patterns[37708] = 29'b1_001001101001_100_1_100100110100;
      patterns[37709] = 29'b1_001001101001_101_0_110010011010;
      patterns[37710] = 29'b1_001001101001_110_1_001001101001;
      patterns[37711] = 29'b1_001001101001_111_1_001001101001;
      patterns[37712] = 29'b1_001001101010_000_1_001001101010;
      patterns[37713] = 29'b1_001001101010_001_1_101010001001;
      patterns[37714] = 29'b1_001001101010_010_0_010011010101;
      patterns[37715] = 29'b1_001001101010_011_0_100110101010;
      patterns[37716] = 29'b1_001001101010_100_0_100100110101;
      patterns[37717] = 29'b1_001001101010_101_1_010010011010;
      patterns[37718] = 29'b1_001001101010_110_1_001001101010;
      patterns[37719] = 29'b1_001001101010_111_1_001001101010;
      patterns[37720] = 29'b1_001001101011_000_1_001001101011;
      patterns[37721] = 29'b1_001001101011_001_1_101011001001;
      patterns[37722] = 29'b1_001001101011_010_0_010011010111;
      patterns[37723] = 29'b1_001001101011_011_0_100110101110;
      patterns[37724] = 29'b1_001001101011_100_1_100100110101;
      patterns[37725] = 29'b1_001001101011_101_1_110010011010;
      patterns[37726] = 29'b1_001001101011_110_1_001001101011;
      patterns[37727] = 29'b1_001001101011_111_1_001001101011;
      patterns[37728] = 29'b1_001001101100_000_1_001001101100;
      patterns[37729] = 29'b1_001001101100_001_1_101100001001;
      patterns[37730] = 29'b1_001001101100_010_0_010011011001;
      patterns[37731] = 29'b1_001001101100_011_0_100110110010;
      patterns[37732] = 29'b1_001001101100_100_0_100100110110;
      patterns[37733] = 29'b1_001001101100_101_0_010010011011;
      patterns[37734] = 29'b1_001001101100_110_1_001001101100;
      patterns[37735] = 29'b1_001001101100_111_1_001001101100;
      patterns[37736] = 29'b1_001001101101_000_1_001001101101;
      patterns[37737] = 29'b1_001001101101_001_1_101101001001;
      patterns[37738] = 29'b1_001001101101_010_0_010011011011;
      patterns[37739] = 29'b1_001001101101_011_0_100110110110;
      patterns[37740] = 29'b1_001001101101_100_1_100100110110;
      patterns[37741] = 29'b1_001001101101_101_0_110010011011;
      patterns[37742] = 29'b1_001001101101_110_1_001001101101;
      patterns[37743] = 29'b1_001001101101_111_1_001001101101;
      patterns[37744] = 29'b1_001001101110_000_1_001001101110;
      patterns[37745] = 29'b1_001001101110_001_1_101110001001;
      patterns[37746] = 29'b1_001001101110_010_0_010011011101;
      patterns[37747] = 29'b1_001001101110_011_0_100110111010;
      patterns[37748] = 29'b1_001001101110_100_0_100100110111;
      patterns[37749] = 29'b1_001001101110_101_1_010010011011;
      patterns[37750] = 29'b1_001001101110_110_1_001001101110;
      patterns[37751] = 29'b1_001001101110_111_1_001001101110;
      patterns[37752] = 29'b1_001001101111_000_1_001001101111;
      patterns[37753] = 29'b1_001001101111_001_1_101111001001;
      patterns[37754] = 29'b1_001001101111_010_0_010011011111;
      patterns[37755] = 29'b1_001001101111_011_0_100110111110;
      patterns[37756] = 29'b1_001001101111_100_1_100100110111;
      patterns[37757] = 29'b1_001001101111_101_1_110010011011;
      patterns[37758] = 29'b1_001001101111_110_1_001001101111;
      patterns[37759] = 29'b1_001001101111_111_1_001001101111;
      patterns[37760] = 29'b1_001001110000_000_1_001001110000;
      patterns[37761] = 29'b1_001001110000_001_1_110000001001;
      patterns[37762] = 29'b1_001001110000_010_0_010011100001;
      patterns[37763] = 29'b1_001001110000_011_0_100111000010;
      patterns[37764] = 29'b1_001001110000_100_0_100100111000;
      patterns[37765] = 29'b1_001001110000_101_0_010010011100;
      patterns[37766] = 29'b1_001001110000_110_1_001001110000;
      patterns[37767] = 29'b1_001001110000_111_1_001001110000;
      patterns[37768] = 29'b1_001001110001_000_1_001001110001;
      patterns[37769] = 29'b1_001001110001_001_1_110001001001;
      patterns[37770] = 29'b1_001001110001_010_0_010011100011;
      patterns[37771] = 29'b1_001001110001_011_0_100111000110;
      patterns[37772] = 29'b1_001001110001_100_1_100100111000;
      patterns[37773] = 29'b1_001001110001_101_0_110010011100;
      patterns[37774] = 29'b1_001001110001_110_1_001001110001;
      patterns[37775] = 29'b1_001001110001_111_1_001001110001;
      patterns[37776] = 29'b1_001001110010_000_1_001001110010;
      patterns[37777] = 29'b1_001001110010_001_1_110010001001;
      patterns[37778] = 29'b1_001001110010_010_0_010011100101;
      patterns[37779] = 29'b1_001001110010_011_0_100111001010;
      patterns[37780] = 29'b1_001001110010_100_0_100100111001;
      patterns[37781] = 29'b1_001001110010_101_1_010010011100;
      patterns[37782] = 29'b1_001001110010_110_1_001001110010;
      patterns[37783] = 29'b1_001001110010_111_1_001001110010;
      patterns[37784] = 29'b1_001001110011_000_1_001001110011;
      patterns[37785] = 29'b1_001001110011_001_1_110011001001;
      patterns[37786] = 29'b1_001001110011_010_0_010011100111;
      patterns[37787] = 29'b1_001001110011_011_0_100111001110;
      patterns[37788] = 29'b1_001001110011_100_1_100100111001;
      patterns[37789] = 29'b1_001001110011_101_1_110010011100;
      patterns[37790] = 29'b1_001001110011_110_1_001001110011;
      patterns[37791] = 29'b1_001001110011_111_1_001001110011;
      patterns[37792] = 29'b1_001001110100_000_1_001001110100;
      patterns[37793] = 29'b1_001001110100_001_1_110100001001;
      patterns[37794] = 29'b1_001001110100_010_0_010011101001;
      patterns[37795] = 29'b1_001001110100_011_0_100111010010;
      patterns[37796] = 29'b1_001001110100_100_0_100100111010;
      patterns[37797] = 29'b1_001001110100_101_0_010010011101;
      patterns[37798] = 29'b1_001001110100_110_1_001001110100;
      patterns[37799] = 29'b1_001001110100_111_1_001001110100;
      patterns[37800] = 29'b1_001001110101_000_1_001001110101;
      patterns[37801] = 29'b1_001001110101_001_1_110101001001;
      patterns[37802] = 29'b1_001001110101_010_0_010011101011;
      patterns[37803] = 29'b1_001001110101_011_0_100111010110;
      patterns[37804] = 29'b1_001001110101_100_1_100100111010;
      patterns[37805] = 29'b1_001001110101_101_0_110010011101;
      patterns[37806] = 29'b1_001001110101_110_1_001001110101;
      patterns[37807] = 29'b1_001001110101_111_1_001001110101;
      patterns[37808] = 29'b1_001001110110_000_1_001001110110;
      patterns[37809] = 29'b1_001001110110_001_1_110110001001;
      patterns[37810] = 29'b1_001001110110_010_0_010011101101;
      patterns[37811] = 29'b1_001001110110_011_0_100111011010;
      patterns[37812] = 29'b1_001001110110_100_0_100100111011;
      patterns[37813] = 29'b1_001001110110_101_1_010010011101;
      patterns[37814] = 29'b1_001001110110_110_1_001001110110;
      patterns[37815] = 29'b1_001001110110_111_1_001001110110;
      patterns[37816] = 29'b1_001001110111_000_1_001001110111;
      patterns[37817] = 29'b1_001001110111_001_1_110111001001;
      patterns[37818] = 29'b1_001001110111_010_0_010011101111;
      patterns[37819] = 29'b1_001001110111_011_0_100111011110;
      patterns[37820] = 29'b1_001001110111_100_1_100100111011;
      patterns[37821] = 29'b1_001001110111_101_1_110010011101;
      patterns[37822] = 29'b1_001001110111_110_1_001001110111;
      patterns[37823] = 29'b1_001001110111_111_1_001001110111;
      patterns[37824] = 29'b1_001001111000_000_1_001001111000;
      patterns[37825] = 29'b1_001001111000_001_1_111000001001;
      patterns[37826] = 29'b1_001001111000_010_0_010011110001;
      patterns[37827] = 29'b1_001001111000_011_0_100111100010;
      patterns[37828] = 29'b1_001001111000_100_0_100100111100;
      patterns[37829] = 29'b1_001001111000_101_0_010010011110;
      patterns[37830] = 29'b1_001001111000_110_1_001001111000;
      patterns[37831] = 29'b1_001001111000_111_1_001001111000;
      patterns[37832] = 29'b1_001001111001_000_1_001001111001;
      patterns[37833] = 29'b1_001001111001_001_1_111001001001;
      patterns[37834] = 29'b1_001001111001_010_0_010011110011;
      patterns[37835] = 29'b1_001001111001_011_0_100111100110;
      patterns[37836] = 29'b1_001001111001_100_1_100100111100;
      patterns[37837] = 29'b1_001001111001_101_0_110010011110;
      patterns[37838] = 29'b1_001001111001_110_1_001001111001;
      patterns[37839] = 29'b1_001001111001_111_1_001001111001;
      patterns[37840] = 29'b1_001001111010_000_1_001001111010;
      patterns[37841] = 29'b1_001001111010_001_1_111010001001;
      patterns[37842] = 29'b1_001001111010_010_0_010011110101;
      patterns[37843] = 29'b1_001001111010_011_0_100111101010;
      patterns[37844] = 29'b1_001001111010_100_0_100100111101;
      patterns[37845] = 29'b1_001001111010_101_1_010010011110;
      patterns[37846] = 29'b1_001001111010_110_1_001001111010;
      patterns[37847] = 29'b1_001001111010_111_1_001001111010;
      patterns[37848] = 29'b1_001001111011_000_1_001001111011;
      patterns[37849] = 29'b1_001001111011_001_1_111011001001;
      patterns[37850] = 29'b1_001001111011_010_0_010011110111;
      patterns[37851] = 29'b1_001001111011_011_0_100111101110;
      patterns[37852] = 29'b1_001001111011_100_1_100100111101;
      patterns[37853] = 29'b1_001001111011_101_1_110010011110;
      patterns[37854] = 29'b1_001001111011_110_1_001001111011;
      patterns[37855] = 29'b1_001001111011_111_1_001001111011;
      patterns[37856] = 29'b1_001001111100_000_1_001001111100;
      patterns[37857] = 29'b1_001001111100_001_1_111100001001;
      patterns[37858] = 29'b1_001001111100_010_0_010011111001;
      patterns[37859] = 29'b1_001001111100_011_0_100111110010;
      patterns[37860] = 29'b1_001001111100_100_0_100100111110;
      patterns[37861] = 29'b1_001001111100_101_0_010010011111;
      patterns[37862] = 29'b1_001001111100_110_1_001001111100;
      patterns[37863] = 29'b1_001001111100_111_1_001001111100;
      patterns[37864] = 29'b1_001001111101_000_1_001001111101;
      patterns[37865] = 29'b1_001001111101_001_1_111101001001;
      patterns[37866] = 29'b1_001001111101_010_0_010011111011;
      patterns[37867] = 29'b1_001001111101_011_0_100111110110;
      patterns[37868] = 29'b1_001001111101_100_1_100100111110;
      patterns[37869] = 29'b1_001001111101_101_0_110010011111;
      patterns[37870] = 29'b1_001001111101_110_1_001001111101;
      patterns[37871] = 29'b1_001001111101_111_1_001001111101;
      patterns[37872] = 29'b1_001001111110_000_1_001001111110;
      patterns[37873] = 29'b1_001001111110_001_1_111110001001;
      patterns[37874] = 29'b1_001001111110_010_0_010011111101;
      patterns[37875] = 29'b1_001001111110_011_0_100111111010;
      patterns[37876] = 29'b1_001001111110_100_0_100100111111;
      patterns[37877] = 29'b1_001001111110_101_1_010010011111;
      patterns[37878] = 29'b1_001001111110_110_1_001001111110;
      patterns[37879] = 29'b1_001001111110_111_1_001001111110;
      patterns[37880] = 29'b1_001001111111_000_1_001001111111;
      patterns[37881] = 29'b1_001001111111_001_1_111111001001;
      patterns[37882] = 29'b1_001001111111_010_0_010011111111;
      patterns[37883] = 29'b1_001001111111_011_0_100111111110;
      patterns[37884] = 29'b1_001001111111_100_1_100100111111;
      patterns[37885] = 29'b1_001001111111_101_1_110010011111;
      patterns[37886] = 29'b1_001001111111_110_1_001001111111;
      patterns[37887] = 29'b1_001001111111_111_1_001001111111;
      patterns[37888] = 29'b1_001010000000_000_1_001010000000;
      patterns[37889] = 29'b1_001010000000_001_1_000000001010;
      patterns[37890] = 29'b1_001010000000_010_0_010100000001;
      patterns[37891] = 29'b1_001010000000_011_0_101000000010;
      patterns[37892] = 29'b1_001010000000_100_0_100101000000;
      patterns[37893] = 29'b1_001010000000_101_0_010010100000;
      patterns[37894] = 29'b1_001010000000_110_1_001010000000;
      patterns[37895] = 29'b1_001010000000_111_1_001010000000;
      patterns[37896] = 29'b1_001010000001_000_1_001010000001;
      patterns[37897] = 29'b1_001010000001_001_1_000001001010;
      patterns[37898] = 29'b1_001010000001_010_0_010100000011;
      patterns[37899] = 29'b1_001010000001_011_0_101000000110;
      patterns[37900] = 29'b1_001010000001_100_1_100101000000;
      patterns[37901] = 29'b1_001010000001_101_0_110010100000;
      patterns[37902] = 29'b1_001010000001_110_1_001010000001;
      patterns[37903] = 29'b1_001010000001_111_1_001010000001;
      patterns[37904] = 29'b1_001010000010_000_1_001010000010;
      patterns[37905] = 29'b1_001010000010_001_1_000010001010;
      patterns[37906] = 29'b1_001010000010_010_0_010100000101;
      patterns[37907] = 29'b1_001010000010_011_0_101000001010;
      patterns[37908] = 29'b1_001010000010_100_0_100101000001;
      patterns[37909] = 29'b1_001010000010_101_1_010010100000;
      patterns[37910] = 29'b1_001010000010_110_1_001010000010;
      patterns[37911] = 29'b1_001010000010_111_1_001010000010;
      patterns[37912] = 29'b1_001010000011_000_1_001010000011;
      patterns[37913] = 29'b1_001010000011_001_1_000011001010;
      patterns[37914] = 29'b1_001010000011_010_0_010100000111;
      patterns[37915] = 29'b1_001010000011_011_0_101000001110;
      patterns[37916] = 29'b1_001010000011_100_1_100101000001;
      patterns[37917] = 29'b1_001010000011_101_1_110010100000;
      patterns[37918] = 29'b1_001010000011_110_1_001010000011;
      patterns[37919] = 29'b1_001010000011_111_1_001010000011;
      patterns[37920] = 29'b1_001010000100_000_1_001010000100;
      patterns[37921] = 29'b1_001010000100_001_1_000100001010;
      patterns[37922] = 29'b1_001010000100_010_0_010100001001;
      patterns[37923] = 29'b1_001010000100_011_0_101000010010;
      patterns[37924] = 29'b1_001010000100_100_0_100101000010;
      patterns[37925] = 29'b1_001010000100_101_0_010010100001;
      patterns[37926] = 29'b1_001010000100_110_1_001010000100;
      patterns[37927] = 29'b1_001010000100_111_1_001010000100;
      patterns[37928] = 29'b1_001010000101_000_1_001010000101;
      patterns[37929] = 29'b1_001010000101_001_1_000101001010;
      patterns[37930] = 29'b1_001010000101_010_0_010100001011;
      patterns[37931] = 29'b1_001010000101_011_0_101000010110;
      patterns[37932] = 29'b1_001010000101_100_1_100101000010;
      patterns[37933] = 29'b1_001010000101_101_0_110010100001;
      patterns[37934] = 29'b1_001010000101_110_1_001010000101;
      patterns[37935] = 29'b1_001010000101_111_1_001010000101;
      patterns[37936] = 29'b1_001010000110_000_1_001010000110;
      patterns[37937] = 29'b1_001010000110_001_1_000110001010;
      patterns[37938] = 29'b1_001010000110_010_0_010100001101;
      patterns[37939] = 29'b1_001010000110_011_0_101000011010;
      patterns[37940] = 29'b1_001010000110_100_0_100101000011;
      patterns[37941] = 29'b1_001010000110_101_1_010010100001;
      patterns[37942] = 29'b1_001010000110_110_1_001010000110;
      patterns[37943] = 29'b1_001010000110_111_1_001010000110;
      patterns[37944] = 29'b1_001010000111_000_1_001010000111;
      patterns[37945] = 29'b1_001010000111_001_1_000111001010;
      patterns[37946] = 29'b1_001010000111_010_0_010100001111;
      patterns[37947] = 29'b1_001010000111_011_0_101000011110;
      patterns[37948] = 29'b1_001010000111_100_1_100101000011;
      patterns[37949] = 29'b1_001010000111_101_1_110010100001;
      patterns[37950] = 29'b1_001010000111_110_1_001010000111;
      patterns[37951] = 29'b1_001010000111_111_1_001010000111;
      patterns[37952] = 29'b1_001010001000_000_1_001010001000;
      patterns[37953] = 29'b1_001010001000_001_1_001000001010;
      patterns[37954] = 29'b1_001010001000_010_0_010100010001;
      patterns[37955] = 29'b1_001010001000_011_0_101000100010;
      patterns[37956] = 29'b1_001010001000_100_0_100101000100;
      patterns[37957] = 29'b1_001010001000_101_0_010010100010;
      patterns[37958] = 29'b1_001010001000_110_1_001010001000;
      patterns[37959] = 29'b1_001010001000_111_1_001010001000;
      patterns[37960] = 29'b1_001010001001_000_1_001010001001;
      patterns[37961] = 29'b1_001010001001_001_1_001001001010;
      patterns[37962] = 29'b1_001010001001_010_0_010100010011;
      patterns[37963] = 29'b1_001010001001_011_0_101000100110;
      patterns[37964] = 29'b1_001010001001_100_1_100101000100;
      patterns[37965] = 29'b1_001010001001_101_0_110010100010;
      patterns[37966] = 29'b1_001010001001_110_1_001010001001;
      patterns[37967] = 29'b1_001010001001_111_1_001010001001;
      patterns[37968] = 29'b1_001010001010_000_1_001010001010;
      patterns[37969] = 29'b1_001010001010_001_1_001010001010;
      patterns[37970] = 29'b1_001010001010_010_0_010100010101;
      patterns[37971] = 29'b1_001010001010_011_0_101000101010;
      patterns[37972] = 29'b1_001010001010_100_0_100101000101;
      patterns[37973] = 29'b1_001010001010_101_1_010010100010;
      patterns[37974] = 29'b1_001010001010_110_1_001010001010;
      patterns[37975] = 29'b1_001010001010_111_1_001010001010;
      patterns[37976] = 29'b1_001010001011_000_1_001010001011;
      patterns[37977] = 29'b1_001010001011_001_1_001011001010;
      patterns[37978] = 29'b1_001010001011_010_0_010100010111;
      patterns[37979] = 29'b1_001010001011_011_0_101000101110;
      patterns[37980] = 29'b1_001010001011_100_1_100101000101;
      patterns[37981] = 29'b1_001010001011_101_1_110010100010;
      patterns[37982] = 29'b1_001010001011_110_1_001010001011;
      patterns[37983] = 29'b1_001010001011_111_1_001010001011;
      patterns[37984] = 29'b1_001010001100_000_1_001010001100;
      patterns[37985] = 29'b1_001010001100_001_1_001100001010;
      patterns[37986] = 29'b1_001010001100_010_0_010100011001;
      patterns[37987] = 29'b1_001010001100_011_0_101000110010;
      patterns[37988] = 29'b1_001010001100_100_0_100101000110;
      patterns[37989] = 29'b1_001010001100_101_0_010010100011;
      patterns[37990] = 29'b1_001010001100_110_1_001010001100;
      patterns[37991] = 29'b1_001010001100_111_1_001010001100;
      patterns[37992] = 29'b1_001010001101_000_1_001010001101;
      patterns[37993] = 29'b1_001010001101_001_1_001101001010;
      patterns[37994] = 29'b1_001010001101_010_0_010100011011;
      patterns[37995] = 29'b1_001010001101_011_0_101000110110;
      patterns[37996] = 29'b1_001010001101_100_1_100101000110;
      patterns[37997] = 29'b1_001010001101_101_0_110010100011;
      patterns[37998] = 29'b1_001010001101_110_1_001010001101;
      patterns[37999] = 29'b1_001010001101_111_1_001010001101;
      patterns[38000] = 29'b1_001010001110_000_1_001010001110;
      patterns[38001] = 29'b1_001010001110_001_1_001110001010;
      patterns[38002] = 29'b1_001010001110_010_0_010100011101;
      patterns[38003] = 29'b1_001010001110_011_0_101000111010;
      patterns[38004] = 29'b1_001010001110_100_0_100101000111;
      patterns[38005] = 29'b1_001010001110_101_1_010010100011;
      patterns[38006] = 29'b1_001010001110_110_1_001010001110;
      patterns[38007] = 29'b1_001010001110_111_1_001010001110;
      patterns[38008] = 29'b1_001010001111_000_1_001010001111;
      patterns[38009] = 29'b1_001010001111_001_1_001111001010;
      patterns[38010] = 29'b1_001010001111_010_0_010100011111;
      patterns[38011] = 29'b1_001010001111_011_0_101000111110;
      patterns[38012] = 29'b1_001010001111_100_1_100101000111;
      patterns[38013] = 29'b1_001010001111_101_1_110010100011;
      patterns[38014] = 29'b1_001010001111_110_1_001010001111;
      patterns[38015] = 29'b1_001010001111_111_1_001010001111;
      patterns[38016] = 29'b1_001010010000_000_1_001010010000;
      patterns[38017] = 29'b1_001010010000_001_1_010000001010;
      patterns[38018] = 29'b1_001010010000_010_0_010100100001;
      patterns[38019] = 29'b1_001010010000_011_0_101001000010;
      patterns[38020] = 29'b1_001010010000_100_0_100101001000;
      patterns[38021] = 29'b1_001010010000_101_0_010010100100;
      patterns[38022] = 29'b1_001010010000_110_1_001010010000;
      patterns[38023] = 29'b1_001010010000_111_1_001010010000;
      patterns[38024] = 29'b1_001010010001_000_1_001010010001;
      patterns[38025] = 29'b1_001010010001_001_1_010001001010;
      patterns[38026] = 29'b1_001010010001_010_0_010100100011;
      patterns[38027] = 29'b1_001010010001_011_0_101001000110;
      patterns[38028] = 29'b1_001010010001_100_1_100101001000;
      patterns[38029] = 29'b1_001010010001_101_0_110010100100;
      patterns[38030] = 29'b1_001010010001_110_1_001010010001;
      patterns[38031] = 29'b1_001010010001_111_1_001010010001;
      patterns[38032] = 29'b1_001010010010_000_1_001010010010;
      patterns[38033] = 29'b1_001010010010_001_1_010010001010;
      patterns[38034] = 29'b1_001010010010_010_0_010100100101;
      patterns[38035] = 29'b1_001010010010_011_0_101001001010;
      patterns[38036] = 29'b1_001010010010_100_0_100101001001;
      patterns[38037] = 29'b1_001010010010_101_1_010010100100;
      patterns[38038] = 29'b1_001010010010_110_1_001010010010;
      patterns[38039] = 29'b1_001010010010_111_1_001010010010;
      patterns[38040] = 29'b1_001010010011_000_1_001010010011;
      patterns[38041] = 29'b1_001010010011_001_1_010011001010;
      patterns[38042] = 29'b1_001010010011_010_0_010100100111;
      patterns[38043] = 29'b1_001010010011_011_0_101001001110;
      patterns[38044] = 29'b1_001010010011_100_1_100101001001;
      patterns[38045] = 29'b1_001010010011_101_1_110010100100;
      patterns[38046] = 29'b1_001010010011_110_1_001010010011;
      patterns[38047] = 29'b1_001010010011_111_1_001010010011;
      patterns[38048] = 29'b1_001010010100_000_1_001010010100;
      patterns[38049] = 29'b1_001010010100_001_1_010100001010;
      patterns[38050] = 29'b1_001010010100_010_0_010100101001;
      patterns[38051] = 29'b1_001010010100_011_0_101001010010;
      patterns[38052] = 29'b1_001010010100_100_0_100101001010;
      patterns[38053] = 29'b1_001010010100_101_0_010010100101;
      patterns[38054] = 29'b1_001010010100_110_1_001010010100;
      patterns[38055] = 29'b1_001010010100_111_1_001010010100;
      patterns[38056] = 29'b1_001010010101_000_1_001010010101;
      patterns[38057] = 29'b1_001010010101_001_1_010101001010;
      patterns[38058] = 29'b1_001010010101_010_0_010100101011;
      patterns[38059] = 29'b1_001010010101_011_0_101001010110;
      patterns[38060] = 29'b1_001010010101_100_1_100101001010;
      patterns[38061] = 29'b1_001010010101_101_0_110010100101;
      patterns[38062] = 29'b1_001010010101_110_1_001010010101;
      patterns[38063] = 29'b1_001010010101_111_1_001010010101;
      patterns[38064] = 29'b1_001010010110_000_1_001010010110;
      patterns[38065] = 29'b1_001010010110_001_1_010110001010;
      patterns[38066] = 29'b1_001010010110_010_0_010100101101;
      patterns[38067] = 29'b1_001010010110_011_0_101001011010;
      patterns[38068] = 29'b1_001010010110_100_0_100101001011;
      patterns[38069] = 29'b1_001010010110_101_1_010010100101;
      patterns[38070] = 29'b1_001010010110_110_1_001010010110;
      patterns[38071] = 29'b1_001010010110_111_1_001010010110;
      patterns[38072] = 29'b1_001010010111_000_1_001010010111;
      patterns[38073] = 29'b1_001010010111_001_1_010111001010;
      patterns[38074] = 29'b1_001010010111_010_0_010100101111;
      patterns[38075] = 29'b1_001010010111_011_0_101001011110;
      patterns[38076] = 29'b1_001010010111_100_1_100101001011;
      patterns[38077] = 29'b1_001010010111_101_1_110010100101;
      patterns[38078] = 29'b1_001010010111_110_1_001010010111;
      patterns[38079] = 29'b1_001010010111_111_1_001010010111;
      patterns[38080] = 29'b1_001010011000_000_1_001010011000;
      patterns[38081] = 29'b1_001010011000_001_1_011000001010;
      patterns[38082] = 29'b1_001010011000_010_0_010100110001;
      patterns[38083] = 29'b1_001010011000_011_0_101001100010;
      patterns[38084] = 29'b1_001010011000_100_0_100101001100;
      patterns[38085] = 29'b1_001010011000_101_0_010010100110;
      patterns[38086] = 29'b1_001010011000_110_1_001010011000;
      patterns[38087] = 29'b1_001010011000_111_1_001010011000;
      patterns[38088] = 29'b1_001010011001_000_1_001010011001;
      patterns[38089] = 29'b1_001010011001_001_1_011001001010;
      patterns[38090] = 29'b1_001010011001_010_0_010100110011;
      patterns[38091] = 29'b1_001010011001_011_0_101001100110;
      patterns[38092] = 29'b1_001010011001_100_1_100101001100;
      patterns[38093] = 29'b1_001010011001_101_0_110010100110;
      patterns[38094] = 29'b1_001010011001_110_1_001010011001;
      patterns[38095] = 29'b1_001010011001_111_1_001010011001;
      patterns[38096] = 29'b1_001010011010_000_1_001010011010;
      patterns[38097] = 29'b1_001010011010_001_1_011010001010;
      patterns[38098] = 29'b1_001010011010_010_0_010100110101;
      patterns[38099] = 29'b1_001010011010_011_0_101001101010;
      patterns[38100] = 29'b1_001010011010_100_0_100101001101;
      patterns[38101] = 29'b1_001010011010_101_1_010010100110;
      patterns[38102] = 29'b1_001010011010_110_1_001010011010;
      patterns[38103] = 29'b1_001010011010_111_1_001010011010;
      patterns[38104] = 29'b1_001010011011_000_1_001010011011;
      patterns[38105] = 29'b1_001010011011_001_1_011011001010;
      patterns[38106] = 29'b1_001010011011_010_0_010100110111;
      patterns[38107] = 29'b1_001010011011_011_0_101001101110;
      patterns[38108] = 29'b1_001010011011_100_1_100101001101;
      patterns[38109] = 29'b1_001010011011_101_1_110010100110;
      patterns[38110] = 29'b1_001010011011_110_1_001010011011;
      patterns[38111] = 29'b1_001010011011_111_1_001010011011;
      patterns[38112] = 29'b1_001010011100_000_1_001010011100;
      patterns[38113] = 29'b1_001010011100_001_1_011100001010;
      patterns[38114] = 29'b1_001010011100_010_0_010100111001;
      patterns[38115] = 29'b1_001010011100_011_0_101001110010;
      patterns[38116] = 29'b1_001010011100_100_0_100101001110;
      patterns[38117] = 29'b1_001010011100_101_0_010010100111;
      patterns[38118] = 29'b1_001010011100_110_1_001010011100;
      patterns[38119] = 29'b1_001010011100_111_1_001010011100;
      patterns[38120] = 29'b1_001010011101_000_1_001010011101;
      patterns[38121] = 29'b1_001010011101_001_1_011101001010;
      patterns[38122] = 29'b1_001010011101_010_0_010100111011;
      patterns[38123] = 29'b1_001010011101_011_0_101001110110;
      patterns[38124] = 29'b1_001010011101_100_1_100101001110;
      patterns[38125] = 29'b1_001010011101_101_0_110010100111;
      patterns[38126] = 29'b1_001010011101_110_1_001010011101;
      patterns[38127] = 29'b1_001010011101_111_1_001010011101;
      patterns[38128] = 29'b1_001010011110_000_1_001010011110;
      patterns[38129] = 29'b1_001010011110_001_1_011110001010;
      patterns[38130] = 29'b1_001010011110_010_0_010100111101;
      patterns[38131] = 29'b1_001010011110_011_0_101001111010;
      patterns[38132] = 29'b1_001010011110_100_0_100101001111;
      patterns[38133] = 29'b1_001010011110_101_1_010010100111;
      patterns[38134] = 29'b1_001010011110_110_1_001010011110;
      patterns[38135] = 29'b1_001010011110_111_1_001010011110;
      patterns[38136] = 29'b1_001010011111_000_1_001010011111;
      patterns[38137] = 29'b1_001010011111_001_1_011111001010;
      patterns[38138] = 29'b1_001010011111_010_0_010100111111;
      patterns[38139] = 29'b1_001010011111_011_0_101001111110;
      patterns[38140] = 29'b1_001010011111_100_1_100101001111;
      patterns[38141] = 29'b1_001010011111_101_1_110010100111;
      patterns[38142] = 29'b1_001010011111_110_1_001010011111;
      patterns[38143] = 29'b1_001010011111_111_1_001010011111;
      patterns[38144] = 29'b1_001010100000_000_1_001010100000;
      patterns[38145] = 29'b1_001010100000_001_1_100000001010;
      patterns[38146] = 29'b1_001010100000_010_0_010101000001;
      patterns[38147] = 29'b1_001010100000_011_0_101010000010;
      patterns[38148] = 29'b1_001010100000_100_0_100101010000;
      patterns[38149] = 29'b1_001010100000_101_0_010010101000;
      patterns[38150] = 29'b1_001010100000_110_1_001010100000;
      patterns[38151] = 29'b1_001010100000_111_1_001010100000;
      patterns[38152] = 29'b1_001010100001_000_1_001010100001;
      patterns[38153] = 29'b1_001010100001_001_1_100001001010;
      patterns[38154] = 29'b1_001010100001_010_0_010101000011;
      patterns[38155] = 29'b1_001010100001_011_0_101010000110;
      patterns[38156] = 29'b1_001010100001_100_1_100101010000;
      patterns[38157] = 29'b1_001010100001_101_0_110010101000;
      patterns[38158] = 29'b1_001010100001_110_1_001010100001;
      patterns[38159] = 29'b1_001010100001_111_1_001010100001;
      patterns[38160] = 29'b1_001010100010_000_1_001010100010;
      patterns[38161] = 29'b1_001010100010_001_1_100010001010;
      patterns[38162] = 29'b1_001010100010_010_0_010101000101;
      patterns[38163] = 29'b1_001010100010_011_0_101010001010;
      patterns[38164] = 29'b1_001010100010_100_0_100101010001;
      patterns[38165] = 29'b1_001010100010_101_1_010010101000;
      patterns[38166] = 29'b1_001010100010_110_1_001010100010;
      patterns[38167] = 29'b1_001010100010_111_1_001010100010;
      patterns[38168] = 29'b1_001010100011_000_1_001010100011;
      patterns[38169] = 29'b1_001010100011_001_1_100011001010;
      patterns[38170] = 29'b1_001010100011_010_0_010101000111;
      patterns[38171] = 29'b1_001010100011_011_0_101010001110;
      patterns[38172] = 29'b1_001010100011_100_1_100101010001;
      patterns[38173] = 29'b1_001010100011_101_1_110010101000;
      patterns[38174] = 29'b1_001010100011_110_1_001010100011;
      patterns[38175] = 29'b1_001010100011_111_1_001010100011;
      patterns[38176] = 29'b1_001010100100_000_1_001010100100;
      patterns[38177] = 29'b1_001010100100_001_1_100100001010;
      patterns[38178] = 29'b1_001010100100_010_0_010101001001;
      patterns[38179] = 29'b1_001010100100_011_0_101010010010;
      patterns[38180] = 29'b1_001010100100_100_0_100101010010;
      patterns[38181] = 29'b1_001010100100_101_0_010010101001;
      patterns[38182] = 29'b1_001010100100_110_1_001010100100;
      patterns[38183] = 29'b1_001010100100_111_1_001010100100;
      patterns[38184] = 29'b1_001010100101_000_1_001010100101;
      patterns[38185] = 29'b1_001010100101_001_1_100101001010;
      patterns[38186] = 29'b1_001010100101_010_0_010101001011;
      patterns[38187] = 29'b1_001010100101_011_0_101010010110;
      patterns[38188] = 29'b1_001010100101_100_1_100101010010;
      patterns[38189] = 29'b1_001010100101_101_0_110010101001;
      patterns[38190] = 29'b1_001010100101_110_1_001010100101;
      patterns[38191] = 29'b1_001010100101_111_1_001010100101;
      patterns[38192] = 29'b1_001010100110_000_1_001010100110;
      patterns[38193] = 29'b1_001010100110_001_1_100110001010;
      patterns[38194] = 29'b1_001010100110_010_0_010101001101;
      patterns[38195] = 29'b1_001010100110_011_0_101010011010;
      patterns[38196] = 29'b1_001010100110_100_0_100101010011;
      patterns[38197] = 29'b1_001010100110_101_1_010010101001;
      patterns[38198] = 29'b1_001010100110_110_1_001010100110;
      patterns[38199] = 29'b1_001010100110_111_1_001010100110;
      patterns[38200] = 29'b1_001010100111_000_1_001010100111;
      patterns[38201] = 29'b1_001010100111_001_1_100111001010;
      patterns[38202] = 29'b1_001010100111_010_0_010101001111;
      patterns[38203] = 29'b1_001010100111_011_0_101010011110;
      patterns[38204] = 29'b1_001010100111_100_1_100101010011;
      patterns[38205] = 29'b1_001010100111_101_1_110010101001;
      patterns[38206] = 29'b1_001010100111_110_1_001010100111;
      patterns[38207] = 29'b1_001010100111_111_1_001010100111;
      patterns[38208] = 29'b1_001010101000_000_1_001010101000;
      patterns[38209] = 29'b1_001010101000_001_1_101000001010;
      patterns[38210] = 29'b1_001010101000_010_0_010101010001;
      patterns[38211] = 29'b1_001010101000_011_0_101010100010;
      patterns[38212] = 29'b1_001010101000_100_0_100101010100;
      patterns[38213] = 29'b1_001010101000_101_0_010010101010;
      patterns[38214] = 29'b1_001010101000_110_1_001010101000;
      patterns[38215] = 29'b1_001010101000_111_1_001010101000;
      patterns[38216] = 29'b1_001010101001_000_1_001010101001;
      patterns[38217] = 29'b1_001010101001_001_1_101001001010;
      patterns[38218] = 29'b1_001010101001_010_0_010101010011;
      patterns[38219] = 29'b1_001010101001_011_0_101010100110;
      patterns[38220] = 29'b1_001010101001_100_1_100101010100;
      patterns[38221] = 29'b1_001010101001_101_0_110010101010;
      patterns[38222] = 29'b1_001010101001_110_1_001010101001;
      patterns[38223] = 29'b1_001010101001_111_1_001010101001;
      patterns[38224] = 29'b1_001010101010_000_1_001010101010;
      patterns[38225] = 29'b1_001010101010_001_1_101010001010;
      patterns[38226] = 29'b1_001010101010_010_0_010101010101;
      patterns[38227] = 29'b1_001010101010_011_0_101010101010;
      patterns[38228] = 29'b1_001010101010_100_0_100101010101;
      patterns[38229] = 29'b1_001010101010_101_1_010010101010;
      patterns[38230] = 29'b1_001010101010_110_1_001010101010;
      patterns[38231] = 29'b1_001010101010_111_1_001010101010;
      patterns[38232] = 29'b1_001010101011_000_1_001010101011;
      patterns[38233] = 29'b1_001010101011_001_1_101011001010;
      patterns[38234] = 29'b1_001010101011_010_0_010101010111;
      patterns[38235] = 29'b1_001010101011_011_0_101010101110;
      patterns[38236] = 29'b1_001010101011_100_1_100101010101;
      patterns[38237] = 29'b1_001010101011_101_1_110010101010;
      patterns[38238] = 29'b1_001010101011_110_1_001010101011;
      patterns[38239] = 29'b1_001010101011_111_1_001010101011;
      patterns[38240] = 29'b1_001010101100_000_1_001010101100;
      patterns[38241] = 29'b1_001010101100_001_1_101100001010;
      patterns[38242] = 29'b1_001010101100_010_0_010101011001;
      patterns[38243] = 29'b1_001010101100_011_0_101010110010;
      patterns[38244] = 29'b1_001010101100_100_0_100101010110;
      patterns[38245] = 29'b1_001010101100_101_0_010010101011;
      patterns[38246] = 29'b1_001010101100_110_1_001010101100;
      patterns[38247] = 29'b1_001010101100_111_1_001010101100;
      patterns[38248] = 29'b1_001010101101_000_1_001010101101;
      patterns[38249] = 29'b1_001010101101_001_1_101101001010;
      patterns[38250] = 29'b1_001010101101_010_0_010101011011;
      patterns[38251] = 29'b1_001010101101_011_0_101010110110;
      patterns[38252] = 29'b1_001010101101_100_1_100101010110;
      patterns[38253] = 29'b1_001010101101_101_0_110010101011;
      patterns[38254] = 29'b1_001010101101_110_1_001010101101;
      patterns[38255] = 29'b1_001010101101_111_1_001010101101;
      patterns[38256] = 29'b1_001010101110_000_1_001010101110;
      patterns[38257] = 29'b1_001010101110_001_1_101110001010;
      patterns[38258] = 29'b1_001010101110_010_0_010101011101;
      patterns[38259] = 29'b1_001010101110_011_0_101010111010;
      patterns[38260] = 29'b1_001010101110_100_0_100101010111;
      patterns[38261] = 29'b1_001010101110_101_1_010010101011;
      patterns[38262] = 29'b1_001010101110_110_1_001010101110;
      patterns[38263] = 29'b1_001010101110_111_1_001010101110;
      patterns[38264] = 29'b1_001010101111_000_1_001010101111;
      patterns[38265] = 29'b1_001010101111_001_1_101111001010;
      patterns[38266] = 29'b1_001010101111_010_0_010101011111;
      patterns[38267] = 29'b1_001010101111_011_0_101010111110;
      patterns[38268] = 29'b1_001010101111_100_1_100101010111;
      patterns[38269] = 29'b1_001010101111_101_1_110010101011;
      patterns[38270] = 29'b1_001010101111_110_1_001010101111;
      patterns[38271] = 29'b1_001010101111_111_1_001010101111;
      patterns[38272] = 29'b1_001010110000_000_1_001010110000;
      patterns[38273] = 29'b1_001010110000_001_1_110000001010;
      patterns[38274] = 29'b1_001010110000_010_0_010101100001;
      patterns[38275] = 29'b1_001010110000_011_0_101011000010;
      patterns[38276] = 29'b1_001010110000_100_0_100101011000;
      patterns[38277] = 29'b1_001010110000_101_0_010010101100;
      patterns[38278] = 29'b1_001010110000_110_1_001010110000;
      patterns[38279] = 29'b1_001010110000_111_1_001010110000;
      patterns[38280] = 29'b1_001010110001_000_1_001010110001;
      patterns[38281] = 29'b1_001010110001_001_1_110001001010;
      patterns[38282] = 29'b1_001010110001_010_0_010101100011;
      patterns[38283] = 29'b1_001010110001_011_0_101011000110;
      patterns[38284] = 29'b1_001010110001_100_1_100101011000;
      patterns[38285] = 29'b1_001010110001_101_0_110010101100;
      patterns[38286] = 29'b1_001010110001_110_1_001010110001;
      patterns[38287] = 29'b1_001010110001_111_1_001010110001;
      patterns[38288] = 29'b1_001010110010_000_1_001010110010;
      patterns[38289] = 29'b1_001010110010_001_1_110010001010;
      patterns[38290] = 29'b1_001010110010_010_0_010101100101;
      patterns[38291] = 29'b1_001010110010_011_0_101011001010;
      patterns[38292] = 29'b1_001010110010_100_0_100101011001;
      patterns[38293] = 29'b1_001010110010_101_1_010010101100;
      patterns[38294] = 29'b1_001010110010_110_1_001010110010;
      patterns[38295] = 29'b1_001010110010_111_1_001010110010;
      patterns[38296] = 29'b1_001010110011_000_1_001010110011;
      patterns[38297] = 29'b1_001010110011_001_1_110011001010;
      patterns[38298] = 29'b1_001010110011_010_0_010101100111;
      patterns[38299] = 29'b1_001010110011_011_0_101011001110;
      patterns[38300] = 29'b1_001010110011_100_1_100101011001;
      patterns[38301] = 29'b1_001010110011_101_1_110010101100;
      patterns[38302] = 29'b1_001010110011_110_1_001010110011;
      patterns[38303] = 29'b1_001010110011_111_1_001010110011;
      patterns[38304] = 29'b1_001010110100_000_1_001010110100;
      patterns[38305] = 29'b1_001010110100_001_1_110100001010;
      patterns[38306] = 29'b1_001010110100_010_0_010101101001;
      patterns[38307] = 29'b1_001010110100_011_0_101011010010;
      patterns[38308] = 29'b1_001010110100_100_0_100101011010;
      patterns[38309] = 29'b1_001010110100_101_0_010010101101;
      patterns[38310] = 29'b1_001010110100_110_1_001010110100;
      patterns[38311] = 29'b1_001010110100_111_1_001010110100;
      patterns[38312] = 29'b1_001010110101_000_1_001010110101;
      patterns[38313] = 29'b1_001010110101_001_1_110101001010;
      patterns[38314] = 29'b1_001010110101_010_0_010101101011;
      patterns[38315] = 29'b1_001010110101_011_0_101011010110;
      patterns[38316] = 29'b1_001010110101_100_1_100101011010;
      patterns[38317] = 29'b1_001010110101_101_0_110010101101;
      patterns[38318] = 29'b1_001010110101_110_1_001010110101;
      patterns[38319] = 29'b1_001010110101_111_1_001010110101;
      patterns[38320] = 29'b1_001010110110_000_1_001010110110;
      patterns[38321] = 29'b1_001010110110_001_1_110110001010;
      patterns[38322] = 29'b1_001010110110_010_0_010101101101;
      patterns[38323] = 29'b1_001010110110_011_0_101011011010;
      patterns[38324] = 29'b1_001010110110_100_0_100101011011;
      patterns[38325] = 29'b1_001010110110_101_1_010010101101;
      patterns[38326] = 29'b1_001010110110_110_1_001010110110;
      patterns[38327] = 29'b1_001010110110_111_1_001010110110;
      patterns[38328] = 29'b1_001010110111_000_1_001010110111;
      patterns[38329] = 29'b1_001010110111_001_1_110111001010;
      patterns[38330] = 29'b1_001010110111_010_0_010101101111;
      patterns[38331] = 29'b1_001010110111_011_0_101011011110;
      patterns[38332] = 29'b1_001010110111_100_1_100101011011;
      patterns[38333] = 29'b1_001010110111_101_1_110010101101;
      patterns[38334] = 29'b1_001010110111_110_1_001010110111;
      patterns[38335] = 29'b1_001010110111_111_1_001010110111;
      patterns[38336] = 29'b1_001010111000_000_1_001010111000;
      patterns[38337] = 29'b1_001010111000_001_1_111000001010;
      patterns[38338] = 29'b1_001010111000_010_0_010101110001;
      patterns[38339] = 29'b1_001010111000_011_0_101011100010;
      patterns[38340] = 29'b1_001010111000_100_0_100101011100;
      patterns[38341] = 29'b1_001010111000_101_0_010010101110;
      patterns[38342] = 29'b1_001010111000_110_1_001010111000;
      patterns[38343] = 29'b1_001010111000_111_1_001010111000;
      patterns[38344] = 29'b1_001010111001_000_1_001010111001;
      patterns[38345] = 29'b1_001010111001_001_1_111001001010;
      patterns[38346] = 29'b1_001010111001_010_0_010101110011;
      patterns[38347] = 29'b1_001010111001_011_0_101011100110;
      patterns[38348] = 29'b1_001010111001_100_1_100101011100;
      patterns[38349] = 29'b1_001010111001_101_0_110010101110;
      patterns[38350] = 29'b1_001010111001_110_1_001010111001;
      patterns[38351] = 29'b1_001010111001_111_1_001010111001;
      patterns[38352] = 29'b1_001010111010_000_1_001010111010;
      patterns[38353] = 29'b1_001010111010_001_1_111010001010;
      patterns[38354] = 29'b1_001010111010_010_0_010101110101;
      patterns[38355] = 29'b1_001010111010_011_0_101011101010;
      patterns[38356] = 29'b1_001010111010_100_0_100101011101;
      patterns[38357] = 29'b1_001010111010_101_1_010010101110;
      patterns[38358] = 29'b1_001010111010_110_1_001010111010;
      patterns[38359] = 29'b1_001010111010_111_1_001010111010;
      patterns[38360] = 29'b1_001010111011_000_1_001010111011;
      patterns[38361] = 29'b1_001010111011_001_1_111011001010;
      patterns[38362] = 29'b1_001010111011_010_0_010101110111;
      patterns[38363] = 29'b1_001010111011_011_0_101011101110;
      patterns[38364] = 29'b1_001010111011_100_1_100101011101;
      patterns[38365] = 29'b1_001010111011_101_1_110010101110;
      patterns[38366] = 29'b1_001010111011_110_1_001010111011;
      patterns[38367] = 29'b1_001010111011_111_1_001010111011;
      patterns[38368] = 29'b1_001010111100_000_1_001010111100;
      patterns[38369] = 29'b1_001010111100_001_1_111100001010;
      patterns[38370] = 29'b1_001010111100_010_0_010101111001;
      patterns[38371] = 29'b1_001010111100_011_0_101011110010;
      patterns[38372] = 29'b1_001010111100_100_0_100101011110;
      patterns[38373] = 29'b1_001010111100_101_0_010010101111;
      patterns[38374] = 29'b1_001010111100_110_1_001010111100;
      patterns[38375] = 29'b1_001010111100_111_1_001010111100;
      patterns[38376] = 29'b1_001010111101_000_1_001010111101;
      patterns[38377] = 29'b1_001010111101_001_1_111101001010;
      patterns[38378] = 29'b1_001010111101_010_0_010101111011;
      patterns[38379] = 29'b1_001010111101_011_0_101011110110;
      patterns[38380] = 29'b1_001010111101_100_1_100101011110;
      patterns[38381] = 29'b1_001010111101_101_0_110010101111;
      patterns[38382] = 29'b1_001010111101_110_1_001010111101;
      patterns[38383] = 29'b1_001010111101_111_1_001010111101;
      patterns[38384] = 29'b1_001010111110_000_1_001010111110;
      patterns[38385] = 29'b1_001010111110_001_1_111110001010;
      patterns[38386] = 29'b1_001010111110_010_0_010101111101;
      patterns[38387] = 29'b1_001010111110_011_0_101011111010;
      patterns[38388] = 29'b1_001010111110_100_0_100101011111;
      patterns[38389] = 29'b1_001010111110_101_1_010010101111;
      patterns[38390] = 29'b1_001010111110_110_1_001010111110;
      patterns[38391] = 29'b1_001010111110_111_1_001010111110;
      patterns[38392] = 29'b1_001010111111_000_1_001010111111;
      patterns[38393] = 29'b1_001010111111_001_1_111111001010;
      patterns[38394] = 29'b1_001010111111_010_0_010101111111;
      patterns[38395] = 29'b1_001010111111_011_0_101011111110;
      patterns[38396] = 29'b1_001010111111_100_1_100101011111;
      patterns[38397] = 29'b1_001010111111_101_1_110010101111;
      patterns[38398] = 29'b1_001010111111_110_1_001010111111;
      patterns[38399] = 29'b1_001010111111_111_1_001010111111;
      patterns[38400] = 29'b1_001011000000_000_1_001011000000;
      patterns[38401] = 29'b1_001011000000_001_1_000000001011;
      patterns[38402] = 29'b1_001011000000_010_0_010110000001;
      patterns[38403] = 29'b1_001011000000_011_0_101100000010;
      patterns[38404] = 29'b1_001011000000_100_0_100101100000;
      patterns[38405] = 29'b1_001011000000_101_0_010010110000;
      patterns[38406] = 29'b1_001011000000_110_1_001011000000;
      patterns[38407] = 29'b1_001011000000_111_1_001011000000;
      patterns[38408] = 29'b1_001011000001_000_1_001011000001;
      patterns[38409] = 29'b1_001011000001_001_1_000001001011;
      patterns[38410] = 29'b1_001011000001_010_0_010110000011;
      patterns[38411] = 29'b1_001011000001_011_0_101100000110;
      patterns[38412] = 29'b1_001011000001_100_1_100101100000;
      patterns[38413] = 29'b1_001011000001_101_0_110010110000;
      patterns[38414] = 29'b1_001011000001_110_1_001011000001;
      patterns[38415] = 29'b1_001011000001_111_1_001011000001;
      patterns[38416] = 29'b1_001011000010_000_1_001011000010;
      patterns[38417] = 29'b1_001011000010_001_1_000010001011;
      patterns[38418] = 29'b1_001011000010_010_0_010110000101;
      patterns[38419] = 29'b1_001011000010_011_0_101100001010;
      patterns[38420] = 29'b1_001011000010_100_0_100101100001;
      patterns[38421] = 29'b1_001011000010_101_1_010010110000;
      patterns[38422] = 29'b1_001011000010_110_1_001011000010;
      patterns[38423] = 29'b1_001011000010_111_1_001011000010;
      patterns[38424] = 29'b1_001011000011_000_1_001011000011;
      patterns[38425] = 29'b1_001011000011_001_1_000011001011;
      patterns[38426] = 29'b1_001011000011_010_0_010110000111;
      patterns[38427] = 29'b1_001011000011_011_0_101100001110;
      patterns[38428] = 29'b1_001011000011_100_1_100101100001;
      patterns[38429] = 29'b1_001011000011_101_1_110010110000;
      patterns[38430] = 29'b1_001011000011_110_1_001011000011;
      patterns[38431] = 29'b1_001011000011_111_1_001011000011;
      patterns[38432] = 29'b1_001011000100_000_1_001011000100;
      patterns[38433] = 29'b1_001011000100_001_1_000100001011;
      patterns[38434] = 29'b1_001011000100_010_0_010110001001;
      patterns[38435] = 29'b1_001011000100_011_0_101100010010;
      patterns[38436] = 29'b1_001011000100_100_0_100101100010;
      patterns[38437] = 29'b1_001011000100_101_0_010010110001;
      patterns[38438] = 29'b1_001011000100_110_1_001011000100;
      patterns[38439] = 29'b1_001011000100_111_1_001011000100;
      patterns[38440] = 29'b1_001011000101_000_1_001011000101;
      patterns[38441] = 29'b1_001011000101_001_1_000101001011;
      patterns[38442] = 29'b1_001011000101_010_0_010110001011;
      patterns[38443] = 29'b1_001011000101_011_0_101100010110;
      patterns[38444] = 29'b1_001011000101_100_1_100101100010;
      patterns[38445] = 29'b1_001011000101_101_0_110010110001;
      patterns[38446] = 29'b1_001011000101_110_1_001011000101;
      patterns[38447] = 29'b1_001011000101_111_1_001011000101;
      patterns[38448] = 29'b1_001011000110_000_1_001011000110;
      patterns[38449] = 29'b1_001011000110_001_1_000110001011;
      patterns[38450] = 29'b1_001011000110_010_0_010110001101;
      patterns[38451] = 29'b1_001011000110_011_0_101100011010;
      patterns[38452] = 29'b1_001011000110_100_0_100101100011;
      patterns[38453] = 29'b1_001011000110_101_1_010010110001;
      patterns[38454] = 29'b1_001011000110_110_1_001011000110;
      patterns[38455] = 29'b1_001011000110_111_1_001011000110;
      patterns[38456] = 29'b1_001011000111_000_1_001011000111;
      patterns[38457] = 29'b1_001011000111_001_1_000111001011;
      patterns[38458] = 29'b1_001011000111_010_0_010110001111;
      patterns[38459] = 29'b1_001011000111_011_0_101100011110;
      patterns[38460] = 29'b1_001011000111_100_1_100101100011;
      patterns[38461] = 29'b1_001011000111_101_1_110010110001;
      patterns[38462] = 29'b1_001011000111_110_1_001011000111;
      patterns[38463] = 29'b1_001011000111_111_1_001011000111;
      patterns[38464] = 29'b1_001011001000_000_1_001011001000;
      patterns[38465] = 29'b1_001011001000_001_1_001000001011;
      patterns[38466] = 29'b1_001011001000_010_0_010110010001;
      patterns[38467] = 29'b1_001011001000_011_0_101100100010;
      patterns[38468] = 29'b1_001011001000_100_0_100101100100;
      patterns[38469] = 29'b1_001011001000_101_0_010010110010;
      patterns[38470] = 29'b1_001011001000_110_1_001011001000;
      patterns[38471] = 29'b1_001011001000_111_1_001011001000;
      patterns[38472] = 29'b1_001011001001_000_1_001011001001;
      patterns[38473] = 29'b1_001011001001_001_1_001001001011;
      patterns[38474] = 29'b1_001011001001_010_0_010110010011;
      patterns[38475] = 29'b1_001011001001_011_0_101100100110;
      patterns[38476] = 29'b1_001011001001_100_1_100101100100;
      patterns[38477] = 29'b1_001011001001_101_0_110010110010;
      patterns[38478] = 29'b1_001011001001_110_1_001011001001;
      patterns[38479] = 29'b1_001011001001_111_1_001011001001;
      patterns[38480] = 29'b1_001011001010_000_1_001011001010;
      patterns[38481] = 29'b1_001011001010_001_1_001010001011;
      patterns[38482] = 29'b1_001011001010_010_0_010110010101;
      patterns[38483] = 29'b1_001011001010_011_0_101100101010;
      patterns[38484] = 29'b1_001011001010_100_0_100101100101;
      patterns[38485] = 29'b1_001011001010_101_1_010010110010;
      patterns[38486] = 29'b1_001011001010_110_1_001011001010;
      patterns[38487] = 29'b1_001011001010_111_1_001011001010;
      patterns[38488] = 29'b1_001011001011_000_1_001011001011;
      patterns[38489] = 29'b1_001011001011_001_1_001011001011;
      patterns[38490] = 29'b1_001011001011_010_0_010110010111;
      patterns[38491] = 29'b1_001011001011_011_0_101100101110;
      patterns[38492] = 29'b1_001011001011_100_1_100101100101;
      patterns[38493] = 29'b1_001011001011_101_1_110010110010;
      patterns[38494] = 29'b1_001011001011_110_1_001011001011;
      patterns[38495] = 29'b1_001011001011_111_1_001011001011;
      patterns[38496] = 29'b1_001011001100_000_1_001011001100;
      patterns[38497] = 29'b1_001011001100_001_1_001100001011;
      patterns[38498] = 29'b1_001011001100_010_0_010110011001;
      patterns[38499] = 29'b1_001011001100_011_0_101100110010;
      patterns[38500] = 29'b1_001011001100_100_0_100101100110;
      patterns[38501] = 29'b1_001011001100_101_0_010010110011;
      patterns[38502] = 29'b1_001011001100_110_1_001011001100;
      patterns[38503] = 29'b1_001011001100_111_1_001011001100;
      patterns[38504] = 29'b1_001011001101_000_1_001011001101;
      patterns[38505] = 29'b1_001011001101_001_1_001101001011;
      patterns[38506] = 29'b1_001011001101_010_0_010110011011;
      patterns[38507] = 29'b1_001011001101_011_0_101100110110;
      patterns[38508] = 29'b1_001011001101_100_1_100101100110;
      patterns[38509] = 29'b1_001011001101_101_0_110010110011;
      patterns[38510] = 29'b1_001011001101_110_1_001011001101;
      patterns[38511] = 29'b1_001011001101_111_1_001011001101;
      patterns[38512] = 29'b1_001011001110_000_1_001011001110;
      patterns[38513] = 29'b1_001011001110_001_1_001110001011;
      patterns[38514] = 29'b1_001011001110_010_0_010110011101;
      patterns[38515] = 29'b1_001011001110_011_0_101100111010;
      patterns[38516] = 29'b1_001011001110_100_0_100101100111;
      patterns[38517] = 29'b1_001011001110_101_1_010010110011;
      patterns[38518] = 29'b1_001011001110_110_1_001011001110;
      patterns[38519] = 29'b1_001011001110_111_1_001011001110;
      patterns[38520] = 29'b1_001011001111_000_1_001011001111;
      patterns[38521] = 29'b1_001011001111_001_1_001111001011;
      patterns[38522] = 29'b1_001011001111_010_0_010110011111;
      patterns[38523] = 29'b1_001011001111_011_0_101100111110;
      patterns[38524] = 29'b1_001011001111_100_1_100101100111;
      patterns[38525] = 29'b1_001011001111_101_1_110010110011;
      patterns[38526] = 29'b1_001011001111_110_1_001011001111;
      patterns[38527] = 29'b1_001011001111_111_1_001011001111;
      patterns[38528] = 29'b1_001011010000_000_1_001011010000;
      patterns[38529] = 29'b1_001011010000_001_1_010000001011;
      patterns[38530] = 29'b1_001011010000_010_0_010110100001;
      patterns[38531] = 29'b1_001011010000_011_0_101101000010;
      patterns[38532] = 29'b1_001011010000_100_0_100101101000;
      patterns[38533] = 29'b1_001011010000_101_0_010010110100;
      patterns[38534] = 29'b1_001011010000_110_1_001011010000;
      patterns[38535] = 29'b1_001011010000_111_1_001011010000;
      patterns[38536] = 29'b1_001011010001_000_1_001011010001;
      patterns[38537] = 29'b1_001011010001_001_1_010001001011;
      patterns[38538] = 29'b1_001011010001_010_0_010110100011;
      patterns[38539] = 29'b1_001011010001_011_0_101101000110;
      patterns[38540] = 29'b1_001011010001_100_1_100101101000;
      patterns[38541] = 29'b1_001011010001_101_0_110010110100;
      patterns[38542] = 29'b1_001011010001_110_1_001011010001;
      patterns[38543] = 29'b1_001011010001_111_1_001011010001;
      patterns[38544] = 29'b1_001011010010_000_1_001011010010;
      patterns[38545] = 29'b1_001011010010_001_1_010010001011;
      patterns[38546] = 29'b1_001011010010_010_0_010110100101;
      patterns[38547] = 29'b1_001011010010_011_0_101101001010;
      patterns[38548] = 29'b1_001011010010_100_0_100101101001;
      patterns[38549] = 29'b1_001011010010_101_1_010010110100;
      patterns[38550] = 29'b1_001011010010_110_1_001011010010;
      patterns[38551] = 29'b1_001011010010_111_1_001011010010;
      patterns[38552] = 29'b1_001011010011_000_1_001011010011;
      patterns[38553] = 29'b1_001011010011_001_1_010011001011;
      patterns[38554] = 29'b1_001011010011_010_0_010110100111;
      patterns[38555] = 29'b1_001011010011_011_0_101101001110;
      patterns[38556] = 29'b1_001011010011_100_1_100101101001;
      patterns[38557] = 29'b1_001011010011_101_1_110010110100;
      patterns[38558] = 29'b1_001011010011_110_1_001011010011;
      patterns[38559] = 29'b1_001011010011_111_1_001011010011;
      patterns[38560] = 29'b1_001011010100_000_1_001011010100;
      patterns[38561] = 29'b1_001011010100_001_1_010100001011;
      patterns[38562] = 29'b1_001011010100_010_0_010110101001;
      patterns[38563] = 29'b1_001011010100_011_0_101101010010;
      patterns[38564] = 29'b1_001011010100_100_0_100101101010;
      patterns[38565] = 29'b1_001011010100_101_0_010010110101;
      patterns[38566] = 29'b1_001011010100_110_1_001011010100;
      patterns[38567] = 29'b1_001011010100_111_1_001011010100;
      patterns[38568] = 29'b1_001011010101_000_1_001011010101;
      patterns[38569] = 29'b1_001011010101_001_1_010101001011;
      patterns[38570] = 29'b1_001011010101_010_0_010110101011;
      patterns[38571] = 29'b1_001011010101_011_0_101101010110;
      patterns[38572] = 29'b1_001011010101_100_1_100101101010;
      patterns[38573] = 29'b1_001011010101_101_0_110010110101;
      patterns[38574] = 29'b1_001011010101_110_1_001011010101;
      patterns[38575] = 29'b1_001011010101_111_1_001011010101;
      patterns[38576] = 29'b1_001011010110_000_1_001011010110;
      patterns[38577] = 29'b1_001011010110_001_1_010110001011;
      patterns[38578] = 29'b1_001011010110_010_0_010110101101;
      patterns[38579] = 29'b1_001011010110_011_0_101101011010;
      patterns[38580] = 29'b1_001011010110_100_0_100101101011;
      patterns[38581] = 29'b1_001011010110_101_1_010010110101;
      patterns[38582] = 29'b1_001011010110_110_1_001011010110;
      patterns[38583] = 29'b1_001011010110_111_1_001011010110;
      patterns[38584] = 29'b1_001011010111_000_1_001011010111;
      patterns[38585] = 29'b1_001011010111_001_1_010111001011;
      patterns[38586] = 29'b1_001011010111_010_0_010110101111;
      patterns[38587] = 29'b1_001011010111_011_0_101101011110;
      patterns[38588] = 29'b1_001011010111_100_1_100101101011;
      patterns[38589] = 29'b1_001011010111_101_1_110010110101;
      patterns[38590] = 29'b1_001011010111_110_1_001011010111;
      patterns[38591] = 29'b1_001011010111_111_1_001011010111;
      patterns[38592] = 29'b1_001011011000_000_1_001011011000;
      patterns[38593] = 29'b1_001011011000_001_1_011000001011;
      patterns[38594] = 29'b1_001011011000_010_0_010110110001;
      patterns[38595] = 29'b1_001011011000_011_0_101101100010;
      patterns[38596] = 29'b1_001011011000_100_0_100101101100;
      patterns[38597] = 29'b1_001011011000_101_0_010010110110;
      patterns[38598] = 29'b1_001011011000_110_1_001011011000;
      patterns[38599] = 29'b1_001011011000_111_1_001011011000;
      patterns[38600] = 29'b1_001011011001_000_1_001011011001;
      patterns[38601] = 29'b1_001011011001_001_1_011001001011;
      patterns[38602] = 29'b1_001011011001_010_0_010110110011;
      patterns[38603] = 29'b1_001011011001_011_0_101101100110;
      patterns[38604] = 29'b1_001011011001_100_1_100101101100;
      patterns[38605] = 29'b1_001011011001_101_0_110010110110;
      patterns[38606] = 29'b1_001011011001_110_1_001011011001;
      patterns[38607] = 29'b1_001011011001_111_1_001011011001;
      patterns[38608] = 29'b1_001011011010_000_1_001011011010;
      patterns[38609] = 29'b1_001011011010_001_1_011010001011;
      patterns[38610] = 29'b1_001011011010_010_0_010110110101;
      patterns[38611] = 29'b1_001011011010_011_0_101101101010;
      patterns[38612] = 29'b1_001011011010_100_0_100101101101;
      patterns[38613] = 29'b1_001011011010_101_1_010010110110;
      patterns[38614] = 29'b1_001011011010_110_1_001011011010;
      patterns[38615] = 29'b1_001011011010_111_1_001011011010;
      patterns[38616] = 29'b1_001011011011_000_1_001011011011;
      patterns[38617] = 29'b1_001011011011_001_1_011011001011;
      patterns[38618] = 29'b1_001011011011_010_0_010110110111;
      patterns[38619] = 29'b1_001011011011_011_0_101101101110;
      patterns[38620] = 29'b1_001011011011_100_1_100101101101;
      patterns[38621] = 29'b1_001011011011_101_1_110010110110;
      patterns[38622] = 29'b1_001011011011_110_1_001011011011;
      patterns[38623] = 29'b1_001011011011_111_1_001011011011;
      patterns[38624] = 29'b1_001011011100_000_1_001011011100;
      patterns[38625] = 29'b1_001011011100_001_1_011100001011;
      patterns[38626] = 29'b1_001011011100_010_0_010110111001;
      patterns[38627] = 29'b1_001011011100_011_0_101101110010;
      patterns[38628] = 29'b1_001011011100_100_0_100101101110;
      patterns[38629] = 29'b1_001011011100_101_0_010010110111;
      patterns[38630] = 29'b1_001011011100_110_1_001011011100;
      patterns[38631] = 29'b1_001011011100_111_1_001011011100;
      patterns[38632] = 29'b1_001011011101_000_1_001011011101;
      patterns[38633] = 29'b1_001011011101_001_1_011101001011;
      patterns[38634] = 29'b1_001011011101_010_0_010110111011;
      patterns[38635] = 29'b1_001011011101_011_0_101101110110;
      patterns[38636] = 29'b1_001011011101_100_1_100101101110;
      patterns[38637] = 29'b1_001011011101_101_0_110010110111;
      patterns[38638] = 29'b1_001011011101_110_1_001011011101;
      patterns[38639] = 29'b1_001011011101_111_1_001011011101;
      patterns[38640] = 29'b1_001011011110_000_1_001011011110;
      patterns[38641] = 29'b1_001011011110_001_1_011110001011;
      patterns[38642] = 29'b1_001011011110_010_0_010110111101;
      patterns[38643] = 29'b1_001011011110_011_0_101101111010;
      patterns[38644] = 29'b1_001011011110_100_0_100101101111;
      patterns[38645] = 29'b1_001011011110_101_1_010010110111;
      patterns[38646] = 29'b1_001011011110_110_1_001011011110;
      patterns[38647] = 29'b1_001011011110_111_1_001011011110;
      patterns[38648] = 29'b1_001011011111_000_1_001011011111;
      patterns[38649] = 29'b1_001011011111_001_1_011111001011;
      patterns[38650] = 29'b1_001011011111_010_0_010110111111;
      patterns[38651] = 29'b1_001011011111_011_0_101101111110;
      patterns[38652] = 29'b1_001011011111_100_1_100101101111;
      patterns[38653] = 29'b1_001011011111_101_1_110010110111;
      patterns[38654] = 29'b1_001011011111_110_1_001011011111;
      patterns[38655] = 29'b1_001011011111_111_1_001011011111;
      patterns[38656] = 29'b1_001011100000_000_1_001011100000;
      patterns[38657] = 29'b1_001011100000_001_1_100000001011;
      patterns[38658] = 29'b1_001011100000_010_0_010111000001;
      patterns[38659] = 29'b1_001011100000_011_0_101110000010;
      patterns[38660] = 29'b1_001011100000_100_0_100101110000;
      patterns[38661] = 29'b1_001011100000_101_0_010010111000;
      patterns[38662] = 29'b1_001011100000_110_1_001011100000;
      patterns[38663] = 29'b1_001011100000_111_1_001011100000;
      patterns[38664] = 29'b1_001011100001_000_1_001011100001;
      patterns[38665] = 29'b1_001011100001_001_1_100001001011;
      patterns[38666] = 29'b1_001011100001_010_0_010111000011;
      patterns[38667] = 29'b1_001011100001_011_0_101110000110;
      patterns[38668] = 29'b1_001011100001_100_1_100101110000;
      patterns[38669] = 29'b1_001011100001_101_0_110010111000;
      patterns[38670] = 29'b1_001011100001_110_1_001011100001;
      patterns[38671] = 29'b1_001011100001_111_1_001011100001;
      patterns[38672] = 29'b1_001011100010_000_1_001011100010;
      patterns[38673] = 29'b1_001011100010_001_1_100010001011;
      patterns[38674] = 29'b1_001011100010_010_0_010111000101;
      patterns[38675] = 29'b1_001011100010_011_0_101110001010;
      patterns[38676] = 29'b1_001011100010_100_0_100101110001;
      patterns[38677] = 29'b1_001011100010_101_1_010010111000;
      patterns[38678] = 29'b1_001011100010_110_1_001011100010;
      patterns[38679] = 29'b1_001011100010_111_1_001011100010;
      patterns[38680] = 29'b1_001011100011_000_1_001011100011;
      patterns[38681] = 29'b1_001011100011_001_1_100011001011;
      patterns[38682] = 29'b1_001011100011_010_0_010111000111;
      patterns[38683] = 29'b1_001011100011_011_0_101110001110;
      patterns[38684] = 29'b1_001011100011_100_1_100101110001;
      patterns[38685] = 29'b1_001011100011_101_1_110010111000;
      patterns[38686] = 29'b1_001011100011_110_1_001011100011;
      patterns[38687] = 29'b1_001011100011_111_1_001011100011;
      patterns[38688] = 29'b1_001011100100_000_1_001011100100;
      patterns[38689] = 29'b1_001011100100_001_1_100100001011;
      patterns[38690] = 29'b1_001011100100_010_0_010111001001;
      patterns[38691] = 29'b1_001011100100_011_0_101110010010;
      patterns[38692] = 29'b1_001011100100_100_0_100101110010;
      patterns[38693] = 29'b1_001011100100_101_0_010010111001;
      patterns[38694] = 29'b1_001011100100_110_1_001011100100;
      patterns[38695] = 29'b1_001011100100_111_1_001011100100;
      patterns[38696] = 29'b1_001011100101_000_1_001011100101;
      patterns[38697] = 29'b1_001011100101_001_1_100101001011;
      patterns[38698] = 29'b1_001011100101_010_0_010111001011;
      patterns[38699] = 29'b1_001011100101_011_0_101110010110;
      patterns[38700] = 29'b1_001011100101_100_1_100101110010;
      patterns[38701] = 29'b1_001011100101_101_0_110010111001;
      patterns[38702] = 29'b1_001011100101_110_1_001011100101;
      patterns[38703] = 29'b1_001011100101_111_1_001011100101;
      patterns[38704] = 29'b1_001011100110_000_1_001011100110;
      patterns[38705] = 29'b1_001011100110_001_1_100110001011;
      patterns[38706] = 29'b1_001011100110_010_0_010111001101;
      patterns[38707] = 29'b1_001011100110_011_0_101110011010;
      patterns[38708] = 29'b1_001011100110_100_0_100101110011;
      patterns[38709] = 29'b1_001011100110_101_1_010010111001;
      patterns[38710] = 29'b1_001011100110_110_1_001011100110;
      patterns[38711] = 29'b1_001011100110_111_1_001011100110;
      patterns[38712] = 29'b1_001011100111_000_1_001011100111;
      patterns[38713] = 29'b1_001011100111_001_1_100111001011;
      patterns[38714] = 29'b1_001011100111_010_0_010111001111;
      patterns[38715] = 29'b1_001011100111_011_0_101110011110;
      patterns[38716] = 29'b1_001011100111_100_1_100101110011;
      patterns[38717] = 29'b1_001011100111_101_1_110010111001;
      patterns[38718] = 29'b1_001011100111_110_1_001011100111;
      patterns[38719] = 29'b1_001011100111_111_1_001011100111;
      patterns[38720] = 29'b1_001011101000_000_1_001011101000;
      patterns[38721] = 29'b1_001011101000_001_1_101000001011;
      patterns[38722] = 29'b1_001011101000_010_0_010111010001;
      patterns[38723] = 29'b1_001011101000_011_0_101110100010;
      patterns[38724] = 29'b1_001011101000_100_0_100101110100;
      patterns[38725] = 29'b1_001011101000_101_0_010010111010;
      patterns[38726] = 29'b1_001011101000_110_1_001011101000;
      patterns[38727] = 29'b1_001011101000_111_1_001011101000;
      patterns[38728] = 29'b1_001011101001_000_1_001011101001;
      patterns[38729] = 29'b1_001011101001_001_1_101001001011;
      patterns[38730] = 29'b1_001011101001_010_0_010111010011;
      patterns[38731] = 29'b1_001011101001_011_0_101110100110;
      patterns[38732] = 29'b1_001011101001_100_1_100101110100;
      patterns[38733] = 29'b1_001011101001_101_0_110010111010;
      patterns[38734] = 29'b1_001011101001_110_1_001011101001;
      patterns[38735] = 29'b1_001011101001_111_1_001011101001;
      patterns[38736] = 29'b1_001011101010_000_1_001011101010;
      patterns[38737] = 29'b1_001011101010_001_1_101010001011;
      patterns[38738] = 29'b1_001011101010_010_0_010111010101;
      patterns[38739] = 29'b1_001011101010_011_0_101110101010;
      patterns[38740] = 29'b1_001011101010_100_0_100101110101;
      patterns[38741] = 29'b1_001011101010_101_1_010010111010;
      patterns[38742] = 29'b1_001011101010_110_1_001011101010;
      patterns[38743] = 29'b1_001011101010_111_1_001011101010;
      patterns[38744] = 29'b1_001011101011_000_1_001011101011;
      patterns[38745] = 29'b1_001011101011_001_1_101011001011;
      patterns[38746] = 29'b1_001011101011_010_0_010111010111;
      patterns[38747] = 29'b1_001011101011_011_0_101110101110;
      patterns[38748] = 29'b1_001011101011_100_1_100101110101;
      patterns[38749] = 29'b1_001011101011_101_1_110010111010;
      patterns[38750] = 29'b1_001011101011_110_1_001011101011;
      patterns[38751] = 29'b1_001011101011_111_1_001011101011;
      patterns[38752] = 29'b1_001011101100_000_1_001011101100;
      patterns[38753] = 29'b1_001011101100_001_1_101100001011;
      patterns[38754] = 29'b1_001011101100_010_0_010111011001;
      patterns[38755] = 29'b1_001011101100_011_0_101110110010;
      patterns[38756] = 29'b1_001011101100_100_0_100101110110;
      patterns[38757] = 29'b1_001011101100_101_0_010010111011;
      patterns[38758] = 29'b1_001011101100_110_1_001011101100;
      patterns[38759] = 29'b1_001011101100_111_1_001011101100;
      patterns[38760] = 29'b1_001011101101_000_1_001011101101;
      patterns[38761] = 29'b1_001011101101_001_1_101101001011;
      patterns[38762] = 29'b1_001011101101_010_0_010111011011;
      patterns[38763] = 29'b1_001011101101_011_0_101110110110;
      patterns[38764] = 29'b1_001011101101_100_1_100101110110;
      patterns[38765] = 29'b1_001011101101_101_0_110010111011;
      patterns[38766] = 29'b1_001011101101_110_1_001011101101;
      patterns[38767] = 29'b1_001011101101_111_1_001011101101;
      patterns[38768] = 29'b1_001011101110_000_1_001011101110;
      patterns[38769] = 29'b1_001011101110_001_1_101110001011;
      patterns[38770] = 29'b1_001011101110_010_0_010111011101;
      patterns[38771] = 29'b1_001011101110_011_0_101110111010;
      patterns[38772] = 29'b1_001011101110_100_0_100101110111;
      patterns[38773] = 29'b1_001011101110_101_1_010010111011;
      patterns[38774] = 29'b1_001011101110_110_1_001011101110;
      patterns[38775] = 29'b1_001011101110_111_1_001011101110;
      patterns[38776] = 29'b1_001011101111_000_1_001011101111;
      patterns[38777] = 29'b1_001011101111_001_1_101111001011;
      patterns[38778] = 29'b1_001011101111_010_0_010111011111;
      patterns[38779] = 29'b1_001011101111_011_0_101110111110;
      patterns[38780] = 29'b1_001011101111_100_1_100101110111;
      patterns[38781] = 29'b1_001011101111_101_1_110010111011;
      patterns[38782] = 29'b1_001011101111_110_1_001011101111;
      patterns[38783] = 29'b1_001011101111_111_1_001011101111;
      patterns[38784] = 29'b1_001011110000_000_1_001011110000;
      patterns[38785] = 29'b1_001011110000_001_1_110000001011;
      patterns[38786] = 29'b1_001011110000_010_0_010111100001;
      patterns[38787] = 29'b1_001011110000_011_0_101111000010;
      patterns[38788] = 29'b1_001011110000_100_0_100101111000;
      patterns[38789] = 29'b1_001011110000_101_0_010010111100;
      patterns[38790] = 29'b1_001011110000_110_1_001011110000;
      patterns[38791] = 29'b1_001011110000_111_1_001011110000;
      patterns[38792] = 29'b1_001011110001_000_1_001011110001;
      patterns[38793] = 29'b1_001011110001_001_1_110001001011;
      patterns[38794] = 29'b1_001011110001_010_0_010111100011;
      patterns[38795] = 29'b1_001011110001_011_0_101111000110;
      patterns[38796] = 29'b1_001011110001_100_1_100101111000;
      patterns[38797] = 29'b1_001011110001_101_0_110010111100;
      patterns[38798] = 29'b1_001011110001_110_1_001011110001;
      patterns[38799] = 29'b1_001011110001_111_1_001011110001;
      patterns[38800] = 29'b1_001011110010_000_1_001011110010;
      patterns[38801] = 29'b1_001011110010_001_1_110010001011;
      patterns[38802] = 29'b1_001011110010_010_0_010111100101;
      patterns[38803] = 29'b1_001011110010_011_0_101111001010;
      patterns[38804] = 29'b1_001011110010_100_0_100101111001;
      patterns[38805] = 29'b1_001011110010_101_1_010010111100;
      patterns[38806] = 29'b1_001011110010_110_1_001011110010;
      patterns[38807] = 29'b1_001011110010_111_1_001011110010;
      patterns[38808] = 29'b1_001011110011_000_1_001011110011;
      patterns[38809] = 29'b1_001011110011_001_1_110011001011;
      patterns[38810] = 29'b1_001011110011_010_0_010111100111;
      patterns[38811] = 29'b1_001011110011_011_0_101111001110;
      patterns[38812] = 29'b1_001011110011_100_1_100101111001;
      patterns[38813] = 29'b1_001011110011_101_1_110010111100;
      patterns[38814] = 29'b1_001011110011_110_1_001011110011;
      patterns[38815] = 29'b1_001011110011_111_1_001011110011;
      patterns[38816] = 29'b1_001011110100_000_1_001011110100;
      patterns[38817] = 29'b1_001011110100_001_1_110100001011;
      patterns[38818] = 29'b1_001011110100_010_0_010111101001;
      patterns[38819] = 29'b1_001011110100_011_0_101111010010;
      patterns[38820] = 29'b1_001011110100_100_0_100101111010;
      patterns[38821] = 29'b1_001011110100_101_0_010010111101;
      patterns[38822] = 29'b1_001011110100_110_1_001011110100;
      patterns[38823] = 29'b1_001011110100_111_1_001011110100;
      patterns[38824] = 29'b1_001011110101_000_1_001011110101;
      patterns[38825] = 29'b1_001011110101_001_1_110101001011;
      patterns[38826] = 29'b1_001011110101_010_0_010111101011;
      patterns[38827] = 29'b1_001011110101_011_0_101111010110;
      patterns[38828] = 29'b1_001011110101_100_1_100101111010;
      patterns[38829] = 29'b1_001011110101_101_0_110010111101;
      patterns[38830] = 29'b1_001011110101_110_1_001011110101;
      patterns[38831] = 29'b1_001011110101_111_1_001011110101;
      patterns[38832] = 29'b1_001011110110_000_1_001011110110;
      patterns[38833] = 29'b1_001011110110_001_1_110110001011;
      patterns[38834] = 29'b1_001011110110_010_0_010111101101;
      patterns[38835] = 29'b1_001011110110_011_0_101111011010;
      patterns[38836] = 29'b1_001011110110_100_0_100101111011;
      patterns[38837] = 29'b1_001011110110_101_1_010010111101;
      patterns[38838] = 29'b1_001011110110_110_1_001011110110;
      patterns[38839] = 29'b1_001011110110_111_1_001011110110;
      patterns[38840] = 29'b1_001011110111_000_1_001011110111;
      patterns[38841] = 29'b1_001011110111_001_1_110111001011;
      patterns[38842] = 29'b1_001011110111_010_0_010111101111;
      patterns[38843] = 29'b1_001011110111_011_0_101111011110;
      patterns[38844] = 29'b1_001011110111_100_1_100101111011;
      patterns[38845] = 29'b1_001011110111_101_1_110010111101;
      patterns[38846] = 29'b1_001011110111_110_1_001011110111;
      patterns[38847] = 29'b1_001011110111_111_1_001011110111;
      patterns[38848] = 29'b1_001011111000_000_1_001011111000;
      patterns[38849] = 29'b1_001011111000_001_1_111000001011;
      patterns[38850] = 29'b1_001011111000_010_0_010111110001;
      patterns[38851] = 29'b1_001011111000_011_0_101111100010;
      patterns[38852] = 29'b1_001011111000_100_0_100101111100;
      patterns[38853] = 29'b1_001011111000_101_0_010010111110;
      patterns[38854] = 29'b1_001011111000_110_1_001011111000;
      patterns[38855] = 29'b1_001011111000_111_1_001011111000;
      patterns[38856] = 29'b1_001011111001_000_1_001011111001;
      patterns[38857] = 29'b1_001011111001_001_1_111001001011;
      patterns[38858] = 29'b1_001011111001_010_0_010111110011;
      patterns[38859] = 29'b1_001011111001_011_0_101111100110;
      patterns[38860] = 29'b1_001011111001_100_1_100101111100;
      patterns[38861] = 29'b1_001011111001_101_0_110010111110;
      patterns[38862] = 29'b1_001011111001_110_1_001011111001;
      patterns[38863] = 29'b1_001011111001_111_1_001011111001;
      patterns[38864] = 29'b1_001011111010_000_1_001011111010;
      patterns[38865] = 29'b1_001011111010_001_1_111010001011;
      patterns[38866] = 29'b1_001011111010_010_0_010111110101;
      patterns[38867] = 29'b1_001011111010_011_0_101111101010;
      patterns[38868] = 29'b1_001011111010_100_0_100101111101;
      patterns[38869] = 29'b1_001011111010_101_1_010010111110;
      patterns[38870] = 29'b1_001011111010_110_1_001011111010;
      patterns[38871] = 29'b1_001011111010_111_1_001011111010;
      patterns[38872] = 29'b1_001011111011_000_1_001011111011;
      patterns[38873] = 29'b1_001011111011_001_1_111011001011;
      patterns[38874] = 29'b1_001011111011_010_0_010111110111;
      patterns[38875] = 29'b1_001011111011_011_0_101111101110;
      patterns[38876] = 29'b1_001011111011_100_1_100101111101;
      patterns[38877] = 29'b1_001011111011_101_1_110010111110;
      patterns[38878] = 29'b1_001011111011_110_1_001011111011;
      patterns[38879] = 29'b1_001011111011_111_1_001011111011;
      patterns[38880] = 29'b1_001011111100_000_1_001011111100;
      patterns[38881] = 29'b1_001011111100_001_1_111100001011;
      patterns[38882] = 29'b1_001011111100_010_0_010111111001;
      patterns[38883] = 29'b1_001011111100_011_0_101111110010;
      patterns[38884] = 29'b1_001011111100_100_0_100101111110;
      patterns[38885] = 29'b1_001011111100_101_0_010010111111;
      patterns[38886] = 29'b1_001011111100_110_1_001011111100;
      patterns[38887] = 29'b1_001011111100_111_1_001011111100;
      patterns[38888] = 29'b1_001011111101_000_1_001011111101;
      patterns[38889] = 29'b1_001011111101_001_1_111101001011;
      patterns[38890] = 29'b1_001011111101_010_0_010111111011;
      patterns[38891] = 29'b1_001011111101_011_0_101111110110;
      patterns[38892] = 29'b1_001011111101_100_1_100101111110;
      patterns[38893] = 29'b1_001011111101_101_0_110010111111;
      patterns[38894] = 29'b1_001011111101_110_1_001011111101;
      patterns[38895] = 29'b1_001011111101_111_1_001011111101;
      patterns[38896] = 29'b1_001011111110_000_1_001011111110;
      patterns[38897] = 29'b1_001011111110_001_1_111110001011;
      patterns[38898] = 29'b1_001011111110_010_0_010111111101;
      patterns[38899] = 29'b1_001011111110_011_0_101111111010;
      patterns[38900] = 29'b1_001011111110_100_0_100101111111;
      patterns[38901] = 29'b1_001011111110_101_1_010010111111;
      patterns[38902] = 29'b1_001011111110_110_1_001011111110;
      patterns[38903] = 29'b1_001011111110_111_1_001011111110;
      patterns[38904] = 29'b1_001011111111_000_1_001011111111;
      patterns[38905] = 29'b1_001011111111_001_1_111111001011;
      patterns[38906] = 29'b1_001011111111_010_0_010111111111;
      patterns[38907] = 29'b1_001011111111_011_0_101111111110;
      patterns[38908] = 29'b1_001011111111_100_1_100101111111;
      patterns[38909] = 29'b1_001011111111_101_1_110010111111;
      patterns[38910] = 29'b1_001011111111_110_1_001011111111;
      patterns[38911] = 29'b1_001011111111_111_1_001011111111;
      patterns[38912] = 29'b1_001100000000_000_1_001100000000;
      patterns[38913] = 29'b1_001100000000_001_1_000000001100;
      patterns[38914] = 29'b1_001100000000_010_0_011000000001;
      patterns[38915] = 29'b1_001100000000_011_0_110000000010;
      patterns[38916] = 29'b1_001100000000_100_0_100110000000;
      patterns[38917] = 29'b1_001100000000_101_0_010011000000;
      patterns[38918] = 29'b1_001100000000_110_1_001100000000;
      patterns[38919] = 29'b1_001100000000_111_1_001100000000;
      patterns[38920] = 29'b1_001100000001_000_1_001100000001;
      patterns[38921] = 29'b1_001100000001_001_1_000001001100;
      patterns[38922] = 29'b1_001100000001_010_0_011000000011;
      patterns[38923] = 29'b1_001100000001_011_0_110000000110;
      patterns[38924] = 29'b1_001100000001_100_1_100110000000;
      patterns[38925] = 29'b1_001100000001_101_0_110011000000;
      patterns[38926] = 29'b1_001100000001_110_1_001100000001;
      patterns[38927] = 29'b1_001100000001_111_1_001100000001;
      patterns[38928] = 29'b1_001100000010_000_1_001100000010;
      patterns[38929] = 29'b1_001100000010_001_1_000010001100;
      patterns[38930] = 29'b1_001100000010_010_0_011000000101;
      patterns[38931] = 29'b1_001100000010_011_0_110000001010;
      patterns[38932] = 29'b1_001100000010_100_0_100110000001;
      patterns[38933] = 29'b1_001100000010_101_1_010011000000;
      patterns[38934] = 29'b1_001100000010_110_1_001100000010;
      patterns[38935] = 29'b1_001100000010_111_1_001100000010;
      patterns[38936] = 29'b1_001100000011_000_1_001100000011;
      patterns[38937] = 29'b1_001100000011_001_1_000011001100;
      patterns[38938] = 29'b1_001100000011_010_0_011000000111;
      patterns[38939] = 29'b1_001100000011_011_0_110000001110;
      patterns[38940] = 29'b1_001100000011_100_1_100110000001;
      patterns[38941] = 29'b1_001100000011_101_1_110011000000;
      patterns[38942] = 29'b1_001100000011_110_1_001100000011;
      patterns[38943] = 29'b1_001100000011_111_1_001100000011;
      patterns[38944] = 29'b1_001100000100_000_1_001100000100;
      patterns[38945] = 29'b1_001100000100_001_1_000100001100;
      patterns[38946] = 29'b1_001100000100_010_0_011000001001;
      patterns[38947] = 29'b1_001100000100_011_0_110000010010;
      patterns[38948] = 29'b1_001100000100_100_0_100110000010;
      patterns[38949] = 29'b1_001100000100_101_0_010011000001;
      patterns[38950] = 29'b1_001100000100_110_1_001100000100;
      patterns[38951] = 29'b1_001100000100_111_1_001100000100;
      patterns[38952] = 29'b1_001100000101_000_1_001100000101;
      patterns[38953] = 29'b1_001100000101_001_1_000101001100;
      patterns[38954] = 29'b1_001100000101_010_0_011000001011;
      patterns[38955] = 29'b1_001100000101_011_0_110000010110;
      patterns[38956] = 29'b1_001100000101_100_1_100110000010;
      patterns[38957] = 29'b1_001100000101_101_0_110011000001;
      patterns[38958] = 29'b1_001100000101_110_1_001100000101;
      patterns[38959] = 29'b1_001100000101_111_1_001100000101;
      patterns[38960] = 29'b1_001100000110_000_1_001100000110;
      patterns[38961] = 29'b1_001100000110_001_1_000110001100;
      patterns[38962] = 29'b1_001100000110_010_0_011000001101;
      patterns[38963] = 29'b1_001100000110_011_0_110000011010;
      patterns[38964] = 29'b1_001100000110_100_0_100110000011;
      patterns[38965] = 29'b1_001100000110_101_1_010011000001;
      patterns[38966] = 29'b1_001100000110_110_1_001100000110;
      patterns[38967] = 29'b1_001100000110_111_1_001100000110;
      patterns[38968] = 29'b1_001100000111_000_1_001100000111;
      patterns[38969] = 29'b1_001100000111_001_1_000111001100;
      patterns[38970] = 29'b1_001100000111_010_0_011000001111;
      patterns[38971] = 29'b1_001100000111_011_0_110000011110;
      patterns[38972] = 29'b1_001100000111_100_1_100110000011;
      patterns[38973] = 29'b1_001100000111_101_1_110011000001;
      patterns[38974] = 29'b1_001100000111_110_1_001100000111;
      patterns[38975] = 29'b1_001100000111_111_1_001100000111;
      patterns[38976] = 29'b1_001100001000_000_1_001100001000;
      patterns[38977] = 29'b1_001100001000_001_1_001000001100;
      patterns[38978] = 29'b1_001100001000_010_0_011000010001;
      patterns[38979] = 29'b1_001100001000_011_0_110000100010;
      patterns[38980] = 29'b1_001100001000_100_0_100110000100;
      patterns[38981] = 29'b1_001100001000_101_0_010011000010;
      patterns[38982] = 29'b1_001100001000_110_1_001100001000;
      patterns[38983] = 29'b1_001100001000_111_1_001100001000;
      patterns[38984] = 29'b1_001100001001_000_1_001100001001;
      patterns[38985] = 29'b1_001100001001_001_1_001001001100;
      patterns[38986] = 29'b1_001100001001_010_0_011000010011;
      patterns[38987] = 29'b1_001100001001_011_0_110000100110;
      patterns[38988] = 29'b1_001100001001_100_1_100110000100;
      patterns[38989] = 29'b1_001100001001_101_0_110011000010;
      patterns[38990] = 29'b1_001100001001_110_1_001100001001;
      patterns[38991] = 29'b1_001100001001_111_1_001100001001;
      patterns[38992] = 29'b1_001100001010_000_1_001100001010;
      patterns[38993] = 29'b1_001100001010_001_1_001010001100;
      patterns[38994] = 29'b1_001100001010_010_0_011000010101;
      patterns[38995] = 29'b1_001100001010_011_0_110000101010;
      patterns[38996] = 29'b1_001100001010_100_0_100110000101;
      patterns[38997] = 29'b1_001100001010_101_1_010011000010;
      patterns[38998] = 29'b1_001100001010_110_1_001100001010;
      patterns[38999] = 29'b1_001100001010_111_1_001100001010;
      patterns[39000] = 29'b1_001100001011_000_1_001100001011;
      patterns[39001] = 29'b1_001100001011_001_1_001011001100;
      patterns[39002] = 29'b1_001100001011_010_0_011000010111;
      patterns[39003] = 29'b1_001100001011_011_0_110000101110;
      patterns[39004] = 29'b1_001100001011_100_1_100110000101;
      patterns[39005] = 29'b1_001100001011_101_1_110011000010;
      patterns[39006] = 29'b1_001100001011_110_1_001100001011;
      patterns[39007] = 29'b1_001100001011_111_1_001100001011;
      patterns[39008] = 29'b1_001100001100_000_1_001100001100;
      patterns[39009] = 29'b1_001100001100_001_1_001100001100;
      patterns[39010] = 29'b1_001100001100_010_0_011000011001;
      patterns[39011] = 29'b1_001100001100_011_0_110000110010;
      patterns[39012] = 29'b1_001100001100_100_0_100110000110;
      patterns[39013] = 29'b1_001100001100_101_0_010011000011;
      patterns[39014] = 29'b1_001100001100_110_1_001100001100;
      patterns[39015] = 29'b1_001100001100_111_1_001100001100;
      patterns[39016] = 29'b1_001100001101_000_1_001100001101;
      patterns[39017] = 29'b1_001100001101_001_1_001101001100;
      patterns[39018] = 29'b1_001100001101_010_0_011000011011;
      patterns[39019] = 29'b1_001100001101_011_0_110000110110;
      patterns[39020] = 29'b1_001100001101_100_1_100110000110;
      patterns[39021] = 29'b1_001100001101_101_0_110011000011;
      patterns[39022] = 29'b1_001100001101_110_1_001100001101;
      patterns[39023] = 29'b1_001100001101_111_1_001100001101;
      patterns[39024] = 29'b1_001100001110_000_1_001100001110;
      patterns[39025] = 29'b1_001100001110_001_1_001110001100;
      patterns[39026] = 29'b1_001100001110_010_0_011000011101;
      patterns[39027] = 29'b1_001100001110_011_0_110000111010;
      patterns[39028] = 29'b1_001100001110_100_0_100110000111;
      patterns[39029] = 29'b1_001100001110_101_1_010011000011;
      patterns[39030] = 29'b1_001100001110_110_1_001100001110;
      patterns[39031] = 29'b1_001100001110_111_1_001100001110;
      patterns[39032] = 29'b1_001100001111_000_1_001100001111;
      patterns[39033] = 29'b1_001100001111_001_1_001111001100;
      patterns[39034] = 29'b1_001100001111_010_0_011000011111;
      patterns[39035] = 29'b1_001100001111_011_0_110000111110;
      patterns[39036] = 29'b1_001100001111_100_1_100110000111;
      patterns[39037] = 29'b1_001100001111_101_1_110011000011;
      patterns[39038] = 29'b1_001100001111_110_1_001100001111;
      patterns[39039] = 29'b1_001100001111_111_1_001100001111;
      patterns[39040] = 29'b1_001100010000_000_1_001100010000;
      patterns[39041] = 29'b1_001100010000_001_1_010000001100;
      patterns[39042] = 29'b1_001100010000_010_0_011000100001;
      patterns[39043] = 29'b1_001100010000_011_0_110001000010;
      patterns[39044] = 29'b1_001100010000_100_0_100110001000;
      patterns[39045] = 29'b1_001100010000_101_0_010011000100;
      patterns[39046] = 29'b1_001100010000_110_1_001100010000;
      patterns[39047] = 29'b1_001100010000_111_1_001100010000;
      patterns[39048] = 29'b1_001100010001_000_1_001100010001;
      patterns[39049] = 29'b1_001100010001_001_1_010001001100;
      patterns[39050] = 29'b1_001100010001_010_0_011000100011;
      patterns[39051] = 29'b1_001100010001_011_0_110001000110;
      patterns[39052] = 29'b1_001100010001_100_1_100110001000;
      patterns[39053] = 29'b1_001100010001_101_0_110011000100;
      patterns[39054] = 29'b1_001100010001_110_1_001100010001;
      patterns[39055] = 29'b1_001100010001_111_1_001100010001;
      patterns[39056] = 29'b1_001100010010_000_1_001100010010;
      patterns[39057] = 29'b1_001100010010_001_1_010010001100;
      patterns[39058] = 29'b1_001100010010_010_0_011000100101;
      patterns[39059] = 29'b1_001100010010_011_0_110001001010;
      patterns[39060] = 29'b1_001100010010_100_0_100110001001;
      patterns[39061] = 29'b1_001100010010_101_1_010011000100;
      patterns[39062] = 29'b1_001100010010_110_1_001100010010;
      patterns[39063] = 29'b1_001100010010_111_1_001100010010;
      patterns[39064] = 29'b1_001100010011_000_1_001100010011;
      patterns[39065] = 29'b1_001100010011_001_1_010011001100;
      patterns[39066] = 29'b1_001100010011_010_0_011000100111;
      patterns[39067] = 29'b1_001100010011_011_0_110001001110;
      patterns[39068] = 29'b1_001100010011_100_1_100110001001;
      patterns[39069] = 29'b1_001100010011_101_1_110011000100;
      patterns[39070] = 29'b1_001100010011_110_1_001100010011;
      patterns[39071] = 29'b1_001100010011_111_1_001100010011;
      patterns[39072] = 29'b1_001100010100_000_1_001100010100;
      patterns[39073] = 29'b1_001100010100_001_1_010100001100;
      patterns[39074] = 29'b1_001100010100_010_0_011000101001;
      patterns[39075] = 29'b1_001100010100_011_0_110001010010;
      patterns[39076] = 29'b1_001100010100_100_0_100110001010;
      patterns[39077] = 29'b1_001100010100_101_0_010011000101;
      patterns[39078] = 29'b1_001100010100_110_1_001100010100;
      patterns[39079] = 29'b1_001100010100_111_1_001100010100;
      patterns[39080] = 29'b1_001100010101_000_1_001100010101;
      patterns[39081] = 29'b1_001100010101_001_1_010101001100;
      patterns[39082] = 29'b1_001100010101_010_0_011000101011;
      patterns[39083] = 29'b1_001100010101_011_0_110001010110;
      patterns[39084] = 29'b1_001100010101_100_1_100110001010;
      patterns[39085] = 29'b1_001100010101_101_0_110011000101;
      patterns[39086] = 29'b1_001100010101_110_1_001100010101;
      patterns[39087] = 29'b1_001100010101_111_1_001100010101;
      patterns[39088] = 29'b1_001100010110_000_1_001100010110;
      patterns[39089] = 29'b1_001100010110_001_1_010110001100;
      patterns[39090] = 29'b1_001100010110_010_0_011000101101;
      patterns[39091] = 29'b1_001100010110_011_0_110001011010;
      patterns[39092] = 29'b1_001100010110_100_0_100110001011;
      patterns[39093] = 29'b1_001100010110_101_1_010011000101;
      patterns[39094] = 29'b1_001100010110_110_1_001100010110;
      patterns[39095] = 29'b1_001100010110_111_1_001100010110;
      patterns[39096] = 29'b1_001100010111_000_1_001100010111;
      patterns[39097] = 29'b1_001100010111_001_1_010111001100;
      patterns[39098] = 29'b1_001100010111_010_0_011000101111;
      patterns[39099] = 29'b1_001100010111_011_0_110001011110;
      patterns[39100] = 29'b1_001100010111_100_1_100110001011;
      patterns[39101] = 29'b1_001100010111_101_1_110011000101;
      patterns[39102] = 29'b1_001100010111_110_1_001100010111;
      patterns[39103] = 29'b1_001100010111_111_1_001100010111;
      patterns[39104] = 29'b1_001100011000_000_1_001100011000;
      patterns[39105] = 29'b1_001100011000_001_1_011000001100;
      patterns[39106] = 29'b1_001100011000_010_0_011000110001;
      patterns[39107] = 29'b1_001100011000_011_0_110001100010;
      patterns[39108] = 29'b1_001100011000_100_0_100110001100;
      patterns[39109] = 29'b1_001100011000_101_0_010011000110;
      patterns[39110] = 29'b1_001100011000_110_1_001100011000;
      patterns[39111] = 29'b1_001100011000_111_1_001100011000;
      patterns[39112] = 29'b1_001100011001_000_1_001100011001;
      patterns[39113] = 29'b1_001100011001_001_1_011001001100;
      patterns[39114] = 29'b1_001100011001_010_0_011000110011;
      patterns[39115] = 29'b1_001100011001_011_0_110001100110;
      patterns[39116] = 29'b1_001100011001_100_1_100110001100;
      patterns[39117] = 29'b1_001100011001_101_0_110011000110;
      patterns[39118] = 29'b1_001100011001_110_1_001100011001;
      patterns[39119] = 29'b1_001100011001_111_1_001100011001;
      patterns[39120] = 29'b1_001100011010_000_1_001100011010;
      patterns[39121] = 29'b1_001100011010_001_1_011010001100;
      patterns[39122] = 29'b1_001100011010_010_0_011000110101;
      patterns[39123] = 29'b1_001100011010_011_0_110001101010;
      patterns[39124] = 29'b1_001100011010_100_0_100110001101;
      patterns[39125] = 29'b1_001100011010_101_1_010011000110;
      patterns[39126] = 29'b1_001100011010_110_1_001100011010;
      patterns[39127] = 29'b1_001100011010_111_1_001100011010;
      patterns[39128] = 29'b1_001100011011_000_1_001100011011;
      patterns[39129] = 29'b1_001100011011_001_1_011011001100;
      patterns[39130] = 29'b1_001100011011_010_0_011000110111;
      patterns[39131] = 29'b1_001100011011_011_0_110001101110;
      patterns[39132] = 29'b1_001100011011_100_1_100110001101;
      patterns[39133] = 29'b1_001100011011_101_1_110011000110;
      patterns[39134] = 29'b1_001100011011_110_1_001100011011;
      patterns[39135] = 29'b1_001100011011_111_1_001100011011;
      patterns[39136] = 29'b1_001100011100_000_1_001100011100;
      patterns[39137] = 29'b1_001100011100_001_1_011100001100;
      patterns[39138] = 29'b1_001100011100_010_0_011000111001;
      patterns[39139] = 29'b1_001100011100_011_0_110001110010;
      patterns[39140] = 29'b1_001100011100_100_0_100110001110;
      patterns[39141] = 29'b1_001100011100_101_0_010011000111;
      patterns[39142] = 29'b1_001100011100_110_1_001100011100;
      patterns[39143] = 29'b1_001100011100_111_1_001100011100;
      patterns[39144] = 29'b1_001100011101_000_1_001100011101;
      patterns[39145] = 29'b1_001100011101_001_1_011101001100;
      patterns[39146] = 29'b1_001100011101_010_0_011000111011;
      patterns[39147] = 29'b1_001100011101_011_0_110001110110;
      patterns[39148] = 29'b1_001100011101_100_1_100110001110;
      patterns[39149] = 29'b1_001100011101_101_0_110011000111;
      patterns[39150] = 29'b1_001100011101_110_1_001100011101;
      patterns[39151] = 29'b1_001100011101_111_1_001100011101;
      patterns[39152] = 29'b1_001100011110_000_1_001100011110;
      patterns[39153] = 29'b1_001100011110_001_1_011110001100;
      patterns[39154] = 29'b1_001100011110_010_0_011000111101;
      patterns[39155] = 29'b1_001100011110_011_0_110001111010;
      patterns[39156] = 29'b1_001100011110_100_0_100110001111;
      patterns[39157] = 29'b1_001100011110_101_1_010011000111;
      patterns[39158] = 29'b1_001100011110_110_1_001100011110;
      patterns[39159] = 29'b1_001100011110_111_1_001100011110;
      patterns[39160] = 29'b1_001100011111_000_1_001100011111;
      patterns[39161] = 29'b1_001100011111_001_1_011111001100;
      patterns[39162] = 29'b1_001100011111_010_0_011000111111;
      patterns[39163] = 29'b1_001100011111_011_0_110001111110;
      patterns[39164] = 29'b1_001100011111_100_1_100110001111;
      patterns[39165] = 29'b1_001100011111_101_1_110011000111;
      patterns[39166] = 29'b1_001100011111_110_1_001100011111;
      patterns[39167] = 29'b1_001100011111_111_1_001100011111;
      patterns[39168] = 29'b1_001100100000_000_1_001100100000;
      patterns[39169] = 29'b1_001100100000_001_1_100000001100;
      patterns[39170] = 29'b1_001100100000_010_0_011001000001;
      patterns[39171] = 29'b1_001100100000_011_0_110010000010;
      patterns[39172] = 29'b1_001100100000_100_0_100110010000;
      patterns[39173] = 29'b1_001100100000_101_0_010011001000;
      patterns[39174] = 29'b1_001100100000_110_1_001100100000;
      patterns[39175] = 29'b1_001100100000_111_1_001100100000;
      patterns[39176] = 29'b1_001100100001_000_1_001100100001;
      patterns[39177] = 29'b1_001100100001_001_1_100001001100;
      patterns[39178] = 29'b1_001100100001_010_0_011001000011;
      patterns[39179] = 29'b1_001100100001_011_0_110010000110;
      patterns[39180] = 29'b1_001100100001_100_1_100110010000;
      patterns[39181] = 29'b1_001100100001_101_0_110011001000;
      patterns[39182] = 29'b1_001100100001_110_1_001100100001;
      patterns[39183] = 29'b1_001100100001_111_1_001100100001;
      patterns[39184] = 29'b1_001100100010_000_1_001100100010;
      patterns[39185] = 29'b1_001100100010_001_1_100010001100;
      patterns[39186] = 29'b1_001100100010_010_0_011001000101;
      patterns[39187] = 29'b1_001100100010_011_0_110010001010;
      patterns[39188] = 29'b1_001100100010_100_0_100110010001;
      patterns[39189] = 29'b1_001100100010_101_1_010011001000;
      patterns[39190] = 29'b1_001100100010_110_1_001100100010;
      patterns[39191] = 29'b1_001100100010_111_1_001100100010;
      patterns[39192] = 29'b1_001100100011_000_1_001100100011;
      patterns[39193] = 29'b1_001100100011_001_1_100011001100;
      patterns[39194] = 29'b1_001100100011_010_0_011001000111;
      patterns[39195] = 29'b1_001100100011_011_0_110010001110;
      patterns[39196] = 29'b1_001100100011_100_1_100110010001;
      patterns[39197] = 29'b1_001100100011_101_1_110011001000;
      patterns[39198] = 29'b1_001100100011_110_1_001100100011;
      patterns[39199] = 29'b1_001100100011_111_1_001100100011;
      patterns[39200] = 29'b1_001100100100_000_1_001100100100;
      patterns[39201] = 29'b1_001100100100_001_1_100100001100;
      patterns[39202] = 29'b1_001100100100_010_0_011001001001;
      patterns[39203] = 29'b1_001100100100_011_0_110010010010;
      patterns[39204] = 29'b1_001100100100_100_0_100110010010;
      patterns[39205] = 29'b1_001100100100_101_0_010011001001;
      patterns[39206] = 29'b1_001100100100_110_1_001100100100;
      patterns[39207] = 29'b1_001100100100_111_1_001100100100;
      patterns[39208] = 29'b1_001100100101_000_1_001100100101;
      patterns[39209] = 29'b1_001100100101_001_1_100101001100;
      patterns[39210] = 29'b1_001100100101_010_0_011001001011;
      patterns[39211] = 29'b1_001100100101_011_0_110010010110;
      patterns[39212] = 29'b1_001100100101_100_1_100110010010;
      patterns[39213] = 29'b1_001100100101_101_0_110011001001;
      patterns[39214] = 29'b1_001100100101_110_1_001100100101;
      patterns[39215] = 29'b1_001100100101_111_1_001100100101;
      patterns[39216] = 29'b1_001100100110_000_1_001100100110;
      patterns[39217] = 29'b1_001100100110_001_1_100110001100;
      patterns[39218] = 29'b1_001100100110_010_0_011001001101;
      patterns[39219] = 29'b1_001100100110_011_0_110010011010;
      patterns[39220] = 29'b1_001100100110_100_0_100110010011;
      patterns[39221] = 29'b1_001100100110_101_1_010011001001;
      patterns[39222] = 29'b1_001100100110_110_1_001100100110;
      patterns[39223] = 29'b1_001100100110_111_1_001100100110;
      patterns[39224] = 29'b1_001100100111_000_1_001100100111;
      patterns[39225] = 29'b1_001100100111_001_1_100111001100;
      patterns[39226] = 29'b1_001100100111_010_0_011001001111;
      patterns[39227] = 29'b1_001100100111_011_0_110010011110;
      patterns[39228] = 29'b1_001100100111_100_1_100110010011;
      patterns[39229] = 29'b1_001100100111_101_1_110011001001;
      patterns[39230] = 29'b1_001100100111_110_1_001100100111;
      patterns[39231] = 29'b1_001100100111_111_1_001100100111;
      patterns[39232] = 29'b1_001100101000_000_1_001100101000;
      patterns[39233] = 29'b1_001100101000_001_1_101000001100;
      patterns[39234] = 29'b1_001100101000_010_0_011001010001;
      patterns[39235] = 29'b1_001100101000_011_0_110010100010;
      patterns[39236] = 29'b1_001100101000_100_0_100110010100;
      patterns[39237] = 29'b1_001100101000_101_0_010011001010;
      patterns[39238] = 29'b1_001100101000_110_1_001100101000;
      patterns[39239] = 29'b1_001100101000_111_1_001100101000;
      patterns[39240] = 29'b1_001100101001_000_1_001100101001;
      patterns[39241] = 29'b1_001100101001_001_1_101001001100;
      patterns[39242] = 29'b1_001100101001_010_0_011001010011;
      patterns[39243] = 29'b1_001100101001_011_0_110010100110;
      patterns[39244] = 29'b1_001100101001_100_1_100110010100;
      patterns[39245] = 29'b1_001100101001_101_0_110011001010;
      patterns[39246] = 29'b1_001100101001_110_1_001100101001;
      patterns[39247] = 29'b1_001100101001_111_1_001100101001;
      patterns[39248] = 29'b1_001100101010_000_1_001100101010;
      patterns[39249] = 29'b1_001100101010_001_1_101010001100;
      patterns[39250] = 29'b1_001100101010_010_0_011001010101;
      patterns[39251] = 29'b1_001100101010_011_0_110010101010;
      patterns[39252] = 29'b1_001100101010_100_0_100110010101;
      patterns[39253] = 29'b1_001100101010_101_1_010011001010;
      patterns[39254] = 29'b1_001100101010_110_1_001100101010;
      patterns[39255] = 29'b1_001100101010_111_1_001100101010;
      patterns[39256] = 29'b1_001100101011_000_1_001100101011;
      patterns[39257] = 29'b1_001100101011_001_1_101011001100;
      patterns[39258] = 29'b1_001100101011_010_0_011001010111;
      patterns[39259] = 29'b1_001100101011_011_0_110010101110;
      patterns[39260] = 29'b1_001100101011_100_1_100110010101;
      patterns[39261] = 29'b1_001100101011_101_1_110011001010;
      patterns[39262] = 29'b1_001100101011_110_1_001100101011;
      patterns[39263] = 29'b1_001100101011_111_1_001100101011;
      patterns[39264] = 29'b1_001100101100_000_1_001100101100;
      patterns[39265] = 29'b1_001100101100_001_1_101100001100;
      patterns[39266] = 29'b1_001100101100_010_0_011001011001;
      patterns[39267] = 29'b1_001100101100_011_0_110010110010;
      patterns[39268] = 29'b1_001100101100_100_0_100110010110;
      patterns[39269] = 29'b1_001100101100_101_0_010011001011;
      patterns[39270] = 29'b1_001100101100_110_1_001100101100;
      patterns[39271] = 29'b1_001100101100_111_1_001100101100;
      patterns[39272] = 29'b1_001100101101_000_1_001100101101;
      patterns[39273] = 29'b1_001100101101_001_1_101101001100;
      patterns[39274] = 29'b1_001100101101_010_0_011001011011;
      patterns[39275] = 29'b1_001100101101_011_0_110010110110;
      patterns[39276] = 29'b1_001100101101_100_1_100110010110;
      patterns[39277] = 29'b1_001100101101_101_0_110011001011;
      patterns[39278] = 29'b1_001100101101_110_1_001100101101;
      patterns[39279] = 29'b1_001100101101_111_1_001100101101;
      patterns[39280] = 29'b1_001100101110_000_1_001100101110;
      patterns[39281] = 29'b1_001100101110_001_1_101110001100;
      patterns[39282] = 29'b1_001100101110_010_0_011001011101;
      patterns[39283] = 29'b1_001100101110_011_0_110010111010;
      patterns[39284] = 29'b1_001100101110_100_0_100110010111;
      patterns[39285] = 29'b1_001100101110_101_1_010011001011;
      patterns[39286] = 29'b1_001100101110_110_1_001100101110;
      patterns[39287] = 29'b1_001100101110_111_1_001100101110;
      patterns[39288] = 29'b1_001100101111_000_1_001100101111;
      patterns[39289] = 29'b1_001100101111_001_1_101111001100;
      patterns[39290] = 29'b1_001100101111_010_0_011001011111;
      patterns[39291] = 29'b1_001100101111_011_0_110010111110;
      patterns[39292] = 29'b1_001100101111_100_1_100110010111;
      patterns[39293] = 29'b1_001100101111_101_1_110011001011;
      patterns[39294] = 29'b1_001100101111_110_1_001100101111;
      patterns[39295] = 29'b1_001100101111_111_1_001100101111;
      patterns[39296] = 29'b1_001100110000_000_1_001100110000;
      patterns[39297] = 29'b1_001100110000_001_1_110000001100;
      patterns[39298] = 29'b1_001100110000_010_0_011001100001;
      patterns[39299] = 29'b1_001100110000_011_0_110011000010;
      patterns[39300] = 29'b1_001100110000_100_0_100110011000;
      patterns[39301] = 29'b1_001100110000_101_0_010011001100;
      patterns[39302] = 29'b1_001100110000_110_1_001100110000;
      patterns[39303] = 29'b1_001100110000_111_1_001100110000;
      patterns[39304] = 29'b1_001100110001_000_1_001100110001;
      patterns[39305] = 29'b1_001100110001_001_1_110001001100;
      patterns[39306] = 29'b1_001100110001_010_0_011001100011;
      patterns[39307] = 29'b1_001100110001_011_0_110011000110;
      patterns[39308] = 29'b1_001100110001_100_1_100110011000;
      patterns[39309] = 29'b1_001100110001_101_0_110011001100;
      patterns[39310] = 29'b1_001100110001_110_1_001100110001;
      patterns[39311] = 29'b1_001100110001_111_1_001100110001;
      patterns[39312] = 29'b1_001100110010_000_1_001100110010;
      patterns[39313] = 29'b1_001100110010_001_1_110010001100;
      patterns[39314] = 29'b1_001100110010_010_0_011001100101;
      patterns[39315] = 29'b1_001100110010_011_0_110011001010;
      patterns[39316] = 29'b1_001100110010_100_0_100110011001;
      patterns[39317] = 29'b1_001100110010_101_1_010011001100;
      patterns[39318] = 29'b1_001100110010_110_1_001100110010;
      patterns[39319] = 29'b1_001100110010_111_1_001100110010;
      patterns[39320] = 29'b1_001100110011_000_1_001100110011;
      patterns[39321] = 29'b1_001100110011_001_1_110011001100;
      patterns[39322] = 29'b1_001100110011_010_0_011001100111;
      patterns[39323] = 29'b1_001100110011_011_0_110011001110;
      patterns[39324] = 29'b1_001100110011_100_1_100110011001;
      patterns[39325] = 29'b1_001100110011_101_1_110011001100;
      patterns[39326] = 29'b1_001100110011_110_1_001100110011;
      patterns[39327] = 29'b1_001100110011_111_1_001100110011;
      patterns[39328] = 29'b1_001100110100_000_1_001100110100;
      patterns[39329] = 29'b1_001100110100_001_1_110100001100;
      patterns[39330] = 29'b1_001100110100_010_0_011001101001;
      patterns[39331] = 29'b1_001100110100_011_0_110011010010;
      patterns[39332] = 29'b1_001100110100_100_0_100110011010;
      patterns[39333] = 29'b1_001100110100_101_0_010011001101;
      patterns[39334] = 29'b1_001100110100_110_1_001100110100;
      patterns[39335] = 29'b1_001100110100_111_1_001100110100;
      patterns[39336] = 29'b1_001100110101_000_1_001100110101;
      patterns[39337] = 29'b1_001100110101_001_1_110101001100;
      patterns[39338] = 29'b1_001100110101_010_0_011001101011;
      patterns[39339] = 29'b1_001100110101_011_0_110011010110;
      patterns[39340] = 29'b1_001100110101_100_1_100110011010;
      patterns[39341] = 29'b1_001100110101_101_0_110011001101;
      patterns[39342] = 29'b1_001100110101_110_1_001100110101;
      patterns[39343] = 29'b1_001100110101_111_1_001100110101;
      patterns[39344] = 29'b1_001100110110_000_1_001100110110;
      patterns[39345] = 29'b1_001100110110_001_1_110110001100;
      patterns[39346] = 29'b1_001100110110_010_0_011001101101;
      patterns[39347] = 29'b1_001100110110_011_0_110011011010;
      patterns[39348] = 29'b1_001100110110_100_0_100110011011;
      patterns[39349] = 29'b1_001100110110_101_1_010011001101;
      patterns[39350] = 29'b1_001100110110_110_1_001100110110;
      patterns[39351] = 29'b1_001100110110_111_1_001100110110;
      patterns[39352] = 29'b1_001100110111_000_1_001100110111;
      patterns[39353] = 29'b1_001100110111_001_1_110111001100;
      patterns[39354] = 29'b1_001100110111_010_0_011001101111;
      patterns[39355] = 29'b1_001100110111_011_0_110011011110;
      patterns[39356] = 29'b1_001100110111_100_1_100110011011;
      patterns[39357] = 29'b1_001100110111_101_1_110011001101;
      patterns[39358] = 29'b1_001100110111_110_1_001100110111;
      patterns[39359] = 29'b1_001100110111_111_1_001100110111;
      patterns[39360] = 29'b1_001100111000_000_1_001100111000;
      patterns[39361] = 29'b1_001100111000_001_1_111000001100;
      patterns[39362] = 29'b1_001100111000_010_0_011001110001;
      patterns[39363] = 29'b1_001100111000_011_0_110011100010;
      patterns[39364] = 29'b1_001100111000_100_0_100110011100;
      patterns[39365] = 29'b1_001100111000_101_0_010011001110;
      patterns[39366] = 29'b1_001100111000_110_1_001100111000;
      patterns[39367] = 29'b1_001100111000_111_1_001100111000;
      patterns[39368] = 29'b1_001100111001_000_1_001100111001;
      patterns[39369] = 29'b1_001100111001_001_1_111001001100;
      patterns[39370] = 29'b1_001100111001_010_0_011001110011;
      patterns[39371] = 29'b1_001100111001_011_0_110011100110;
      patterns[39372] = 29'b1_001100111001_100_1_100110011100;
      patterns[39373] = 29'b1_001100111001_101_0_110011001110;
      patterns[39374] = 29'b1_001100111001_110_1_001100111001;
      patterns[39375] = 29'b1_001100111001_111_1_001100111001;
      patterns[39376] = 29'b1_001100111010_000_1_001100111010;
      patterns[39377] = 29'b1_001100111010_001_1_111010001100;
      patterns[39378] = 29'b1_001100111010_010_0_011001110101;
      patterns[39379] = 29'b1_001100111010_011_0_110011101010;
      patterns[39380] = 29'b1_001100111010_100_0_100110011101;
      patterns[39381] = 29'b1_001100111010_101_1_010011001110;
      patterns[39382] = 29'b1_001100111010_110_1_001100111010;
      patterns[39383] = 29'b1_001100111010_111_1_001100111010;
      patterns[39384] = 29'b1_001100111011_000_1_001100111011;
      patterns[39385] = 29'b1_001100111011_001_1_111011001100;
      patterns[39386] = 29'b1_001100111011_010_0_011001110111;
      patterns[39387] = 29'b1_001100111011_011_0_110011101110;
      patterns[39388] = 29'b1_001100111011_100_1_100110011101;
      patterns[39389] = 29'b1_001100111011_101_1_110011001110;
      patterns[39390] = 29'b1_001100111011_110_1_001100111011;
      patterns[39391] = 29'b1_001100111011_111_1_001100111011;
      patterns[39392] = 29'b1_001100111100_000_1_001100111100;
      patterns[39393] = 29'b1_001100111100_001_1_111100001100;
      patterns[39394] = 29'b1_001100111100_010_0_011001111001;
      patterns[39395] = 29'b1_001100111100_011_0_110011110010;
      patterns[39396] = 29'b1_001100111100_100_0_100110011110;
      patterns[39397] = 29'b1_001100111100_101_0_010011001111;
      patterns[39398] = 29'b1_001100111100_110_1_001100111100;
      patterns[39399] = 29'b1_001100111100_111_1_001100111100;
      patterns[39400] = 29'b1_001100111101_000_1_001100111101;
      patterns[39401] = 29'b1_001100111101_001_1_111101001100;
      patterns[39402] = 29'b1_001100111101_010_0_011001111011;
      patterns[39403] = 29'b1_001100111101_011_0_110011110110;
      patterns[39404] = 29'b1_001100111101_100_1_100110011110;
      patterns[39405] = 29'b1_001100111101_101_0_110011001111;
      patterns[39406] = 29'b1_001100111101_110_1_001100111101;
      patterns[39407] = 29'b1_001100111101_111_1_001100111101;
      patterns[39408] = 29'b1_001100111110_000_1_001100111110;
      patterns[39409] = 29'b1_001100111110_001_1_111110001100;
      patterns[39410] = 29'b1_001100111110_010_0_011001111101;
      patterns[39411] = 29'b1_001100111110_011_0_110011111010;
      patterns[39412] = 29'b1_001100111110_100_0_100110011111;
      patterns[39413] = 29'b1_001100111110_101_1_010011001111;
      patterns[39414] = 29'b1_001100111110_110_1_001100111110;
      patterns[39415] = 29'b1_001100111110_111_1_001100111110;
      patterns[39416] = 29'b1_001100111111_000_1_001100111111;
      patterns[39417] = 29'b1_001100111111_001_1_111111001100;
      patterns[39418] = 29'b1_001100111111_010_0_011001111111;
      patterns[39419] = 29'b1_001100111111_011_0_110011111110;
      patterns[39420] = 29'b1_001100111111_100_1_100110011111;
      patterns[39421] = 29'b1_001100111111_101_1_110011001111;
      patterns[39422] = 29'b1_001100111111_110_1_001100111111;
      patterns[39423] = 29'b1_001100111111_111_1_001100111111;
      patterns[39424] = 29'b1_001101000000_000_1_001101000000;
      patterns[39425] = 29'b1_001101000000_001_1_000000001101;
      patterns[39426] = 29'b1_001101000000_010_0_011010000001;
      patterns[39427] = 29'b1_001101000000_011_0_110100000010;
      patterns[39428] = 29'b1_001101000000_100_0_100110100000;
      patterns[39429] = 29'b1_001101000000_101_0_010011010000;
      patterns[39430] = 29'b1_001101000000_110_1_001101000000;
      patterns[39431] = 29'b1_001101000000_111_1_001101000000;
      patterns[39432] = 29'b1_001101000001_000_1_001101000001;
      patterns[39433] = 29'b1_001101000001_001_1_000001001101;
      patterns[39434] = 29'b1_001101000001_010_0_011010000011;
      patterns[39435] = 29'b1_001101000001_011_0_110100000110;
      patterns[39436] = 29'b1_001101000001_100_1_100110100000;
      patterns[39437] = 29'b1_001101000001_101_0_110011010000;
      patterns[39438] = 29'b1_001101000001_110_1_001101000001;
      patterns[39439] = 29'b1_001101000001_111_1_001101000001;
      patterns[39440] = 29'b1_001101000010_000_1_001101000010;
      patterns[39441] = 29'b1_001101000010_001_1_000010001101;
      patterns[39442] = 29'b1_001101000010_010_0_011010000101;
      patterns[39443] = 29'b1_001101000010_011_0_110100001010;
      patterns[39444] = 29'b1_001101000010_100_0_100110100001;
      patterns[39445] = 29'b1_001101000010_101_1_010011010000;
      patterns[39446] = 29'b1_001101000010_110_1_001101000010;
      patterns[39447] = 29'b1_001101000010_111_1_001101000010;
      patterns[39448] = 29'b1_001101000011_000_1_001101000011;
      patterns[39449] = 29'b1_001101000011_001_1_000011001101;
      patterns[39450] = 29'b1_001101000011_010_0_011010000111;
      patterns[39451] = 29'b1_001101000011_011_0_110100001110;
      patterns[39452] = 29'b1_001101000011_100_1_100110100001;
      patterns[39453] = 29'b1_001101000011_101_1_110011010000;
      patterns[39454] = 29'b1_001101000011_110_1_001101000011;
      patterns[39455] = 29'b1_001101000011_111_1_001101000011;
      patterns[39456] = 29'b1_001101000100_000_1_001101000100;
      patterns[39457] = 29'b1_001101000100_001_1_000100001101;
      patterns[39458] = 29'b1_001101000100_010_0_011010001001;
      patterns[39459] = 29'b1_001101000100_011_0_110100010010;
      patterns[39460] = 29'b1_001101000100_100_0_100110100010;
      patterns[39461] = 29'b1_001101000100_101_0_010011010001;
      patterns[39462] = 29'b1_001101000100_110_1_001101000100;
      patterns[39463] = 29'b1_001101000100_111_1_001101000100;
      patterns[39464] = 29'b1_001101000101_000_1_001101000101;
      patterns[39465] = 29'b1_001101000101_001_1_000101001101;
      patterns[39466] = 29'b1_001101000101_010_0_011010001011;
      patterns[39467] = 29'b1_001101000101_011_0_110100010110;
      patterns[39468] = 29'b1_001101000101_100_1_100110100010;
      patterns[39469] = 29'b1_001101000101_101_0_110011010001;
      patterns[39470] = 29'b1_001101000101_110_1_001101000101;
      patterns[39471] = 29'b1_001101000101_111_1_001101000101;
      patterns[39472] = 29'b1_001101000110_000_1_001101000110;
      patterns[39473] = 29'b1_001101000110_001_1_000110001101;
      patterns[39474] = 29'b1_001101000110_010_0_011010001101;
      patterns[39475] = 29'b1_001101000110_011_0_110100011010;
      patterns[39476] = 29'b1_001101000110_100_0_100110100011;
      patterns[39477] = 29'b1_001101000110_101_1_010011010001;
      patterns[39478] = 29'b1_001101000110_110_1_001101000110;
      patterns[39479] = 29'b1_001101000110_111_1_001101000110;
      patterns[39480] = 29'b1_001101000111_000_1_001101000111;
      patterns[39481] = 29'b1_001101000111_001_1_000111001101;
      patterns[39482] = 29'b1_001101000111_010_0_011010001111;
      patterns[39483] = 29'b1_001101000111_011_0_110100011110;
      patterns[39484] = 29'b1_001101000111_100_1_100110100011;
      patterns[39485] = 29'b1_001101000111_101_1_110011010001;
      patterns[39486] = 29'b1_001101000111_110_1_001101000111;
      patterns[39487] = 29'b1_001101000111_111_1_001101000111;
      patterns[39488] = 29'b1_001101001000_000_1_001101001000;
      patterns[39489] = 29'b1_001101001000_001_1_001000001101;
      patterns[39490] = 29'b1_001101001000_010_0_011010010001;
      patterns[39491] = 29'b1_001101001000_011_0_110100100010;
      patterns[39492] = 29'b1_001101001000_100_0_100110100100;
      patterns[39493] = 29'b1_001101001000_101_0_010011010010;
      patterns[39494] = 29'b1_001101001000_110_1_001101001000;
      patterns[39495] = 29'b1_001101001000_111_1_001101001000;
      patterns[39496] = 29'b1_001101001001_000_1_001101001001;
      patterns[39497] = 29'b1_001101001001_001_1_001001001101;
      patterns[39498] = 29'b1_001101001001_010_0_011010010011;
      patterns[39499] = 29'b1_001101001001_011_0_110100100110;
      patterns[39500] = 29'b1_001101001001_100_1_100110100100;
      patterns[39501] = 29'b1_001101001001_101_0_110011010010;
      patterns[39502] = 29'b1_001101001001_110_1_001101001001;
      patterns[39503] = 29'b1_001101001001_111_1_001101001001;
      patterns[39504] = 29'b1_001101001010_000_1_001101001010;
      patterns[39505] = 29'b1_001101001010_001_1_001010001101;
      patterns[39506] = 29'b1_001101001010_010_0_011010010101;
      patterns[39507] = 29'b1_001101001010_011_0_110100101010;
      patterns[39508] = 29'b1_001101001010_100_0_100110100101;
      patterns[39509] = 29'b1_001101001010_101_1_010011010010;
      patterns[39510] = 29'b1_001101001010_110_1_001101001010;
      patterns[39511] = 29'b1_001101001010_111_1_001101001010;
      patterns[39512] = 29'b1_001101001011_000_1_001101001011;
      patterns[39513] = 29'b1_001101001011_001_1_001011001101;
      patterns[39514] = 29'b1_001101001011_010_0_011010010111;
      patterns[39515] = 29'b1_001101001011_011_0_110100101110;
      patterns[39516] = 29'b1_001101001011_100_1_100110100101;
      patterns[39517] = 29'b1_001101001011_101_1_110011010010;
      patterns[39518] = 29'b1_001101001011_110_1_001101001011;
      patterns[39519] = 29'b1_001101001011_111_1_001101001011;
      patterns[39520] = 29'b1_001101001100_000_1_001101001100;
      patterns[39521] = 29'b1_001101001100_001_1_001100001101;
      patterns[39522] = 29'b1_001101001100_010_0_011010011001;
      patterns[39523] = 29'b1_001101001100_011_0_110100110010;
      patterns[39524] = 29'b1_001101001100_100_0_100110100110;
      patterns[39525] = 29'b1_001101001100_101_0_010011010011;
      patterns[39526] = 29'b1_001101001100_110_1_001101001100;
      patterns[39527] = 29'b1_001101001100_111_1_001101001100;
      patterns[39528] = 29'b1_001101001101_000_1_001101001101;
      patterns[39529] = 29'b1_001101001101_001_1_001101001101;
      patterns[39530] = 29'b1_001101001101_010_0_011010011011;
      patterns[39531] = 29'b1_001101001101_011_0_110100110110;
      patterns[39532] = 29'b1_001101001101_100_1_100110100110;
      patterns[39533] = 29'b1_001101001101_101_0_110011010011;
      patterns[39534] = 29'b1_001101001101_110_1_001101001101;
      patterns[39535] = 29'b1_001101001101_111_1_001101001101;
      patterns[39536] = 29'b1_001101001110_000_1_001101001110;
      patterns[39537] = 29'b1_001101001110_001_1_001110001101;
      patterns[39538] = 29'b1_001101001110_010_0_011010011101;
      patterns[39539] = 29'b1_001101001110_011_0_110100111010;
      patterns[39540] = 29'b1_001101001110_100_0_100110100111;
      patterns[39541] = 29'b1_001101001110_101_1_010011010011;
      patterns[39542] = 29'b1_001101001110_110_1_001101001110;
      patterns[39543] = 29'b1_001101001110_111_1_001101001110;
      patterns[39544] = 29'b1_001101001111_000_1_001101001111;
      patterns[39545] = 29'b1_001101001111_001_1_001111001101;
      patterns[39546] = 29'b1_001101001111_010_0_011010011111;
      patterns[39547] = 29'b1_001101001111_011_0_110100111110;
      patterns[39548] = 29'b1_001101001111_100_1_100110100111;
      patterns[39549] = 29'b1_001101001111_101_1_110011010011;
      patterns[39550] = 29'b1_001101001111_110_1_001101001111;
      patterns[39551] = 29'b1_001101001111_111_1_001101001111;
      patterns[39552] = 29'b1_001101010000_000_1_001101010000;
      patterns[39553] = 29'b1_001101010000_001_1_010000001101;
      patterns[39554] = 29'b1_001101010000_010_0_011010100001;
      patterns[39555] = 29'b1_001101010000_011_0_110101000010;
      patterns[39556] = 29'b1_001101010000_100_0_100110101000;
      patterns[39557] = 29'b1_001101010000_101_0_010011010100;
      patterns[39558] = 29'b1_001101010000_110_1_001101010000;
      patterns[39559] = 29'b1_001101010000_111_1_001101010000;
      patterns[39560] = 29'b1_001101010001_000_1_001101010001;
      patterns[39561] = 29'b1_001101010001_001_1_010001001101;
      patterns[39562] = 29'b1_001101010001_010_0_011010100011;
      patterns[39563] = 29'b1_001101010001_011_0_110101000110;
      patterns[39564] = 29'b1_001101010001_100_1_100110101000;
      patterns[39565] = 29'b1_001101010001_101_0_110011010100;
      patterns[39566] = 29'b1_001101010001_110_1_001101010001;
      patterns[39567] = 29'b1_001101010001_111_1_001101010001;
      patterns[39568] = 29'b1_001101010010_000_1_001101010010;
      patterns[39569] = 29'b1_001101010010_001_1_010010001101;
      patterns[39570] = 29'b1_001101010010_010_0_011010100101;
      patterns[39571] = 29'b1_001101010010_011_0_110101001010;
      patterns[39572] = 29'b1_001101010010_100_0_100110101001;
      patterns[39573] = 29'b1_001101010010_101_1_010011010100;
      patterns[39574] = 29'b1_001101010010_110_1_001101010010;
      patterns[39575] = 29'b1_001101010010_111_1_001101010010;
      patterns[39576] = 29'b1_001101010011_000_1_001101010011;
      patterns[39577] = 29'b1_001101010011_001_1_010011001101;
      patterns[39578] = 29'b1_001101010011_010_0_011010100111;
      patterns[39579] = 29'b1_001101010011_011_0_110101001110;
      patterns[39580] = 29'b1_001101010011_100_1_100110101001;
      patterns[39581] = 29'b1_001101010011_101_1_110011010100;
      patterns[39582] = 29'b1_001101010011_110_1_001101010011;
      patterns[39583] = 29'b1_001101010011_111_1_001101010011;
      patterns[39584] = 29'b1_001101010100_000_1_001101010100;
      patterns[39585] = 29'b1_001101010100_001_1_010100001101;
      patterns[39586] = 29'b1_001101010100_010_0_011010101001;
      patterns[39587] = 29'b1_001101010100_011_0_110101010010;
      patterns[39588] = 29'b1_001101010100_100_0_100110101010;
      patterns[39589] = 29'b1_001101010100_101_0_010011010101;
      patterns[39590] = 29'b1_001101010100_110_1_001101010100;
      patterns[39591] = 29'b1_001101010100_111_1_001101010100;
      patterns[39592] = 29'b1_001101010101_000_1_001101010101;
      patterns[39593] = 29'b1_001101010101_001_1_010101001101;
      patterns[39594] = 29'b1_001101010101_010_0_011010101011;
      patterns[39595] = 29'b1_001101010101_011_0_110101010110;
      patterns[39596] = 29'b1_001101010101_100_1_100110101010;
      patterns[39597] = 29'b1_001101010101_101_0_110011010101;
      patterns[39598] = 29'b1_001101010101_110_1_001101010101;
      patterns[39599] = 29'b1_001101010101_111_1_001101010101;
      patterns[39600] = 29'b1_001101010110_000_1_001101010110;
      patterns[39601] = 29'b1_001101010110_001_1_010110001101;
      patterns[39602] = 29'b1_001101010110_010_0_011010101101;
      patterns[39603] = 29'b1_001101010110_011_0_110101011010;
      patterns[39604] = 29'b1_001101010110_100_0_100110101011;
      patterns[39605] = 29'b1_001101010110_101_1_010011010101;
      patterns[39606] = 29'b1_001101010110_110_1_001101010110;
      patterns[39607] = 29'b1_001101010110_111_1_001101010110;
      patterns[39608] = 29'b1_001101010111_000_1_001101010111;
      patterns[39609] = 29'b1_001101010111_001_1_010111001101;
      patterns[39610] = 29'b1_001101010111_010_0_011010101111;
      patterns[39611] = 29'b1_001101010111_011_0_110101011110;
      patterns[39612] = 29'b1_001101010111_100_1_100110101011;
      patterns[39613] = 29'b1_001101010111_101_1_110011010101;
      patterns[39614] = 29'b1_001101010111_110_1_001101010111;
      patterns[39615] = 29'b1_001101010111_111_1_001101010111;
      patterns[39616] = 29'b1_001101011000_000_1_001101011000;
      patterns[39617] = 29'b1_001101011000_001_1_011000001101;
      patterns[39618] = 29'b1_001101011000_010_0_011010110001;
      patterns[39619] = 29'b1_001101011000_011_0_110101100010;
      patterns[39620] = 29'b1_001101011000_100_0_100110101100;
      patterns[39621] = 29'b1_001101011000_101_0_010011010110;
      patterns[39622] = 29'b1_001101011000_110_1_001101011000;
      patterns[39623] = 29'b1_001101011000_111_1_001101011000;
      patterns[39624] = 29'b1_001101011001_000_1_001101011001;
      patterns[39625] = 29'b1_001101011001_001_1_011001001101;
      patterns[39626] = 29'b1_001101011001_010_0_011010110011;
      patterns[39627] = 29'b1_001101011001_011_0_110101100110;
      patterns[39628] = 29'b1_001101011001_100_1_100110101100;
      patterns[39629] = 29'b1_001101011001_101_0_110011010110;
      patterns[39630] = 29'b1_001101011001_110_1_001101011001;
      patterns[39631] = 29'b1_001101011001_111_1_001101011001;
      patterns[39632] = 29'b1_001101011010_000_1_001101011010;
      patterns[39633] = 29'b1_001101011010_001_1_011010001101;
      patterns[39634] = 29'b1_001101011010_010_0_011010110101;
      patterns[39635] = 29'b1_001101011010_011_0_110101101010;
      patterns[39636] = 29'b1_001101011010_100_0_100110101101;
      patterns[39637] = 29'b1_001101011010_101_1_010011010110;
      patterns[39638] = 29'b1_001101011010_110_1_001101011010;
      patterns[39639] = 29'b1_001101011010_111_1_001101011010;
      patterns[39640] = 29'b1_001101011011_000_1_001101011011;
      patterns[39641] = 29'b1_001101011011_001_1_011011001101;
      patterns[39642] = 29'b1_001101011011_010_0_011010110111;
      patterns[39643] = 29'b1_001101011011_011_0_110101101110;
      patterns[39644] = 29'b1_001101011011_100_1_100110101101;
      patterns[39645] = 29'b1_001101011011_101_1_110011010110;
      patterns[39646] = 29'b1_001101011011_110_1_001101011011;
      patterns[39647] = 29'b1_001101011011_111_1_001101011011;
      patterns[39648] = 29'b1_001101011100_000_1_001101011100;
      patterns[39649] = 29'b1_001101011100_001_1_011100001101;
      patterns[39650] = 29'b1_001101011100_010_0_011010111001;
      patterns[39651] = 29'b1_001101011100_011_0_110101110010;
      patterns[39652] = 29'b1_001101011100_100_0_100110101110;
      patterns[39653] = 29'b1_001101011100_101_0_010011010111;
      patterns[39654] = 29'b1_001101011100_110_1_001101011100;
      patterns[39655] = 29'b1_001101011100_111_1_001101011100;
      patterns[39656] = 29'b1_001101011101_000_1_001101011101;
      patterns[39657] = 29'b1_001101011101_001_1_011101001101;
      patterns[39658] = 29'b1_001101011101_010_0_011010111011;
      patterns[39659] = 29'b1_001101011101_011_0_110101110110;
      patterns[39660] = 29'b1_001101011101_100_1_100110101110;
      patterns[39661] = 29'b1_001101011101_101_0_110011010111;
      patterns[39662] = 29'b1_001101011101_110_1_001101011101;
      patterns[39663] = 29'b1_001101011101_111_1_001101011101;
      patterns[39664] = 29'b1_001101011110_000_1_001101011110;
      patterns[39665] = 29'b1_001101011110_001_1_011110001101;
      patterns[39666] = 29'b1_001101011110_010_0_011010111101;
      patterns[39667] = 29'b1_001101011110_011_0_110101111010;
      patterns[39668] = 29'b1_001101011110_100_0_100110101111;
      patterns[39669] = 29'b1_001101011110_101_1_010011010111;
      patterns[39670] = 29'b1_001101011110_110_1_001101011110;
      patterns[39671] = 29'b1_001101011110_111_1_001101011110;
      patterns[39672] = 29'b1_001101011111_000_1_001101011111;
      patterns[39673] = 29'b1_001101011111_001_1_011111001101;
      patterns[39674] = 29'b1_001101011111_010_0_011010111111;
      patterns[39675] = 29'b1_001101011111_011_0_110101111110;
      patterns[39676] = 29'b1_001101011111_100_1_100110101111;
      patterns[39677] = 29'b1_001101011111_101_1_110011010111;
      patterns[39678] = 29'b1_001101011111_110_1_001101011111;
      patterns[39679] = 29'b1_001101011111_111_1_001101011111;
      patterns[39680] = 29'b1_001101100000_000_1_001101100000;
      patterns[39681] = 29'b1_001101100000_001_1_100000001101;
      patterns[39682] = 29'b1_001101100000_010_0_011011000001;
      patterns[39683] = 29'b1_001101100000_011_0_110110000010;
      patterns[39684] = 29'b1_001101100000_100_0_100110110000;
      patterns[39685] = 29'b1_001101100000_101_0_010011011000;
      patterns[39686] = 29'b1_001101100000_110_1_001101100000;
      patterns[39687] = 29'b1_001101100000_111_1_001101100000;
      patterns[39688] = 29'b1_001101100001_000_1_001101100001;
      patterns[39689] = 29'b1_001101100001_001_1_100001001101;
      patterns[39690] = 29'b1_001101100001_010_0_011011000011;
      patterns[39691] = 29'b1_001101100001_011_0_110110000110;
      patterns[39692] = 29'b1_001101100001_100_1_100110110000;
      patterns[39693] = 29'b1_001101100001_101_0_110011011000;
      patterns[39694] = 29'b1_001101100001_110_1_001101100001;
      patterns[39695] = 29'b1_001101100001_111_1_001101100001;
      patterns[39696] = 29'b1_001101100010_000_1_001101100010;
      patterns[39697] = 29'b1_001101100010_001_1_100010001101;
      patterns[39698] = 29'b1_001101100010_010_0_011011000101;
      patterns[39699] = 29'b1_001101100010_011_0_110110001010;
      patterns[39700] = 29'b1_001101100010_100_0_100110110001;
      patterns[39701] = 29'b1_001101100010_101_1_010011011000;
      patterns[39702] = 29'b1_001101100010_110_1_001101100010;
      patterns[39703] = 29'b1_001101100010_111_1_001101100010;
      patterns[39704] = 29'b1_001101100011_000_1_001101100011;
      patterns[39705] = 29'b1_001101100011_001_1_100011001101;
      patterns[39706] = 29'b1_001101100011_010_0_011011000111;
      patterns[39707] = 29'b1_001101100011_011_0_110110001110;
      patterns[39708] = 29'b1_001101100011_100_1_100110110001;
      patterns[39709] = 29'b1_001101100011_101_1_110011011000;
      patterns[39710] = 29'b1_001101100011_110_1_001101100011;
      patterns[39711] = 29'b1_001101100011_111_1_001101100011;
      patterns[39712] = 29'b1_001101100100_000_1_001101100100;
      patterns[39713] = 29'b1_001101100100_001_1_100100001101;
      patterns[39714] = 29'b1_001101100100_010_0_011011001001;
      patterns[39715] = 29'b1_001101100100_011_0_110110010010;
      patterns[39716] = 29'b1_001101100100_100_0_100110110010;
      patterns[39717] = 29'b1_001101100100_101_0_010011011001;
      patterns[39718] = 29'b1_001101100100_110_1_001101100100;
      patterns[39719] = 29'b1_001101100100_111_1_001101100100;
      patterns[39720] = 29'b1_001101100101_000_1_001101100101;
      patterns[39721] = 29'b1_001101100101_001_1_100101001101;
      patterns[39722] = 29'b1_001101100101_010_0_011011001011;
      patterns[39723] = 29'b1_001101100101_011_0_110110010110;
      patterns[39724] = 29'b1_001101100101_100_1_100110110010;
      patterns[39725] = 29'b1_001101100101_101_0_110011011001;
      patterns[39726] = 29'b1_001101100101_110_1_001101100101;
      patterns[39727] = 29'b1_001101100101_111_1_001101100101;
      patterns[39728] = 29'b1_001101100110_000_1_001101100110;
      patterns[39729] = 29'b1_001101100110_001_1_100110001101;
      patterns[39730] = 29'b1_001101100110_010_0_011011001101;
      patterns[39731] = 29'b1_001101100110_011_0_110110011010;
      patterns[39732] = 29'b1_001101100110_100_0_100110110011;
      patterns[39733] = 29'b1_001101100110_101_1_010011011001;
      patterns[39734] = 29'b1_001101100110_110_1_001101100110;
      patterns[39735] = 29'b1_001101100110_111_1_001101100110;
      patterns[39736] = 29'b1_001101100111_000_1_001101100111;
      patterns[39737] = 29'b1_001101100111_001_1_100111001101;
      patterns[39738] = 29'b1_001101100111_010_0_011011001111;
      patterns[39739] = 29'b1_001101100111_011_0_110110011110;
      patterns[39740] = 29'b1_001101100111_100_1_100110110011;
      patterns[39741] = 29'b1_001101100111_101_1_110011011001;
      patterns[39742] = 29'b1_001101100111_110_1_001101100111;
      patterns[39743] = 29'b1_001101100111_111_1_001101100111;
      patterns[39744] = 29'b1_001101101000_000_1_001101101000;
      patterns[39745] = 29'b1_001101101000_001_1_101000001101;
      patterns[39746] = 29'b1_001101101000_010_0_011011010001;
      patterns[39747] = 29'b1_001101101000_011_0_110110100010;
      patterns[39748] = 29'b1_001101101000_100_0_100110110100;
      patterns[39749] = 29'b1_001101101000_101_0_010011011010;
      patterns[39750] = 29'b1_001101101000_110_1_001101101000;
      patterns[39751] = 29'b1_001101101000_111_1_001101101000;
      patterns[39752] = 29'b1_001101101001_000_1_001101101001;
      patterns[39753] = 29'b1_001101101001_001_1_101001001101;
      patterns[39754] = 29'b1_001101101001_010_0_011011010011;
      patterns[39755] = 29'b1_001101101001_011_0_110110100110;
      patterns[39756] = 29'b1_001101101001_100_1_100110110100;
      patterns[39757] = 29'b1_001101101001_101_0_110011011010;
      patterns[39758] = 29'b1_001101101001_110_1_001101101001;
      patterns[39759] = 29'b1_001101101001_111_1_001101101001;
      patterns[39760] = 29'b1_001101101010_000_1_001101101010;
      patterns[39761] = 29'b1_001101101010_001_1_101010001101;
      patterns[39762] = 29'b1_001101101010_010_0_011011010101;
      patterns[39763] = 29'b1_001101101010_011_0_110110101010;
      patterns[39764] = 29'b1_001101101010_100_0_100110110101;
      patterns[39765] = 29'b1_001101101010_101_1_010011011010;
      patterns[39766] = 29'b1_001101101010_110_1_001101101010;
      patterns[39767] = 29'b1_001101101010_111_1_001101101010;
      patterns[39768] = 29'b1_001101101011_000_1_001101101011;
      patterns[39769] = 29'b1_001101101011_001_1_101011001101;
      patterns[39770] = 29'b1_001101101011_010_0_011011010111;
      patterns[39771] = 29'b1_001101101011_011_0_110110101110;
      patterns[39772] = 29'b1_001101101011_100_1_100110110101;
      patterns[39773] = 29'b1_001101101011_101_1_110011011010;
      patterns[39774] = 29'b1_001101101011_110_1_001101101011;
      patterns[39775] = 29'b1_001101101011_111_1_001101101011;
      patterns[39776] = 29'b1_001101101100_000_1_001101101100;
      patterns[39777] = 29'b1_001101101100_001_1_101100001101;
      patterns[39778] = 29'b1_001101101100_010_0_011011011001;
      patterns[39779] = 29'b1_001101101100_011_0_110110110010;
      patterns[39780] = 29'b1_001101101100_100_0_100110110110;
      patterns[39781] = 29'b1_001101101100_101_0_010011011011;
      patterns[39782] = 29'b1_001101101100_110_1_001101101100;
      patterns[39783] = 29'b1_001101101100_111_1_001101101100;
      patterns[39784] = 29'b1_001101101101_000_1_001101101101;
      patterns[39785] = 29'b1_001101101101_001_1_101101001101;
      patterns[39786] = 29'b1_001101101101_010_0_011011011011;
      patterns[39787] = 29'b1_001101101101_011_0_110110110110;
      patterns[39788] = 29'b1_001101101101_100_1_100110110110;
      patterns[39789] = 29'b1_001101101101_101_0_110011011011;
      patterns[39790] = 29'b1_001101101101_110_1_001101101101;
      patterns[39791] = 29'b1_001101101101_111_1_001101101101;
      patterns[39792] = 29'b1_001101101110_000_1_001101101110;
      patterns[39793] = 29'b1_001101101110_001_1_101110001101;
      patterns[39794] = 29'b1_001101101110_010_0_011011011101;
      patterns[39795] = 29'b1_001101101110_011_0_110110111010;
      patterns[39796] = 29'b1_001101101110_100_0_100110110111;
      patterns[39797] = 29'b1_001101101110_101_1_010011011011;
      patterns[39798] = 29'b1_001101101110_110_1_001101101110;
      patterns[39799] = 29'b1_001101101110_111_1_001101101110;
      patterns[39800] = 29'b1_001101101111_000_1_001101101111;
      patterns[39801] = 29'b1_001101101111_001_1_101111001101;
      patterns[39802] = 29'b1_001101101111_010_0_011011011111;
      patterns[39803] = 29'b1_001101101111_011_0_110110111110;
      patterns[39804] = 29'b1_001101101111_100_1_100110110111;
      patterns[39805] = 29'b1_001101101111_101_1_110011011011;
      patterns[39806] = 29'b1_001101101111_110_1_001101101111;
      patterns[39807] = 29'b1_001101101111_111_1_001101101111;
      patterns[39808] = 29'b1_001101110000_000_1_001101110000;
      patterns[39809] = 29'b1_001101110000_001_1_110000001101;
      patterns[39810] = 29'b1_001101110000_010_0_011011100001;
      patterns[39811] = 29'b1_001101110000_011_0_110111000010;
      patterns[39812] = 29'b1_001101110000_100_0_100110111000;
      patterns[39813] = 29'b1_001101110000_101_0_010011011100;
      patterns[39814] = 29'b1_001101110000_110_1_001101110000;
      patterns[39815] = 29'b1_001101110000_111_1_001101110000;
      patterns[39816] = 29'b1_001101110001_000_1_001101110001;
      patterns[39817] = 29'b1_001101110001_001_1_110001001101;
      patterns[39818] = 29'b1_001101110001_010_0_011011100011;
      patterns[39819] = 29'b1_001101110001_011_0_110111000110;
      patterns[39820] = 29'b1_001101110001_100_1_100110111000;
      patterns[39821] = 29'b1_001101110001_101_0_110011011100;
      patterns[39822] = 29'b1_001101110001_110_1_001101110001;
      patterns[39823] = 29'b1_001101110001_111_1_001101110001;
      patterns[39824] = 29'b1_001101110010_000_1_001101110010;
      patterns[39825] = 29'b1_001101110010_001_1_110010001101;
      patterns[39826] = 29'b1_001101110010_010_0_011011100101;
      patterns[39827] = 29'b1_001101110010_011_0_110111001010;
      patterns[39828] = 29'b1_001101110010_100_0_100110111001;
      patterns[39829] = 29'b1_001101110010_101_1_010011011100;
      patterns[39830] = 29'b1_001101110010_110_1_001101110010;
      patterns[39831] = 29'b1_001101110010_111_1_001101110010;
      patterns[39832] = 29'b1_001101110011_000_1_001101110011;
      patterns[39833] = 29'b1_001101110011_001_1_110011001101;
      patterns[39834] = 29'b1_001101110011_010_0_011011100111;
      patterns[39835] = 29'b1_001101110011_011_0_110111001110;
      patterns[39836] = 29'b1_001101110011_100_1_100110111001;
      patterns[39837] = 29'b1_001101110011_101_1_110011011100;
      patterns[39838] = 29'b1_001101110011_110_1_001101110011;
      patterns[39839] = 29'b1_001101110011_111_1_001101110011;
      patterns[39840] = 29'b1_001101110100_000_1_001101110100;
      patterns[39841] = 29'b1_001101110100_001_1_110100001101;
      patterns[39842] = 29'b1_001101110100_010_0_011011101001;
      patterns[39843] = 29'b1_001101110100_011_0_110111010010;
      patterns[39844] = 29'b1_001101110100_100_0_100110111010;
      patterns[39845] = 29'b1_001101110100_101_0_010011011101;
      patterns[39846] = 29'b1_001101110100_110_1_001101110100;
      patterns[39847] = 29'b1_001101110100_111_1_001101110100;
      patterns[39848] = 29'b1_001101110101_000_1_001101110101;
      patterns[39849] = 29'b1_001101110101_001_1_110101001101;
      patterns[39850] = 29'b1_001101110101_010_0_011011101011;
      patterns[39851] = 29'b1_001101110101_011_0_110111010110;
      patterns[39852] = 29'b1_001101110101_100_1_100110111010;
      patterns[39853] = 29'b1_001101110101_101_0_110011011101;
      patterns[39854] = 29'b1_001101110101_110_1_001101110101;
      patterns[39855] = 29'b1_001101110101_111_1_001101110101;
      patterns[39856] = 29'b1_001101110110_000_1_001101110110;
      patterns[39857] = 29'b1_001101110110_001_1_110110001101;
      patterns[39858] = 29'b1_001101110110_010_0_011011101101;
      patterns[39859] = 29'b1_001101110110_011_0_110111011010;
      patterns[39860] = 29'b1_001101110110_100_0_100110111011;
      patterns[39861] = 29'b1_001101110110_101_1_010011011101;
      patterns[39862] = 29'b1_001101110110_110_1_001101110110;
      patterns[39863] = 29'b1_001101110110_111_1_001101110110;
      patterns[39864] = 29'b1_001101110111_000_1_001101110111;
      patterns[39865] = 29'b1_001101110111_001_1_110111001101;
      patterns[39866] = 29'b1_001101110111_010_0_011011101111;
      patterns[39867] = 29'b1_001101110111_011_0_110111011110;
      patterns[39868] = 29'b1_001101110111_100_1_100110111011;
      patterns[39869] = 29'b1_001101110111_101_1_110011011101;
      patterns[39870] = 29'b1_001101110111_110_1_001101110111;
      patterns[39871] = 29'b1_001101110111_111_1_001101110111;
      patterns[39872] = 29'b1_001101111000_000_1_001101111000;
      patterns[39873] = 29'b1_001101111000_001_1_111000001101;
      patterns[39874] = 29'b1_001101111000_010_0_011011110001;
      patterns[39875] = 29'b1_001101111000_011_0_110111100010;
      patterns[39876] = 29'b1_001101111000_100_0_100110111100;
      patterns[39877] = 29'b1_001101111000_101_0_010011011110;
      patterns[39878] = 29'b1_001101111000_110_1_001101111000;
      patterns[39879] = 29'b1_001101111000_111_1_001101111000;
      patterns[39880] = 29'b1_001101111001_000_1_001101111001;
      patterns[39881] = 29'b1_001101111001_001_1_111001001101;
      patterns[39882] = 29'b1_001101111001_010_0_011011110011;
      patterns[39883] = 29'b1_001101111001_011_0_110111100110;
      patterns[39884] = 29'b1_001101111001_100_1_100110111100;
      patterns[39885] = 29'b1_001101111001_101_0_110011011110;
      patterns[39886] = 29'b1_001101111001_110_1_001101111001;
      patterns[39887] = 29'b1_001101111001_111_1_001101111001;
      patterns[39888] = 29'b1_001101111010_000_1_001101111010;
      patterns[39889] = 29'b1_001101111010_001_1_111010001101;
      patterns[39890] = 29'b1_001101111010_010_0_011011110101;
      patterns[39891] = 29'b1_001101111010_011_0_110111101010;
      patterns[39892] = 29'b1_001101111010_100_0_100110111101;
      patterns[39893] = 29'b1_001101111010_101_1_010011011110;
      patterns[39894] = 29'b1_001101111010_110_1_001101111010;
      patterns[39895] = 29'b1_001101111010_111_1_001101111010;
      patterns[39896] = 29'b1_001101111011_000_1_001101111011;
      patterns[39897] = 29'b1_001101111011_001_1_111011001101;
      patterns[39898] = 29'b1_001101111011_010_0_011011110111;
      patterns[39899] = 29'b1_001101111011_011_0_110111101110;
      patterns[39900] = 29'b1_001101111011_100_1_100110111101;
      patterns[39901] = 29'b1_001101111011_101_1_110011011110;
      patterns[39902] = 29'b1_001101111011_110_1_001101111011;
      patterns[39903] = 29'b1_001101111011_111_1_001101111011;
      patterns[39904] = 29'b1_001101111100_000_1_001101111100;
      patterns[39905] = 29'b1_001101111100_001_1_111100001101;
      patterns[39906] = 29'b1_001101111100_010_0_011011111001;
      patterns[39907] = 29'b1_001101111100_011_0_110111110010;
      patterns[39908] = 29'b1_001101111100_100_0_100110111110;
      patterns[39909] = 29'b1_001101111100_101_0_010011011111;
      patterns[39910] = 29'b1_001101111100_110_1_001101111100;
      patterns[39911] = 29'b1_001101111100_111_1_001101111100;
      patterns[39912] = 29'b1_001101111101_000_1_001101111101;
      patterns[39913] = 29'b1_001101111101_001_1_111101001101;
      patterns[39914] = 29'b1_001101111101_010_0_011011111011;
      patterns[39915] = 29'b1_001101111101_011_0_110111110110;
      patterns[39916] = 29'b1_001101111101_100_1_100110111110;
      patterns[39917] = 29'b1_001101111101_101_0_110011011111;
      patterns[39918] = 29'b1_001101111101_110_1_001101111101;
      patterns[39919] = 29'b1_001101111101_111_1_001101111101;
      patterns[39920] = 29'b1_001101111110_000_1_001101111110;
      patterns[39921] = 29'b1_001101111110_001_1_111110001101;
      patterns[39922] = 29'b1_001101111110_010_0_011011111101;
      patterns[39923] = 29'b1_001101111110_011_0_110111111010;
      patterns[39924] = 29'b1_001101111110_100_0_100110111111;
      patterns[39925] = 29'b1_001101111110_101_1_010011011111;
      patterns[39926] = 29'b1_001101111110_110_1_001101111110;
      patterns[39927] = 29'b1_001101111110_111_1_001101111110;
      patterns[39928] = 29'b1_001101111111_000_1_001101111111;
      patterns[39929] = 29'b1_001101111111_001_1_111111001101;
      patterns[39930] = 29'b1_001101111111_010_0_011011111111;
      patterns[39931] = 29'b1_001101111111_011_0_110111111110;
      patterns[39932] = 29'b1_001101111111_100_1_100110111111;
      patterns[39933] = 29'b1_001101111111_101_1_110011011111;
      patterns[39934] = 29'b1_001101111111_110_1_001101111111;
      patterns[39935] = 29'b1_001101111111_111_1_001101111111;
      patterns[39936] = 29'b1_001110000000_000_1_001110000000;
      patterns[39937] = 29'b1_001110000000_001_1_000000001110;
      patterns[39938] = 29'b1_001110000000_010_0_011100000001;
      patterns[39939] = 29'b1_001110000000_011_0_111000000010;
      patterns[39940] = 29'b1_001110000000_100_0_100111000000;
      patterns[39941] = 29'b1_001110000000_101_0_010011100000;
      patterns[39942] = 29'b1_001110000000_110_1_001110000000;
      patterns[39943] = 29'b1_001110000000_111_1_001110000000;
      patterns[39944] = 29'b1_001110000001_000_1_001110000001;
      patterns[39945] = 29'b1_001110000001_001_1_000001001110;
      patterns[39946] = 29'b1_001110000001_010_0_011100000011;
      patterns[39947] = 29'b1_001110000001_011_0_111000000110;
      patterns[39948] = 29'b1_001110000001_100_1_100111000000;
      patterns[39949] = 29'b1_001110000001_101_0_110011100000;
      patterns[39950] = 29'b1_001110000001_110_1_001110000001;
      patterns[39951] = 29'b1_001110000001_111_1_001110000001;
      patterns[39952] = 29'b1_001110000010_000_1_001110000010;
      patterns[39953] = 29'b1_001110000010_001_1_000010001110;
      patterns[39954] = 29'b1_001110000010_010_0_011100000101;
      patterns[39955] = 29'b1_001110000010_011_0_111000001010;
      patterns[39956] = 29'b1_001110000010_100_0_100111000001;
      patterns[39957] = 29'b1_001110000010_101_1_010011100000;
      patterns[39958] = 29'b1_001110000010_110_1_001110000010;
      patterns[39959] = 29'b1_001110000010_111_1_001110000010;
      patterns[39960] = 29'b1_001110000011_000_1_001110000011;
      patterns[39961] = 29'b1_001110000011_001_1_000011001110;
      patterns[39962] = 29'b1_001110000011_010_0_011100000111;
      patterns[39963] = 29'b1_001110000011_011_0_111000001110;
      patterns[39964] = 29'b1_001110000011_100_1_100111000001;
      patterns[39965] = 29'b1_001110000011_101_1_110011100000;
      patterns[39966] = 29'b1_001110000011_110_1_001110000011;
      patterns[39967] = 29'b1_001110000011_111_1_001110000011;
      patterns[39968] = 29'b1_001110000100_000_1_001110000100;
      patterns[39969] = 29'b1_001110000100_001_1_000100001110;
      patterns[39970] = 29'b1_001110000100_010_0_011100001001;
      patterns[39971] = 29'b1_001110000100_011_0_111000010010;
      patterns[39972] = 29'b1_001110000100_100_0_100111000010;
      patterns[39973] = 29'b1_001110000100_101_0_010011100001;
      patterns[39974] = 29'b1_001110000100_110_1_001110000100;
      patterns[39975] = 29'b1_001110000100_111_1_001110000100;
      patterns[39976] = 29'b1_001110000101_000_1_001110000101;
      patterns[39977] = 29'b1_001110000101_001_1_000101001110;
      patterns[39978] = 29'b1_001110000101_010_0_011100001011;
      patterns[39979] = 29'b1_001110000101_011_0_111000010110;
      patterns[39980] = 29'b1_001110000101_100_1_100111000010;
      patterns[39981] = 29'b1_001110000101_101_0_110011100001;
      patterns[39982] = 29'b1_001110000101_110_1_001110000101;
      patterns[39983] = 29'b1_001110000101_111_1_001110000101;
      patterns[39984] = 29'b1_001110000110_000_1_001110000110;
      patterns[39985] = 29'b1_001110000110_001_1_000110001110;
      patterns[39986] = 29'b1_001110000110_010_0_011100001101;
      patterns[39987] = 29'b1_001110000110_011_0_111000011010;
      patterns[39988] = 29'b1_001110000110_100_0_100111000011;
      patterns[39989] = 29'b1_001110000110_101_1_010011100001;
      patterns[39990] = 29'b1_001110000110_110_1_001110000110;
      patterns[39991] = 29'b1_001110000110_111_1_001110000110;
      patterns[39992] = 29'b1_001110000111_000_1_001110000111;
      patterns[39993] = 29'b1_001110000111_001_1_000111001110;
      patterns[39994] = 29'b1_001110000111_010_0_011100001111;
      patterns[39995] = 29'b1_001110000111_011_0_111000011110;
      patterns[39996] = 29'b1_001110000111_100_1_100111000011;
      patterns[39997] = 29'b1_001110000111_101_1_110011100001;
      patterns[39998] = 29'b1_001110000111_110_1_001110000111;
      patterns[39999] = 29'b1_001110000111_111_1_001110000111;
      patterns[40000] = 29'b1_001110001000_000_1_001110001000;
      patterns[40001] = 29'b1_001110001000_001_1_001000001110;
      patterns[40002] = 29'b1_001110001000_010_0_011100010001;
      patterns[40003] = 29'b1_001110001000_011_0_111000100010;
      patterns[40004] = 29'b1_001110001000_100_0_100111000100;
      patterns[40005] = 29'b1_001110001000_101_0_010011100010;
      patterns[40006] = 29'b1_001110001000_110_1_001110001000;
      patterns[40007] = 29'b1_001110001000_111_1_001110001000;
      patterns[40008] = 29'b1_001110001001_000_1_001110001001;
      patterns[40009] = 29'b1_001110001001_001_1_001001001110;
      patterns[40010] = 29'b1_001110001001_010_0_011100010011;
      patterns[40011] = 29'b1_001110001001_011_0_111000100110;
      patterns[40012] = 29'b1_001110001001_100_1_100111000100;
      patterns[40013] = 29'b1_001110001001_101_0_110011100010;
      patterns[40014] = 29'b1_001110001001_110_1_001110001001;
      patterns[40015] = 29'b1_001110001001_111_1_001110001001;
      patterns[40016] = 29'b1_001110001010_000_1_001110001010;
      patterns[40017] = 29'b1_001110001010_001_1_001010001110;
      patterns[40018] = 29'b1_001110001010_010_0_011100010101;
      patterns[40019] = 29'b1_001110001010_011_0_111000101010;
      patterns[40020] = 29'b1_001110001010_100_0_100111000101;
      patterns[40021] = 29'b1_001110001010_101_1_010011100010;
      patterns[40022] = 29'b1_001110001010_110_1_001110001010;
      patterns[40023] = 29'b1_001110001010_111_1_001110001010;
      patterns[40024] = 29'b1_001110001011_000_1_001110001011;
      patterns[40025] = 29'b1_001110001011_001_1_001011001110;
      patterns[40026] = 29'b1_001110001011_010_0_011100010111;
      patterns[40027] = 29'b1_001110001011_011_0_111000101110;
      patterns[40028] = 29'b1_001110001011_100_1_100111000101;
      patterns[40029] = 29'b1_001110001011_101_1_110011100010;
      patterns[40030] = 29'b1_001110001011_110_1_001110001011;
      patterns[40031] = 29'b1_001110001011_111_1_001110001011;
      patterns[40032] = 29'b1_001110001100_000_1_001110001100;
      patterns[40033] = 29'b1_001110001100_001_1_001100001110;
      patterns[40034] = 29'b1_001110001100_010_0_011100011001;
      patterns[40035] = 29'b1_001110001100_011_0_111000110010;
      patterns[40036] = 29'b1_001110001100_100_0_100111000110;
      patterns[40037] = 29'b1_001110001100_101_0_010011100011;
      patterns[40038] = 29'b1_001110001100_110_1_001110001100;
      patterns[40039] = 29'b1_001110001100_111_1_001110001100;
      patterns[40040] = 29'b1_001110001101_000_1_001110001101;
      patterns[40041] = 29'b1_001110001101_001_1_001101001110;
      patterns[40042] = 29'b1_001110001101_010_0_011100011011;
      patterns[40043] = 29'b1_001110001101_011_0_111000110110;
      patterns[40044] = 29'b1_001110001101_100_1_100111000110;
      patterns[40045] = 29'b1_001110001101_101_0_110011100011;
      patterns[40046] = 29'b1_001110001101_110_1_001110001101;
      patterns[40047] = 29'b1_001110001101_111_1_001110001101;
      patterns[40048] = 29'b1_001110001110_000_1_001110001110;
      patterns[40049] = 29'b1_001110001110_001_1_001110001110;
      patterns[40050] = 29'b1_001110001110_010_0_011100011101;
      patterns[40051] = 29'b1_001110001110_011_0_111000111010;
      patterns[40052] = 29'b1_001110001110_100_0_100111000111;
      patterns[40053] = 29'b1_001110001110_101_1_010011100011;
      patterns[40054] = 29'b1_001110001110_110_1_001110001110;
      patterns[40055] = 29'b1_001110001110_111_1_001110001110;
      patterns[40056] = 29'b1_001110001111_000_1_001110001111;
      patterns[40057] = 29'b1_001110001111_001_1_001111001110;
      patterns[40058] = 29'b1_001110001111_010_0_011100011111;
      patterns[40059] = 29'b1_001110001111_011_0_111000111110;
      patterns[40060] = 29'b1_001110001111_100_1_100111000111;
      patterns[40061] = 29'b1_001110001111_101_1_110011100011;
      patterns[40062] = 29'b1_001110001111_110_1_001110001111;
      patterns[40063] = 29'b1_001110001111_111_1_001110001111;
      patterns[40064] = 29'b1_001110010000_000_1_001110010000;
      patterns[40065] = 29'b1_001110010000_001_1_010000001110;
      patterns[40066] = 29'b1_001110010000_010_0_011100100001;
      patterns[40067] = 29'b1_001110010000_011_0_111001000010;
      patterns[40068] = 29'b1_001110010000_100_0_100111001000;
      patterns[40069] = 29'b1_001110010000_101_0_010011100100;
      patterns[40070] = 29'b1_001110010000_110_1_001110010000;
      patterns[40071] = 29'b1_001110010000_111_1_001110010000;
      patterns[40072] = 29'b1_001110010001_000_1_001110010001;
      patterns[40073] = 29'b1_001110010001_001_1_010001001110;
      patterns[40074] = 29'b1_001110010001_010_0_011100100011;
      patterns[40075] = 29'b1_001110010001_011_0_111001000110;
      patterns[40076] = 29'b1_001110010001_100_1_100111001000;
      patterns[40077] = 29'b1_001110010001_101_0_110011100100;
      patterns[40078] = 29'b1_001110010001_110_1_001110010001;
      patterns[40079] = 29'b1_001110010001_111_1_001110010001;
      patterns[40080] = 29'b1_001110010010_000_1_001110010010;
      patterns[40081] = 29'b1_001110010010_001_1_010010001110;
      patterns[40082] = 29'b1_001110010010_010_0_011100100101;
      patterns[40083] = 29'b1_001110010010_011_0_111001001010;
      patterns[40084] = 29'b1_001110010010_100_0_100111001001;
      patterns[40085] = 29'b1_001110010010_101_1_010011100100;
      patterns[40086] = 29'b1_001110010010_110_1_001110010010;
      patterns[40087] = 29'b1_001110010010_111_1_001110010010;
      patterns[40088] = 29'b1_001110010011_000_1_001110010011;
      patterns[40089] = 29'b1_001110010011_001_1_010011001110;
      patterns[40090] = 29'b1_001110010011_010_0_011100100111;
      patterns[40091] = 29'b1_001110010011_011_0_111001001110;
      patterns[40092] = 29'b1_001110010011_100_1_100111001001;
      patterns[40093] = 29'b1_001110010011_101_1_110011100100;
      patterns[40094] = 29'b1_001110010011_110_1_001110010011;
      patterns[40095] = 29'b1_001110010011_111_1_001110010011;
      patterns[40096] = 29'b1_001110010100_000_1_001110010100;
      patterns[40097] = 29'b1_001110010100_001_1_010100001110;
      patterns[40098] = 29'b1_001110010100_010_0_011100101001;
      patterns[40099] = 29'b1_001110010100_011_0_111001010010;
      patterns[40100] = 29'b1_001110010100_100_0_100111001010;
      patterns[40101] = 29'b1_001110010100_101_0_010011100101;
      patterns[40102] = 29'b1_001110010100_110_1_001110010100;
      patterns[40103] = 29'b1_001110010100_111_1_001110010100;
      patterns[40104] = 29'b1_001110010101_000_1_001110010101;
      patterns[40105] = 29'b1_001110010101_001_1_010101001110;
      patterns[40106] = 29'b1_001110010101_010_0_011100101011;
      patterns[40107] = 29'b1_001110010101_011_0_111001010110;
      patterns[40108] = 29'b1_001110010101_100_1_100111001010;
      patterns[40109] = 29'b1_001110010101_101_0_110011100101;
      patterns[40110] = 29'b1_001110010101_110_1_001110010101;
      patterns[40111] = 29'b1_001110010101_111_1_001110010101;
      patterns[40112] = 29'b1_001110010110_000_1_001110010110;
      patterns[40113] = 29'b1_001110010110_001_1_010110001110;
      patterns[40114] = 29'b1_001110010110_010_0_011100101101;
      patterns[40115] = 29'b1_001110010110_011_0_111001011010;
      patterns[40116] = 29'b1_001110010110_100_0_100111001011;
      patterns[40117] = 29'b1_001110010110_101_1_010011100101;
      patterns[40118] = 29'b1_001110010110_110_1_001110010110;
      patterns[40119] = 29'b1_001110010110_111_1_001110010110;
      patterns[40120] = 29'b1_001110010111_000_1_001110010111;
      patterns[40121] = 29'b1_001110010111_001_1_010111001110;
      patterns[40122] = 29'b1_001110010111_010_0_011100101111;
      patterns[40123] = 29'b1_001110010111_011_0_111001011110;
      patterns[40124] = 29'b1_001110010111_100_1_100111001011;
      patterns[40125] = 29'b1_001110010111_101_1_110011100101;
      patterns[40126] = 29'b1_001110010111_110_1_001110010111;
      patterns[40127] = 29'b1_001110010111_111_1_001110010111;
      patterns[40128] = 29'b1_001110011000_000_1_001110011000;
      patterns[40129] = 29'b1_001110011000_001_1_011000001110;
      patterns[40130] = 29'b1_001110011000_010_0_011100110001;
      patterns[40131] = 29'b1_001110011000_011_0_111001100010;
      patterns[40132] = 29'b1_001110011000_100_0_100111001100;
      patterns[40133] = 29'b1_001110011000_101_0_010011100110;
      patterns[40134] = 29'b1_001110011000_110_1_001110011000;
      patterns[40135] = 29'b1_001110011000_111_1_001110011000;
      patterns[40136] = 29'b1_001110011001_000_1_001110011001;
      patterns[40137] = 29'b1_001110011001_001_1_011001001110;
      patterns[40138] = 29'b1_001110011001_010_0_011100110011;
      patterns[40139] = 29'b1_001110011001_011_0_111001100110;
      patterns[40140] = 29'b1_001110011001_100_1_100111001100;
      patterns[40141] = 29'b1_001110011001_101_0_110011100110;
      patterns[40142] = 29'b1_001110011001_110_1_001110011001;
      patterns[40143] = 29'b1_001110011001_111_1_001110011001;
      patterns[40144] = 29'b1_001110011010_000_1_001110011010;
      patterns[40145] = 29'b1_001110011010_001_1_011010001110;
      patterns[40146] = 29'b1_001110011010_010_0_011100110101;
      patterns[40147] = 29'b1_001110011010_011_0_111001101010;
      patterns[40148] = 29'b1_001110011010_100_0_100111001101;
      patterns[40149] = 29'b1_001110011010_101_1_010011100110;
      patterns[40150] = 29'b1_001110011010_110_1_001110011010;
      patterns[40151] = 29'b1_001110011010_111_1_001110011010;
      patterns[40152] = 29'b1_001110011011_000_1_001110011011;
      patterns[40153] = 29'b1_001110011011_001_1_011011001110;
      patterns[40154] = 29'b1_001110011011_010_0_011100110111;
      patterns[40155] = 29'b1_001110011011_011_0_111001101110;
      patterns[40156] = 29'b1_001110011011_100_1_100111001101;
      patterns[40157] = 29'b1_001110011011_101_1_110011100110;
      patterns[40158] = 29'b1_001110011011_110_1_001110011011;
      patterns[40159] = 29'b1_001110011011_111_1_001110011011;
      patterns[40160] = 29'b1_001110011100_000_1_001110011100;
      patterns[40161] = 29'b1_001110011100_001_1_011100001110;
      patterns[40162] = 29'b1_001110011100_010_0_011100111001;
      patterns[40163] = 29'b1_001110011100_011_0_111001110010;
      patterns[40164] = 29'b1_001110011100_100_0_100111001110;
      patterns[40165] = 29'b1_001110011100_101_0_010011100111;
      patterns[40166] = 29'b1_001110011100_110_1_001110011100;
      patterns[40167] = 29'b1_001110011100_111_1_001110011100;
      patterns[40168] = 29'b1_001110011101_000_1_001110011101;
      patterns[40169] = 29'b1_001110011101_001_1_011101001110;
      patterns[40170] = 29'b1_001110011101_010_0_011100111011;
      patterns[40171] = 29'b1_001110011101_011_0_111001110110;
      patterns[40172] = 29'b1_001110011101_100_1_100111001110;
      patterns[40173] = 29'b1_001110011101_101_0_110011100111;
      patterns[40174] = 29'b1_001110011101_110_1_001110011101;
      patterns[40175] = 29'b1_001110011101_111_1_001110011101;
      patterns[40176] = 29'b1_001110011110_000_1_001110011110;
      patterns[40177] = 29'b1_001110011110_001_1_011110001110;
      patterns[40178] = 29'b1_001110011110_010_0_011100111101;
      patterns[40179] = 29'b1_001110011110_011_0_111001111010;
      patterns[40180] = 29'b1_001110011110_100_0_100111001111;
      patterns[40181] = 29'b1_001110011110_101_1_010011100111;
      patterns[40182] = 29'b1_001110011110_110_1_001110011110;
      patterns[40183] = 29'b1_001110011110_111_1_001110011110;
      patterns[40184] = 29'b1_001110011111_000_1_001110011111;
      patterns[40185] = 29'b1_001110011111_001_1_011111001110;
      patterns[40186] = 29'b1_001110011111_010_0_011100111111;
      patterns[40187] = 29'b1_001110011111_011_0_111001111110;
      patterns[40188] = 29'b1_001110011111_100_1_100111001111;
      patterns[40189] = 29'b1_001110011111_101_1_110011100111;
      patterns[40190] = 29'b1_001110011111_110_1_001110011111;
      patterns[40191] = 29'b1_001110011111_111_1_001110011111;
      patterns[40192] = 29'b1_001110100000_000_1_001110100000;
      patterns[40193] = 29'b1_001110100000_001_1_100000001110;
      patterns[40194] = 29'b1_001110100000_010_0_011101000001;
      patterns[40195] = 29'b1_001110100000_011_0_111010000010;
      patterns[40196] = 29'b1_001110100000_100_0_100111010000;
      patterns[40197] = 29'b1_001110100000_101_0_010011101000;
      patterns[40198] = 29'b1_001110100000_110_1_001110100000;
      patterns[40199] = 29'b1_001110100000_111_1_001110100000;
      patterns[40200] = 29'b1_001110100001_000_1_001110100001;
      patterns[40201] = 29'b1_001110100001_001_1_100001001110;
      patterns[40202] = 29'b1_001110100001_010_0_011101000011;
      patterns[40203] = 29'b1_001110100001_011_0_111010000110;
      patterns[40204] = 29'b1_001110100001_100_1_100111010000;
      patterns[40205] = 29'b1_001110100001_101_0_110011101000;
      patterns[40206] = 29'b1_001110100001_110_1_001110100001;
      patterns[40207] = 29'b1_001110100001_111_1_001110100001;
      patterns[40208] = 29'b1_001110100010_000_1_001110100010;
      patterns[40209] = 29'b1_001110100010_001_1_100010001110;
      patterns[40210] = 29'b1_001110100010_010_0_011101000101;
      patterns[40211] = 29'b1_001110100010_011_0_111010001010;
      patterns[40212] = 29'b1_001110100010_100_0_100111010001;
      patterns[40213] = 29'b1_001110100010_101_1_010011101000;
      patterns[40214] = 29'b1_001110100010_110_1_001110100010;
      patterns[40215] = 29'b1_001110100010_111_1_001110100010;
      patterns[40216] = 29'b1_001110100011_000_1_001110100011;
      patterns[40217] = 29'b1_001110100011_001_1_100011001110;
      patterns[40218] = 29'b1_001110100011_010_0_011101000111;
      patterns[40219] = 29'b1_001110100011_011_0_111010001110;
      patterns[40220] = 29'b1_001110100011_100_1_100111010001;
      patterns[40221] = 29'b1_001110100011_101_1_110011101000;
      patterns[40222] = 29'b1_001110100011_110_1_001110100011;
      patterns[40223] = 29'b1_001110100011_111_1_001110100011;
      patterns[40224] = 29'b1_001110100100_000_1_001110100100;
      patterns[40225] = 29'b1_001110100100_001_1_100100001110;
      patterns[40226] = 29'b1_001110100100_010_0_011101001001;
      patterns[40227] = 29'b1_001110100100_011_0_111010010010;
      patterns[40228] = 29'b1_001110100100_100_0_100111010010;
      patterns[40229] = 29'b1_001110100100_101_0_010011101001;
      patterns[40230] = 29'b1_001110100100_110_1_001110100100;
      patterns[40231] = 29'b1_001110100100_111_1_001110100100;
      patterns[40232] = 29'b1_001110100101_000_1_001110100101;
      patterns[40233] = 29'b1_001110100101_001_1_100101001110;
      patterns[40234] = 29'b1_001110100101_010_0_011101001011;
      patterns[40235] = 29'b1_001110100101_011_0_111010010110;
      patterns[40236] = 29'b1_001110100101_100_1_100111010010;
      patterns[40237] = 29'b1_001110100101_101_0_110011101001;
      patterns[40238] = 29'b1_001110100101_110_1_001110100101;
      patterns[40239] = 29'b1_001110100101_111_1_001110100101;
      patterns[40240] = 29'b1_001110100110_000_1_001110100110;
      patterns[40241] = 29'b1_001110100110_001_1_100110001110;
      patterns[40242] = 29'b1_001110100110_010_0_011101001101;
      patterns[40243] = 29'b1_001110100110_011_0_111010011010;
      patterns[40244] = 29'b1_001110100110_100_0_100111010011;
      patterns[40245] = 29'b1_001110100110_101_1_010011101001;
      patterns[40246] = 29'b1_001110100110_110_1_001110100110;
      patterns[40247] = 29'b1_001110100110_111_1_001110100110;
      patterns[40248] = 29'b1_001110100111_000_1_001110100111;
      patterns[40249] = 29'b1_001110100111_001_1_100111001110;
      patterns[40250] = 29'b1_001110100111_010_0_011101001111;
      patterns[40251] = 29'b1_001110100111_011_0_111010011110;
      patterns[40252] = 29'b1_001110100111_100_1_100111010011;
      patterns[40253] = 29'b1_001110100111_101_1_110011101001;
      patterns[40254] = 29'b1_001110100111_110_1_001110100111;
      patterns[40255] = 29'b1_001110100111_111_1_001110100111;
      patterns[40256] = 29'b1_001110101000_000_1_001110101000;
      patterns[40257] = 29'b1_001110101000_001_1_101000001110;
      patterns[40258] = 29'b1_001110101000_010_0_011101010001;
      patterns[40259] = 29'b1_001110101000_011_0_111010100010;
      patterns[40260] = 29'b1_001110101000_100_0_100111010100;
      patterns[40261] = 29'b1_001110101000_101_0_010011101010;
      patterns[40262] = 29'b1_001110101000_110_1_001110101000;
      patterns[40263] = 29'b1_001110101000_111_1_001110101000;
      patterns[40264] = 29'b1_001110101001_000_1_001110101001;
      patterns[40265] = 29'b1_001110101001_001_1_101001001110;
      patterns[40266] = 29'b1_001110101001_010_0_011101010011;
      patterns[40267] = 29'b1_001110101001_011_0_111010100110;
      patterns[40268] = 29'b1_001110101001_100_1_100111010100;
      patterns[40269] = 29'b1_001110101001_101_0_110011101010;
      patterns[40270] = 29'b1_001110101001_110_1_001110101001;
      patterns[40271] = 29'b1_001110101001_111_1_001110101001;
      patterns[40272] = 29'b1_001110101010_000_1_001110101010;
      patterns[40273] = 29'b1_001110101010_001_1_101010001110;
      patterns[40274] = 29'b1_001110101010_010_0_011101010101;
      patterns[40275] = 29'b1_001110101010_011_0_111010101010;
      patterns[40276] = 29'b1_001110101010_100_0_100111010101;
      patterns[40277] = 29'b1_001110101010_101_1_010011101010;
      patterns[40278] = 29'b1_001110101010_110_1_001110101010;
      patterns[40279] = 29'b1_001110101010_111_1_001110101010;
      patterns[40280] = 29'b1_001110101011_000_1_001110101011;
      patterns[40281] = 29'b1_001110101011_001_1_101011001110;
      patterns[40282] = 29'b1_001110101011_010_0_011101010111;
      patterns[40283] = 29'b1_001110101011_011_0_111010101110;
      patterns[40284] = 29'b1_001110101011_100_1_100111010101;
      patterns[40285] = 29'b1_001110101011_101_1_110011101010;
      patterns[40286] = 29'b1_001110101011_110_1_001110101011;
      patterns[40287] = 29'b1_001110101011_111_1_001110101011;
      patterns[40288] = 29'b1_001110101100_000_1_001110101100;
      patterns[40289] = 29'b1_001110101100_001_1_101100001110;
      patterns[40290] = 29'b1_001110101100_010_0_011101011001;
      patterns[40291] = 29'b1_001110101100_011_0_111010110010;
      patterns[40292] = 29'b1_001110101100_100_0_100111010110;
      patterns[40293] = 29'b1_001110101100_101_0_010011101011;
      patterns[40294] = 29'b1_001110101100_110_1_001110101100;
      patterns[40295] = 29'b1_001110101100_111_1_001110101100;
      patterns[40296] = 29'b1_001110101101_000_1_001110101101;
      patterns[40297] = 29'b1_001110101101_001_1_101101001110;
      patterns[40298] = 29'b1_001110101101_010_0_011101011011;
      patterns[40299] = 29'b1_001110101101_011_0_111010110110;
      patterns[40300] = 29'b1_001110101101_100_1_100111010110;
      patterns[40301] = 29'b1_001110101101_101_0_110011101011;
      patterns[40302] = 29'b1_001110101101_110_1_001110101101;
      patterns[40303] = 29'b1_001110101101_111_1_001110101101;
      patterns[40304] = 29'b1_001110101110_000_1_001110101110;
      patterns[40305] = 29'b1_001110101110_001_1_101110001110;
      patterns[40306] = 29'b1_001110101110_010_0_011101011101;
      patterns[40307] = 29'b1_001110101110_011_0_111010111010;
      patterns[40308] = 29'b1_001110101110_100_0_100111010111;
      patterns[40309] = 29'b1_001110101110_101_1_010011101011;
      patterns[40310] = 29'b1_001110101110_110_1_001110101110;
      patterns[40311] = 29'b1_001110101110_111_1_001110101110;
      patterns[40312] = 29'b1_001110101111_000_1_001110101111;
      patterns[40313] = 29'b1_001110101111_001_1_101111001110;
      patterns[40314] = 29'b1_001110101111_010_0_011101011111;
      patterns[40315] = 29'b1_001110101111_011_0_111010111110;
      patterns[40316] = 29'b1_001110101111_100_1_100111010111;
      patterns[40317] = 29'b1_001110101111_101_1_110011101011;
      patterns[40318] = 29'b1_001110101111_110_1_001110101111;
      patterns[40319] = 29'b1_001110101111_111_1_001110101111;
      patterns[40320] = 29'b1_001110110000_000_1_001110110000;
      patterns[40321] = 29'b1_001110110000_001_1_110000001110;
      patterns[40322] = 29'b1_001110110000_010_0_011101100001;
      patterns[40323] = 29'b1_001110110000_011_0_111011000010;
      patterns[40324] = 29'b1_001110110000_100_0_100111011000;
      patterns[40325] = 29'b1_001110110000_101_0_010011101100;
      patterns[40326] = 29'b1_001110110000_110_1_001110110000;
      patterns[40327] = 29'b1_001110110000_111_1_001110110000;
      patterns[40328] = 29'b1_001110110001_000_1_001110110001;
      patterns[40329] = 29'b1_001110110001_001_1_110001001110;
      patterns[40330] = 29'b1_001110110001_010_0_011101100011;
      patterns[40331] = 29'b1_001110110001_011_0_111011000110;
      patterns[40332] = 29'b1_001110110001_100_1_100111011000;
      patterns[40333] = 29'b1_001110110001_101_0_110011101100;
      patterns[40334] = 29'b1_001110110001_110_1_001110110001;
      patterns[40335] = 29'b1_001110110001_111_1_001110110001;
      patterns[40336] = 29'b1_001110110010_000_1_001110110010;
      patterns[40337] = 29'b1_001110110010_001_1_110010001110;
      patterns[40338] = 29'b1_001110110010_010_0_011101100101;
      patterns[40339] = 29'b1_001110110010_011_0_111011001010;
      patterns[40340] = 29'b1_001110110010_100_0_100111011001;
      patterns[40341] = 29'b1_001110110010_101_1_010011101100;
      patterns[40342] = 29'b1_001110110010_110_1_001110110010;
      patterns[40343] = 29'b1_001110110010_111_1_001110110010;
      patterns[40344] = 29'b1_001110110011_000_1_001110110011;
      patterns[40345] = 29'b1_001110110011_001_1_110011001110;
      patterns[40346] = 29'b1_001110110011_010_0_011101100111;
      patterns[40347] = 29'b1_001110110011_011_0_111011001110;
      patterns[40348] = 29'b1_001110110011_100_1_100111011001;
      patterns[40349] = 29'b1_001110110011_101_1_110011101100;
      patterns[40350] = 29'b1_001110110011_110_1_001110110011;
      patterns[40351] = 29'b1_001110110011_111_1_001110110011;
      patterns[40352] = 29'b1_001110110100_000_1_001110110100;
      patterns[40353] = 29'b1_001110110100_001_1_110100001110;
      patterns[40354] = 29'b1_001110110100_010_0_011101101001;
      patterns[40355] = 29'b1_001110110100_011_0_111011010010;
      patterns[40356] = 29'b1_001110110100_100_0_100111011010;
      patterns[40357] = 29'b1_001110110100_101_0_010011101101;
      patterns[40358] = 29'b1_001110110100_110_1_001110110100;
      patterns[40359] = 29'b1_001110110100_111_1_001110110100;
      patterns[40360] = 29'b1_001110110101_000_1_001110110101;
      patterns[40361] = 29'b1_001110110101_001_1_110101001110;
      patterns[40362] = 29'b1_001110110101_010_0_011101101011;
      patterns[40363] = 29'b1_001110110101_011_0_111011010110;
      patterns[40364] = 29'b1_001110110101_100_1_100111011010;
      patterns[40365] = 29'b1_001110110101_101_0_110011101101;
      patterns[40366] = 29'b1_001110110101_110_1_001110110101;
      patterns[40367] = 29'b1_001110110101_111_1_001110110101;
      patterns[40368] = 29'b1_001110110110_000_1_001110110110;
      patterns[40369] = 29'b1_001110110110_001_1_110110001110;
      patterns[40370] = 29'b1_001110110110_010_0_011101101101;
      patterns[40371] = 29'b1_001110110110_011_0_111011011010;
      patterns[40372] = 29'b1_001110110110_100_0_100111011011;
      patterns[40373] = 29'b1_001110110110_101_1_010011101101;
      patterns[40374] = 29'b1_001110110110_110_1_001110110110;
      patterns[40375] = 29'b1_001110110110_111_1_001110110110;
      patterns[40376] = 29'b1_001110110111_000_1_001110110111;
      patterns[40377] = 29'b1_001110110111_001_1_110111001110;
      patterns[40378] = 29'b1_001110110111_010_0_011101101111;
      patterns[40379] = 29'b1_001110110111_011_0_111011011110;
      patterns[40380] = 29'b1_001110110111_100_1_100111011011;
      patterns[40381] = 29'b1_001110110111_101_1_110011101101;
      patterns[40382] = 29'b1_001110110111_110_1_001110110111;
      patterns[40383] = 29'b1_001110110111_111_1_001110110111;
      patterns[40384] = 29'b1_001110111000_000_1_001110111000;
      patterns[40385] = 29'b1_001110111000_001_1_111000001110;
      patterns[40386] = 29'b1_001110111000_010_0_011101110001;
      patterns[40387] = 29'b1_001110111000_011_0_111011100010;
      patterns[40388] = 29'b1_001110111000_100_0_100111011100;
      patterns[40389] = 29'b1_001110111000_101_0_010011101110;
      patterns[40390] = 29'b1_001110111000_110_1_001110111000;
      patterns[40391] = 29'b1_001110111000_111_1_001110111000;
      patterns[40392] = 29'b1_001110111001_000_1_001110111001;
      patterns[40393] = 29'b1_001110111001_001_1_111001001110;
      patterns[40394] = 29'b1_001110111001_010_0_011101110011;
      patterns[40395] = 29'b1_001110111001_011_0_111011100110;
      patterns[40396] = 29'b1_001110111001_100_1_100111011100;
      patterns[40397] = 29'b1_001110111001_101_0_110011101110;
      patterns[40398] = 29'b1_001110111001_110_1_001110111001;
      patterns[40399] = 29'b1_001110111001_111_1_001110111001;
      patterns[40400] = 29'b1_001110111010_000_1_001110111010;
      patterns[40401] = 29'b1_001110111010_001_1_111010001110;
      patterns[40402] = 29'b1_001110111010_010_0_011101110101;
      patterns[40403] = 29'b1_001110111010_011_0_111011101010;
      patterns[40404] = 29'b1_001110111010_100_0_100111011101;
      patterns[40405] = 29'b1_001110111010_101_1_010011101110;
      patterns[40406] = 29'b1_001110111010_110_1_001110111010;
      patterns[40407] = 29'b1_001110111010_111_1_001110111010;
      patterns[40408] = 29'b1_001110111011_000_1_001110111011;
      patterns[40409] = 29'b1_001110111011_001_1_111011001110;
      patterns[40410] = 29'b1_001110111011_010_0_011101110111;
      patterns[40411] = 29'b1_001110111011_011_0_111011101110;
      patterns[40412] = 29'b1_001110111011_100_1_100111011101;
      patterns[40413] = 29'b1_001110111011_101_1_110011101110;
      patterns[40414] = 29'b1_001110111011_110_1_001110111011;
      patterns[40415] = 29'b1_001110111011_111_1_001110111011;
      patterns[40416] = 29'b1_001110111100_000_1_001110111100;
      patterns[40417] = 29'b1_001110111100_001_1_111100001110;
      patterns[40418] = 29'b1_001110111100_010_0_011101111001;
      patterns[40419] = 29'b1_001110111100_011_0_111011110010;
      patterns[40420] = 29'b1_001110111100_100_0_100111011110;
      patterns[40421] = 29'b1_001110111100_101_0_010011101111;
      patterns[40422] = 29'b1_001110111100_110_1_001110111100;
      patterns[40423] = 29'b1_001110111100_111_1_001110111100;
      patterns[40424] = 29'b1_001110111101_000_1_001110111101;
      patterns[40425] = 29'b1_001110111101_001_1_111101001110;
      patterns[40426] = 29'b1_001110111101_010_0_011101111011;
      patterns[40427] = 29'b1_001110111101_011_0_111011110110;
      patterns[40428] = 29'b1_001110111101_100_1_100111011110;
      patterns[40429] = 29'b1_001110111101_101_0_110011101111;
      patterns[40430] = 29'b1_001110111101_110_1_001110111101;
      patterns[40431] = 29'b1_001110111101_111_1_001110111101;
      patterns[40432] = 29'b1_001110111110_000_1_001110111110;
      patterns[40433] = 29'b1_001110111110_001_1_111110001110;
      patterns[40434] = 29'b1_001110111110_010_0_011101111101;
      patterns[40435] = 29'b1_001110111110_011_0_111011111010;
      patterns[40436] = 29'b1_001110111110_100_0_100111011111;
      patterns[40437] = 29'b1_001110111110_101_1_010011101111;
      patterns[40438] = 29'b1_001110111110_110_1_001110111110;
      patterns[40439] = 29'b1_001110111110_111_1_001110111110;
      patterns[40440] = 29'b1_001110111111_000_1_001110111111;
      patterns[40441] = 29'b1_001110111111_001_1_111111001110;
      patterns[40442] = 29'b1_001110111111_010_0_011101111111;
      patterns[40443] = 29'b1_001110111111_011_0_111011111110;
      patterns[40444] = 29'b1_001110111111_100_1_100111011111;
      patterns[40445] = 29'b1_001110111111_101_1_110011101111;
      patterns[40446] = 29'b1_001110111111_110_1_001110111111;
      patterns[40447] = 29'b1_001110111111_111_1_001110111111;
      patterns[40448] = 29'b1_001111000000_000_1_001111000000;
      patterns[40449] = 29'b1_001111000000_001_1_000000001111;
      patterns[40450] = 29'b1_001111000000_010_0_011110000001;
      patterns[40451] = 29'b1_001111000000_011_0_111100000010;
      patterns[40452] = 29'b1_001111000000_100_0_100111100000;
      patterns[40453] = 29'b1_001111000000_101_0_010011110000;
      patterns[40454] = 29'b1_001111000000_110_1_001111000000;
      patterns[40455] = 29'b1_001111000000_111_1_001111000000;
      patterns[40456] = 29'b1_001111000001_000_1_001111000001;
      patterns[40457] = 29'b1_001111000001_001_1_000001001111;
      patterns[40458] = 29'b1_001111000001_010_0_011110000011;
      patterns[40459] = 29'b1_001111000001_011_0_111100000110;
      patterns[40460] = 29'b1_001111000001_100_1_100111100000;
      patterns[40461] = 29'b1_001111000001_101_0_110011110000;
      patterns[40462] = 29'b1_001111000001_110_1_001111000001;
      patterns[40463] = 29'b1_001111000001_111_1_001111000001;
      patterns[40464] = 29'b1_001111000010_000_1_001111000010;
      patterns[40465] = 29'b1_001111000010_001_1_000010001111;
      patterns[40466] = 29'b1_001111000010_010_0_011110000101;
      patterns[40467] = 29'b1_001111000010_011_0_111100001010;
      patterns[40468] = 29'b1_001111000010_100_0_100111100001;
      patterns[40469] = 29'b1_001111000010_101_1_010011110000;
      patterns[40470] = 29'b1_001111000010_110_1_001111000010;
      patterns[40471] = 29'b1_001111000010_111_1_001111000010;
      patterns[40472] = 29'b1_001111000011_000_1_001111000011;
      patterns[40473] = 29'b1_001111000011_001_1_000011001111;
      patterns[40474] = 29'b1_001111000011_010_0_011110000111;
      patterns[40475] = 29'b1_001111000011_011_0_111100001110;
      patterns[40476] = 29'b1_001111000011_100_1_100111100001;
      patterns[40477] = 29'b1_001111000011_101_1_110011110000;
      patterns[40478] = 29'b1_001111000011_110_1_001111000011;
      patterns[40479] = 29'b1_001111000011_111_1_001111000011;
      patterns[40480] = 29'b1_001111000100_000_1_001111000100;
      patterns[40481] = 29'b1_001111000100_001_1_000100001111;
      patterns[40482] = 29'b1_001111000100_010_0_011110001001;
      patterns[40483] = 29'b1_001111000100_011_0_111100010010;
      patterns[40484] = 29'b1_001111000100_100_0_100111100010;
      patterns[40485] = 29'b1_001111000100_101_0_010011110001;
      patterns[40486] = 29'b1_001111000100_110_1_001111000100;
      patterns[40487] = 29'b1_001111000100_111_1_001111000100;
      patterns[40488] = 29'b1_001111000101_000_1_001111000101;
      patterns[40489] = 29'b1_001111000101_001_1_000101001111;
      patterns[40490] = 29'b1_001111000101_010_0_011110001011;
      patterns[40491] = 29'b1_001111000101_011_0_111100010110;
      patterns[40492] = 29'b1_001111000101_100_1_100111100010;
      patterns[40493] = 29'b1_001111000101_101_0_110011110001;
      patterns[40494] = 29'b1_001111000101_110_1_001111000101;
      patterns[40495] = 29'b1_001111000101_111_1_001111000101;
      patterns[40496] = 29'b1_001111000110_000_1_001111000110;
      patterns[40497] = 29'b1_001111000110_001_1_000110001111;
      patterns[40498] = 29'b1_001111000110_010_0_011110001101;
      patterns[40499] = 29'b1_001111000110_011_0_111100011010;
      patterns[40500] = 29'b1_001111000110_100_0_100111100011;
      patterns[40501] = 29'b1_001111000110_101_1_010011110001;
      patterns[40502] = 29'b1_001111000110_110_1_001111000110;
      patterns[40503] = 29'b1_001111000110_111_1_001111000110;
      patterns[40504] = 29'b1_001111000111_000_1_001111000111;
      patterns[40505] = 29'b1_001111000111_001_1_000111001111;
      patterns[40506] = 29'b1_001111000111_010_0_011110001111;
      patterns[40507] = 29'b1_001111000111_011_0_111100011110;
      patterns[40508] = 29'b1_001111000111_100_1_100111100011;
      patterns[40509] = 29'b1_001111000111_101_1_110011110001;
      patterns[40510] = 29'b1_001111000111_110_1_001111000111;
      patterns[40511] = 29'b1_001111000111_111_1_001111000111;
      patterns[40512] = 29'b1_001111001000_000_1_001111001000;
      patterns[40513] = 29'b1_001111001000_001_1_001000001111;
      patterns[40514] = 29'b1_001111001000_010_0_011110010001;
      patterns[40515] = 29'b1_001111001000_011_0_111100100010;
      patterns[40516] = 29'b1_001111001000_100_0_100111100100;
      patterns[40517] = 29'b1_001111001000_101_0_010011110010;
      patterns[40518] = 29'b1_001111001000_110_1_001111001000;
      patterns[40519] = 29'b1_001111001000_111_1_001111001000;
      patterns[40520] = 29'b1_001111001001_000_1_001111001001;
      patterns[40521] = 29'b1_001111001001_001_1_001001001111;
      patterns[40522] = 29'b1_001111001001_010_0_011110010011;
      patterns[40523] = 29'b1_001111001001_011_0_111100100110;
      patterns[40524] = 29'b1_001111001001_100_1_100111100100;
      patterns[40525] = 29'b1_001111001001_101_0_110011110010;
      patterns[40526] = 29'b1_001111001001_110_1_001111001001;
      patterns[40527] = 29'b1_001111001001_111_1_001111001001;
      patterns[40528] = 29'b1_001111001010_000_1_001111001010;
      patterns[40529] = 29'b1_001111001010_001_1_001010001111;
      patterns[40530] = 29'b1_001111001010_010_0_011110010101;
      patterns[40531] = 29'b1_001111001010_011_0_111100101010;
      patterns[40532] = 29'b1_001111001010_100_0_100111100101;
      patterns[40533] = 29'b1_001111001010_101_1_010011110010;
      patterns[40534] = 29'b1_001111001010_110_1_001111001010;
      patterns[40535] = 29'b1_001111001010_111_1_001111001010;
      patterns[40536] = 29'b1_001111001011_000_1_001111001011;
      patterns[40537] = 29'b1_001111001011_001_1_001011001111;
      patterns[40538] = 29'b1_001111001011_010_0_011110010111;
      patterns[40539] = 29'b1_001111001011_011_0_111100101110;
      patterns[40540] = 29'b1_001111001011_100_1_100111100101;
      patterns[40541] = 29'b1_001111001011_101_1_110011110010;
      patterns[40542] = 29'b1_001111001011_110_1_001111001011;
      patterns[40543] = 29'b1_001111001011_111_1_001111001011;
      patterns[40544] = 29'b1_001111001100_000_1_001111001100;
      patterns[40545] = 29'b1_001111001100_001_1_001100001111;
      patterns[40546] = 29'b1_001111001100_010_0_011110011001;
      patterns[40547] = 29'b1_001111001100_011_0_111100110010;
      patterns[40548] = 29'b1_001111001100_100_0_100111100110;
      patterns[40549] = 29'b1_001111001100_101_0_010011110011;
      patterns[40550] = 29'b1_001111001100_110_1_001111001100;
      patterns[40551] = 29'b1_001111001100_111_1_001111001100;
      patterns[40552] = 29'b1_001111001101_000_1_001111001101;
      patterns[40553] = 29'b1_001111001101_001_1_001101001111;
      patterns[40554] = 29'b1_001111001101_010_0_011110011011;
      patterns[40555] = 29'b1_001111001101_011_0_111100110110;
      patterns[40556] = 29'b1_001111001101_100_1_100111100110;
      patterns[40557] = 29'b1_001111001101_101_0_110011110011;
      patterns[40558] = 29'b1_001111001101_110_1_001111001101;
      patterns[40559] = 29'b1_001111001101_111_1_001111001101;
      patterns[40560] = 29'b1_001111001110_000_1_001111001110;
      patterns[40561] = 29'b1_001111001110_001_1_001110001111;
      patterns[40562] = 29'b1_001111001110_010_0_011110011101;
      patterns[40563] = 29'b1_001111001110_011_0_111100111010;
      patterns[40564] = 29'b1_001111001110_100_0_100111100111;
      patterns[40565] = 29'b1_001111001110_101_1_010011110011;
      patterns[40566] = 29'b1_001111001110_110_1_001111001110;
      patterns[40567] = 29'b1_001111001110_111_1_001111001110;
      patterns[40568] = 29'b1_001111001111_000_1_001111001111;
      patterns[40569] = 29'b1_001111001111_001_1_001111001111;
      patterns[40570] = 29'b1_001111001111_010_0_011110011111;
      patterns[40571] = 29'b1_001111001111_011_0_111100111110;
      patterns[40572] = 29'b1_001111001111_100_1_100111100111;
      patterns[40573] = 29'b1_001111001111_101_1_110011110011;
      patterns[40574] = 29'b1_001111001111_110_1_001111001111;
      patterns[40575] = 29'b1_001111001111_111_1_001111001111;
      patterns[40576] = 29'b1_001111010000_000_1_001111010000;
      patterns[40577] = 29'b1_001111010000_001_1_010000001111;
      patterns[40578] = 29'b1_001111010000_010_0_011110100001;
      patterns[40579] = 29'b1_001111010000_011_0_111101000010;
      patterns[40580] = 29'b1_001111010000_100_0_100111101000;
      patterns[40581] = 29'b1_001111010000_101_0_010011110100;
      patterns[40582] = 29'b1_001111010000_110_1_001111010000;
      patterns[40583] = 29'b1_001111010000_111_1_001111010000;
      patterns[40584] = 29'b1_001111010001_000_1_001111010001;
      patterns[40585] = 29'b1_001111010001_001_1_010001001111;
      patterns[40586] = 29'b1_001111010001_010_0_011110100011;
      patterns[40587] = 29'b1_001111010001_011_0_111101000110;
      patterns[40588] = 29'b1_001111010001_100_1_100111101000;
      patterns[40589] = 29'b1_001111010001_101_0_110011110100;
      patterns[40590] = 29'b1_001111010001_110_1_001111010001;
      patterns[40591] = 29'b1_001111010001_111_1_001111010001;
      patterns[40592] = 29'b1_001111010010_000_1_001111010010;
      patterns[40593] = 29'b1_001111010010_001_1_010010001111;
      patterns[40594] = 29'b1_001111010010_010_0_011110100101;
      patterns[40595] = 29'b1_001111010010_011_0_111101001010;
      patterns[40596] = 29'b1_001111010010_100_0_100111101001;
      patterns[40597] = 29'b1_001111010010_101_1_010011110100;
      patterns[40598] = 29'b1_001111010010_110_1_001111010010;
      patterns[40599] = 29'b1_001111010010_111_1_001111010010;
      patterns[40600] = 29'b1_001111010011_000_1_001111010011;
      patterns[40601] = 29'b1_001111010011_001_1_010011001111;
      patterns[40602] = 29'b1_001111010011_010_0_011110100111;
      patterns[40603] = 29'b1_001111010011_011_0_111101001110;
      patterns[40604] = 29'b1_001111010011_100_1_100111101001;
      patterns[40605] = 29'b1_001111010011_101_1_110011110100;
      patterns[40606] = 29'b1_001111010011_110_1_001111010011;
      patterns[40607] = 29'b1_001111010011_111_1_001111010011;
      patterns[40608] = 29'b1_001111010100_000_1_001111010100;
      patterns[40609] = 29'b1_001111010100_001_1_010100001111;
      patterns[40610] = 29'b1_001111010100_010_0_011110101001;
      patterns[40611] = 29'b1_001111010100_011_0_111101010010;
      patterns[40612] = 29'b1_001111010100_100_0_100111101010;
      patterns[40613] = 29'b1_001111010100_101_0_010011110101;
      patterns[40614] = 29'b1_001111010100_110_1_001111010100;
      patterns[40615] = 29'b1_001111010100_111_1_001111010100;
      patterns[40616] = 29'b1_001111010101_000_1_001111010101;
      patterns[40617] = 29'b1_001111010101_001_1_010101001111;
      patterns[40618] = 29'b1_001111010101_010_0_011110101011;
      patterns[40619] = 29'b1_001111010101_011_0_111101010110;
      patterns[40620] = 29'b1_001111010101_100_1_100111101010;
      patterns[40621] = 29'b1_001111010101_101_0_110011110101;
      patterns[40622] = 29'b1_001111010101_110_1_001111010101;
      patterns[40623] = 29'b1_001111010101_111_1_001111010101;
      patterns[40624] = 29'b1_001111010110_000_1_001111010110;
      patterns[40625] = 29'b1_001111010110_001_1_010110001111;
      patterns[40626] = 29'b1_001111010110_010_0_011110101101;
      patterns[40627] = 29'b1_001111010110_011_0_111101011010;
      patterns[40628] = 29'b1_001111010110_100_0_100111101011;
      patterns[40629] = 29'b1_001111010110_101_1_010011110101;
      patterns[40630] = 29'b1_001111010110_110_1_001111010110;
      patterns[40631] = 29'b1_001111010110_111_1_001111010110;
      patterns[40632] = 29'b1_001111010111_000_1_001111010111;
      patterns[40633] = 29'b1_001111010111_001_1_010111001111;
      patterns[40634] = 29'b1_001111010111_010_0_011110101111;
      patterns[40635] = 29'b1_001111010111_011_0_111101011110;
      patterns[40636] = 29'b1_001111010111_100_1_100111101011;
      patterns[40637] = 29'b1_001111010111_101_1_110011110101;
      patterns[40638] = 29'b1_001111010111_110_1_001111010111;
      patterns[40639] = 29'b1_001111010111_111_1_001111010111;
      patterns[40640] = 29'b1_001111011000_000_1_001111011000;
      patterns[40641] = 29'b1_001111011000_001_1_011000001111;
      patterns[40642] = 29'b1_001111011000_010_0_011110110001;
      patterns[40643] = 29'b1_001111011000_011_0_111101100010;
      patterns[40644] = 29'b1_001111011000_100_0_100111101100;
      patterns[40645] = 29'b1_001111011000_101_0_010011110110;
      patterns[40646] = 29'b1_001111011000_110_1_001111011000;
      patterns[40647] = 29'b1_001111011000_111_1_001111011000;
      patterns[40648] = 29'b1_001111011001_000_1_001111011001;
      patterns[40649] = 29'b1_001111011001_001_1_011001001111;
      patterns[40650] = 29'b1_001111011001_010_0_011110110011;
      patterns[40651] = 29'b1_001111011001_011_0_111101100110;
      patterns[40652] = 29'b1_001111011001_100_1_100111101100;
      patterns[40653] = 29'b1_001111011001_101_0_110011110110;
      patterns[40654] = 29'b1_001111011001_110_1_001111011001;
      patterns[40655] = 29'b1_001111011001_111_1_001111011001;
      patterns[40656] = 29'b1_001111011010_000_1_001111011010;
      patterns[40657] = 29'b1_001111011010_001_1_011010001111;
      patterns[40658] = 29'b1_001111011010_010_0_011110110101;
      patterns[40659] = 29'b1_001111011010_011_0_111101101010;
      patterns[40660] = 29'b1_001111011010_100_0_100111101101;
      patterns[40661] = 29'b1_001111011010_101_1_010011110110;
      patterns[40662] = 29'b1_001111011010_110_1_001111011010;
      patterns[40663] = 29'b1_001111011010_111_1_001111011010;
      patterns[40664] = 29'b1_001111011011_000_1_001111011011;
      patterns[40665] = 29'b1_001111011011_001_1_011011001111;
      patterns[40666] = 29'b1_001111011011_010_0_011110110111;
      patterns[40667] = 29'b1_001111011011_011_0_111101101110;
      patterns[40668] = 29'b1_001111011011_100_1_100111101101;
      patterns[40669] = 29'b1_001111011011_101_1_110011110110;
      patterns[40670] = 29'b1_001111011011_110_1_001111011011;
      patterns[40671] = 29'b1_001111011011_111_1_001111011011;
      patterns[40672] = 29'b1_001111011100_000_1_001111011100;
      patterns[40673] = 29'b1_001111011100_001_1_011100001111;
      patterns[40674] = 29'b1_001111011100_010_0_011110111001;
      patterns[40675] = 29'b1_001111011100_011_0_111101110010;
      patterns[40676] = 29'b1_001111011100_100_0_100111101110;
      patterns[40677] = 29'b1_001111011100_101_0_010011110111;
      patterns[40678] = 29'b1_001111011100_110_1_001111011100;
      patterns[40679] = 29'b1_001111011100_111_1_001111011100;
      patterns[40680] = 29'b1_001111011101_000_1_001111011101;
      patterns[40681] = 29'b1_001111011101_001_1_011101001111;
      patterns[40682] = 29'b1_001111011101_010_0_011110111011;
      patterns[40683] = 29'b1_001111011101_011_0_111101110110;
      patterns[40684] = 29'b1_001111011101_100_1_100111101110;
      patterns[40685] = 29'b1_001111011101_101_0_110011110111;
      patterns[40686] = 29'b1_001111011101_110_1_001111011101;
      patterns[40687] = 29'b1_001111011101_111_1_001111011101;
      patterns[40688] = 29'b1_001111011110_000_1_001111011110;
      patterns[40689] = 29'b1_001111011110_001_1_011110001111;
      patterns[40690] = 29'b1_001111011110_010_0_011110111101;
      patterns[40691] = 29'b1_001111011110_011_0_111101111010;
      patterns[40692] = 29'b1_001111011110_100_0_100111101111;
      patterns[40693] = 29'b1_001111011110_101_1_010011110111;
      patterns[40694] = 29'b1_001111011110_110_1_001111011110;
      patterns[40695] = 29'b1_001111011110_111_1_001111011110;
      patterns[40696] = 29'b1_001111011111_000_1_001111011111;
      patterns[40697] = 29'b1_001111011111_001_1_011111001111;
      patterns[40698] = 29'b1_001111011111_010_0_011110111111;
      patterns[40699] = 29'b1_001111011111_011_0_111101111110;
      patterns[40700] = 29'b1_001111011111_100_1_100111101111;
      patterns[40701] = 29'b1_001111011111_101_1_110011110111;
      patterns[40702] = 29'b1_001111011111_110_1_001111011111;
      patterns[40703] = 29'b1_001111011111_111_1_001111011111;
      patterns[40704] = 29'b1_001111100000_000_1_001111100000;
      patterns[40705] = 29'b1_001111100000_001_1_100000001111;
      patterns[40706] = 29'b1_001111100000_010_0_011111000001;
      patterns[40707] = 29'b1_001111100000_011_0_111110000010;
      patterns[40708] = 29'b1_001111100000_100_0_100111110000;
      patterns[40709] = 29'b1_001111100000_101_0_010011111000;
      patterns[40710] = 29'b1_001111100000_110_1_001111100000;
      patterns[40711] = 29'b1_001111100000_111_1_001111100000;
      patterns[40712] = 29'b1_001111100001_000_1_001111100001;
      patterns[40713] = 29'b1_001111100001_001_1_100001001111;
      patterns[40714] = 29'b1_001111100001_010_0_011111000011;
      patterns[40715] = 29'b1_001111100001_011_0_111110000110;
      patterns[40716] = 29'b1_001111100001_100_1_100111110000;
      patterns[40717] = 29'b1_001111100001_101_0_110011111000;
      patterns[40718] = 29'b1_001111100001_110_1_001111100001;
      patterns[40719] = 29'b1_001111100001_111_1_001111100001;
      patterns[40720] = 29'b1_001111100010_000_1_001111100010;
      patterns[40721] = 29'b1_001111100010_001_1_100010001111;
      patterns[40722] = 29'b1_001111100010_010_0_011111000101;
      patterns[40723] = 29'b1_001111100010_011_0_111110001010;
      patterns[40724] = 29'b1_001111100010_100_0_100111110001;
      patterns[40725] = 29'b1_001111100010_101_1_010011111000;
      patterns[40726] = 29'b1_001111100010_110_1_001111100010;
      patterns[40727] = 29'b1_001111100010_111_1_001111100010;
      patterns[40728] = 29'b1_001111100011_000_1_001111100011;
      patterns[40729] = 29'b1_001111100011_001_1_100011001111;
      patterns[40730] = 29'b1_001111100011_010_0_011111000111;
      patterns[40731] = 29'b1_001111100011_011_0_111110001110;
      patterns[40732] = 29'b1_001111100011_100_1_100111110001;
      patterns[40733] = 29'b1_001111100011_101_1_110011111000;
      patterns[40734] = 29'b1_001111100011_110_1_001111100011;
      patterns[40735] = 29'b1_001111100011_111_1_001111100011;
      patterns[40736] = 29'b1_001111100100_000_1_001111100100;
      patterns[40737] = 29'b1_001111100100_001_1_100100001111;
      patterns[40738] = 29'b1_001111100100_010_0_011111001001;
      patterns[40739] = 29'b1_001111100100_011_0_111110010010;
      patterns[40740] = 29'b1_001111100100_100_0_100111110010;
      patterns[40741] = 29'b1_001111100100_101_0_010011111001;
      patterns[40742] = 29'b1_001111100100_110_1_001111100100;
      patterns[40743] = 29'b1_001111100100_111_1_001111100100;
      patterns[40744] = 29'b1_001111100101_000_1_001111100101;
      patterns[40745] = 29'b1_001111100101_001_1_100101001111;
      patterns[40746] = 29'b1_001111100101_010_0_011111001011;
      patterns[40747] = 29'b1_001111100101_011_0_111110010110;
      patterns[40748] = 29'b1_001111100101_100_1_100111110010;
      patterns[40749] = 29'b1_001111100101_101_0_110011111001;
      patterns[40750] = 29'b1_001111100101_110_1_001111100101;
      patterns[40751] = 29'b1_001111100101_111_1_001111100101;
      patterns[40752] = 29'b1_001111100110_000_1_001111100110;
      patterns[40753] = 29'b1_001111100110_001_1_100110001111;
      patterns[40754] = 29'b1_001111100110_010_0_011111001101;
      patterns[40755] = 29'b1_001111100110_011_0_111110011010;
      patterns[40756] = 29'b1_001111100110_100_0_100111110011;
      patterns[40757] = 29'b1_001111100110_101_1_010011111001;
      patterns[40758] = 29'b1_001111100110_110_1_001111100110;
      patterns[40759] = 29'b1_001111100110_111_1_001111100110;
      patterns[40760] = 29'b1_001111100111_000_1_001111100111;
      patterns[40761] = 29'b1_001111100111_001_1_100111001111;
      patterns[40762] = 29'b1_001111100111_010_0_011111001111;
      patterns[40763] = 29'b1_001111100111_011_0_111110011110;
      patterns[40764] = 29'b1_001111100111_100_1_100111110011;
      patterns[40765] = 29'b1_001111100111_101_1_110011111001;
      patterns[40766] = 29'b1_001111100111_110_1_001111100111;
      patterns[40767] = 29'b1_001111100111_111_1_001111100111;
      patterns[40768] = 29'b1_001111101000_000_1_001111101000;
      patterns[40769] = 29'b1_001111101000_001_1_101000001111;
      patterns[40770] = 29'b1_001111101000_010_0_011111010001;
      patterns[40771] = 29'b1_001111101000_011_0_111110100010;
      patterns[40772] = 29'b1_001111101000_100_0_100111110100;
      patterns[40773] = 29'b1_001111101000_101_0_010011111010;
      patterns[40774] = 29'b1_001111101000_110_1_001111101000;
      patterns[40775] = 29'b1_001111101000_111_1_001111101000;
      patterns[40776] = 29'b1_001111101001_000_1_001111101001;
      patterns[40777] = 29'b1_001111101001_001_1_101001001111;
      patterns[40778] = 29'b1_001111101001_010_0_011111010011;
      patterns[40779] = 29'b1_001111101001_011_0_111110100110;
      patterns[40780] = 29'b1_001111101001_100_1_100111110100;
      patterns[40781] = 29'b1_001111101001_101_0_110011111010;
      patterns[40782] = 29'b1_001111101001_110_1_001111101001;
      patterns[40783] = 29'b1_001111101001_111_1_001111101001;
      patterns[40784] = 29'b1_001111101010_000_1_001111101010;
      patterns[40785] = 29'b1_001111101010_001_1_101010001111;
      patterns[40786] = 29'b1_001111101010_010_0_011111010101;
      patterns[40787] = 29'b1_001111101010_011_0_111110101010;
      patterns[40788] = 29'b1_001111101010_100_0_100111110101;
      patterns[40789] = 29'b1_001111101010_101_1_010011111010;
      patterns[40790] = 29'b1_001111101010_110_1_001111101010;
      patterns[40791] = 29'b1_001111101010_111_1_001111101010;
      patterns[40792] = 29'b1_001111101011_000_1_001111101011;
      patterns[40793] = 29'b1_001111101011_001_1_101011001111;
      patterns[40794] = 29'b1_001111101011_010_0_011111010111;
      patterns[40795] = 29'b1_001111101011_011_0_111110101110;
      patterns[40796] = 29'b1_001111101011_100_1_100111110101;
      patterns[40797] = 29'b1_001111101011_101_1_110011111010;
      patterns[40798] = 29'b1_001111101011_110_1_001111101011;
      patterns[40799] = 29'b1_001111101011_111_1_001111101011;
      patterns[40800] = 29'b1_001111101100_000_1_001111101100;
      patterns[40801] = 29'b1_001111101100_001_1_101100001111;
      patterns[40802] = 29'b1_001111101100_010_0_011111011001;
      patterns[40803] = 29'b1_001111101100_011_0_111110110010;
      patterns[40804] = 29'b1_001111101100_100_0_100111110110;
      patterns[40805] = 29'b1_001111101100_101_0_010011111011;
      patterns[40806] = 29'b1_001111101100_110_1_001111101100;
      patterns[40807] = 29'b1_001111101100_111_1_001111101100;
      patterns[40808] = 29'b1_001111101101_000_1_001111101101;
      patterns[40809] = 29'b1_001111101101_001_1_101101001111;
      patterns[40810] = 29'b1_001111101101_010_0_011111011011;
      patterns[40811] = 29'b1_001111101101_011_0_111110110110;
      patterns[40812] = 29'b1_001111101101_100_1_100111110110;
      patterns[40813] = 29'b1_001111101101_101_0_110011111011;
      patterns[40814] = 29'b1_001111101101_110_1_001111101101;
      patterns[40815] = 29'b1_001111101101_111_1_001111101101;
      patterns[40816] = 29'b1_001111101110_000_1_001111101110;
      patterns[40817] = 29'b1_001111101110_001_1_101110001111;
      patterns[40818] = 29'b1_001111101110_010_0_011111011101;
      patterns[40819] = 29'b1_001111101110_011_0_111110111010;
      patterns[40820] = 29'b1_001111101110_100_0_100111110111;
      patterns[40821] = 29'b1_001111101110_101_1_010011111011;
      patterns[40822] = 29'b1_001111101110_110_1_001111101110;
      patterns[40823] = 29'b1_001111101110_111_1_001111101110;
      patterns[40824] = 29'b1_001111101111_000_1_001111101111;
      patterns[40825] = 29'b1_001111101111_001_1_101111001111;
      patterns[40826] = 29'b1_001111101111_010_0_011111011111;
      patterns[40827] = 29'b1_001111101111_011_0_111110111110;
      patterns[40828] = 29'b1_001111101111_100_1_100111110111;
      patterns[40829] = 29'b1_001111101111_101_1_110011111011;
      patterns[40830] = 29'b1_001111101111_110_1_001111101111;
      patterns[40831] = 29'b1_001111101111_111_1_001111101111;
      patterns[40832] = 29'b1_001111110000_000_1_001111110000;
      patterns[40833] = 29'b1_001111110000_001_1_110000001111;
      patterns[40834] = 29'b1_001111110000_010_0_011111100001;
      patterns[40835] = 29'b1_001111110000_011_0_111111000010;
      patterns[40836] = 29'b1_001111110000_100_0_100111111000;
      patterns[40837] = 29'b1_001111110000_101_0_010011111100;
      patterns[40838] = 29'b1_001111110000_110_1_001111110000;
      patterns[40839] = 29'b1_001111110000_111_1_001111110000;
      patterns[40840] = 29'b1_001111110001_000_1_001111110001;
      patterns[40841] = 29'b1_001111110001_001_1_110001001111;
      patterns[40842] = 29'b1_001111110001_010_0_011111100011;
      patterns[40843] = 29'b1_001111110001_011_0_111111000110;
      patterns[40844] = 29'b1_001111110001_100_1_100111111000;
      patterns[40845] = 29'b1_001111110001_101_0_110011111100;
      patterns[40846] = 29'b1_001111110001_110_1_001111110001;
      patterns[40847] = 29'b1_001111110001_111_1_001111110001;
      patterns[40848] = 29'b1_001111110010_000_1_001111110010;
      patterns[40849] = 29'b1_001111110010_001_1_110010001111;
      patterns[40850] = 29'b1_001111110010_010_0_011111100101;
      patterns[40851] = 29'b1_001111110010_011_0_111111001010;
      patterns[40852] = 29'b1_001111110010_100_0_100111111001;
      patterns[40853] = 29'b1_001111110010_101_1_010011111100;
      patterns[40854] = 29'b1_001111110010_110_1_001111110010;
      patterns[40855] = 29'b1_001111110010_111_1_001111110010;
      patterns[40856] = 29'b1_001111110011_000_1_001111110011;
      patterns[40857] = 29'b1_001111110011_001_1_110011001111;
      patterns[40858] = 29'b1_001111110011_010_0_011111100111;
      patterns[40859] = 29'b1_001111110011_011_0_111111001110;
      patterns[40860] = 29'b1_001111110011_100_1_100111111001;
      patterns[40861] = 29'b1_001111110011_101_1_110011111100;
      patterns[40862] = 29'b1_001111110011_110_1_001111110011;
      patterns[40863] = 29'b1_001111110011_111_1_001111110011;
      patterns[40864] = 29'b1_001111110100_000_1_001111110100;
      patterns[40865] = 29'b1_001111110100_001_1_110100001111;
      patterns[40866] = 29'b1_001111110100_010_0_011111101001;
      patterns[40867] = 29'b1_001111110100_011_0_111111010010;
      patterns[40868] = 29'b1_001111110100_100_0_100111111010;
      patterns[40869] = 29'b1_001111110100_101_0_010011111101;
      patterns[40870] = 29'b1_001111110100_110_1_001111110100;
      patterns[40871] = 29'b1_001111110100_111_1_001111110100;
      patterns[40872] = 29'b1_001111110101_000_1_001111110101;
      patterns[40873] = 29'b1_001111110101_001_1_110101001111;
      patterns[40874] = 29'b1_001111110101_010_0_011111101011;
      patterns[40875] = 29'b1_001111110101_011_0_111111010110;
      patterns[40876] = 29'b1_001111110101_100_1_100111111010;
      patterns[40877] = 29'b1_001111110101_101_0_110011111101;
      patterns[40878] = 29'b1_001111110101_110_1_001111110101;
      patterns[40879] = 29'b1_001111110101_111_1_001111110101;
      patterns[40880] = 29'b1_001111110110_000_1_001111110110;
      patterns[40881] = 29'b1_001111110110_001_1_110110001111;
      patterns[40882] = 29'b1_001111110110_010_0_011111101101;
      patterns[40883] = 29'b1_001111110110_011_0_111111011010;
      patterns[40884] = 29'b1_001111110110_100_0_100111111011;
      patterns[40885] = 29'b1_001111110110_101_1_010011111101;
      patterns[40886] = 29'b1_001111110110_110_1_001111110110;
      patterns[40887] = 29'b1_001111110110_111_1_001111110110;
      patterns[40888] = 29'b1_001111110111_000_1_001111110111;
      patterns[40889] = 29'b1_001111110111_001_1_110111001111;
      patterns[40890] = 29'b1_001111110111_010_0_011111101111;
      patterns[40891] = 29'b1_001111110111_011_0_111111011110;
      patterns[40892] = 29'b1_001111110111_100_1_100111111011;
      patterns[40893] = 29'b1_001111110111_101_1_110011111101;
      patterns[40894] = 29'b1_001111110111_110_1_001111110111;
      patterns[40895] = 29'b1_001111110111_111_1_001111110111;
      patterns[40896] = 29'b1_001111111000_000_1_001111111000;
      patterns[40897] = 29'b1_001111111000_001_1_111000001111;
      patterns[40898] = 29'b1_001111111000_010_0_011111110001;
      patterns[40899] = 29'b1_001111111000_011_0_111111100010;
      patterns[40900] = 29'b1_001111111000_100_0_100111111100;
      patterns[40901] = 29'b1_001111111000_101_0_010011111110;
      patterns[40902] = 29'b1_001111111000_110_1_001111111000;
      patterns[40903] = 29'b1_001111111000_111_1_001111111000;
      patterns[40904] = 29'b1_001111111001_000_1_001111111001;
      patterns[40905] = 29'b1_001111111001_001_1_111001001111;
      patterns[40906] = 29'b1_001111111001_010_0_011111110011;
      patterns[40907] = 29'b1_001111111001_011_0_111111100110;
      patterns[40908] = 29'b1_001111111001_100_1_100111111100;
      patterns[40909] = 29'b1_001111111001_101_0_110011111110;
      patterns[40910] = 29'b1_001111111001_110_1_001111111001;
      patterns[40911] = 29'b1_001111111001_111_1_001111111001;
      patterns[40912] = 29'b1_001111111010_000_1_001111111010;
      patterns[40913] = 29'b1_001111111010_001_1_111010001111;
      patterns[40914] = 29'b1_001111111010_010_0_011111110101;
      patterns[40915] = 29'b1_001111111010_011_0_111111101010;
      patterns[40916] = 29'b1_001111111010_100_0_100111111101;
      patterns[40917] = 29'b1_001111111010_101_1_010011111110;
      patterns[40918] = 29'b1_001111111010_110_1_001111111010;
      patterns[40919] = 29'b1_001111111010_111_1_001111111010;
      patterns[40920] = 29'b1_001111111011_000_1_001111111011;
      patterns[40921] = 29'b1_001111111011_001_1_111011001111;
      patterns[40922] = 29'b1_001111111011_010_0_011111110111;
      patterns[40923] = 29'b1_001111111011_011_0_111111101110;
      patterns[40924] = 29'b1_001111111011_100_1_100111111101;
      patterns[40925] = 29'b1_001111111011_101_1_110011111110;
      patterns[40926] = 29'b1_001111111011_110_1_001111111011;
      patterns[40927] = 29'b1_001111111011_111_1_001111111011;
      patterns[40928] = 29'b1_001111111100_000_1_001111111100;
      patterns[40929] = 29'b1_001111111100_001_1_111100001111;
      patterns[40930] = 29'b1_001111111100_010_0_011111111001;
      patterns[40931] = 29'b1_001111111100_011_0_111111110010;
      patterns[40932] = 29'b1_001111111100_100_0_100111111110;
      patterns[40933] = 29'b1_001111111100_101_0_010011111111;
      patterns[40934] = 29'b1_001111111100_110_1_001111111100;
      patterns[40935] = 29'b1_001111111100_111_1_001111111100;
      patterns[40936] = 29'b1_001111111101_000_1_001111111101;
      patterns[40937] = 29'b1_001111111101_001_1_111101001111;
      patterns[40938] = 29'b1_001111111101_010_0_011111111011;
      patterns[40939] = 29'b1_001111111101_011_0_111111110110;
      patterns[40940] = 29'b1_001111111101_100_1_100111111110;
      patterns[40941] = 29'b1_001111111101_101_0_110011111111;
      patterns[40942] = 29'b1_001111111101_110_1_001111111101;
      patterns[40943] = 29'b1_001111111101_111_1_001111111101;
      patterns[40944] = 29'b1_001111111110_000_1_001111111110;
      patterns[40945] = 29'b1_001111111110_001_1_111110001111;
      patterns[40946] = 29'b1_001111111110_010_0_011111111101;
      patterns[40947] = 29'b1_001111111110_011_0_111111111010;
      patterns[40948] = 29'b1_001111111110_100_0_100111111111;
      patterns[40949] = 29'b1_001111111110_101_1_010011111111;
      patterns[40950] = 29'b1_001111111110_110_1_001111111110;
      patterns[40951] = 29'b1_001111111110_111_1_001111111110;
      patterns[40952] = 29'b1_001111111111_000_1_001111111111;
      patterns[40953] = 29'b1_001111111111_001_1_111111001111;
      patterns[40954] = 29'b1_001111111111_010_0_011111111111;
      patterns[40955] = 29'b1_001111111111_011_0_111111111110;
      patterns[40956] = 29'b1_001111111111_100_1_100111111111;
      patterns[40957] = 29'b1_001111111111_101_1_110011111111;
      patterns[40958] = 29'b1_001111111111_110_1_001111111111;
      patterns[40959] = 29'b1_001111111111_111_1_001111111111;
      patterns[40960] = 29'b1_010000000000_000_1_010000000000;
      patterns[40961] = 29'b1_010000000000_001_1_000000010000;
      patterns[40962] = 29'b1_010000000000_010_0_100000000001;
      patterns[40963] = 29'b1_010000000000_011_1_000000000010;
      patterns[40964] = 29'b1_010000000000_100_0_101000000000;
      patterns[40965] = 29'b1_010000000000_101_0_010100000000;
      patterns[40966] = 29'b1_010000000000_110_1_010000000000;
      patterns[40967] = 29'b1_010000000000_111_1_010000000000;
      patterns[40968] = 29'b1_010000000001_000_1_010000000001;
      patterns[40969] = 29'b1_010000000001_001_1_000001010000;
      patterns[40970] = 29'b1_010000000001_010_0_100000000011;
      patterns[40971] = 29'b1_010000000001_011_1_000000000110;
      patterns[40972] = 29'b1_010000000001_100_1_101000000000;
      patterns[40973] = 29'b1_010000000001_101_0_110100000000;
      patterns[40974] = 29'b1_010000000001_110_1_010000000001;
      patterns[40975] = 29'b1_010000000001_111_1_010000000001;
      patterns[40976] = 29'b1_010000000010_000_1_010000000010;
      patterns[40977] = 29'b1_010000000010_001_1_000010010000;
      patterns[40978] = 29'b1_010000000010_010_0_100000000101;
      patterns[40979] = 29'b1_010000000010_011_1_000000001010;
      patterns[40980] = 29'b1_010000000010_100_0_101000000001;
      patterns[40981] = 29'b1_010000000010_101_1_010100000000;
      patterns[40982] = 29'b1_010000000010_110_1_010000000010;
      patterns[40983] = 29'b1_010000000010_111_1_010000000010;
      patterns[40984] = 29'b1_010000000011_000_1_010000000011;
      patterns[40985] = 29'b1_010000000011_001_1_000011010000;
      patterns[40986] = 29'b1_010000000011_010_0_100000000111;
      patterns[40987] = 29'b1_010000000011_011_1_000000001110;
      patterns[40988] = 29'b1_010000000011_100_1_101000000001;
      patterns[40989] = 29'b1_010000000011_101_1_110100000000;
      patterns[40990] = 29'b1_010000000011_110_1_010000000011;
      patterns[40991] = 29'b1_010000000011_111_1_010000000011;
      patterns[40992] = 29'b1_010000000100_000_1_010000000100;
      patterns[40993] = 29'b1_010000000100_001_1_000100010000;
      patterns[40994] = 29'b1_010000000100_010_0_100000001001;
      patterns[40995] = 29'b1_010000000100_011_1_000000010010;
      patterns[40996] = 29'b1_010000000100_100_0_101000000010;
      patterns[40997] = 29'b1_010000000100_101_0_010100000001;
      patterns[40998] = 29'b1_010000000100_110_1_010000000100;
      patterns[40999] = 29'b1_010000000100_111_1_010000000100;
      patterns[41000] = 29'b1_010000000101_000_1_010000000101;
      patterns[41001] = 29'b1_010000000101_001_1_000101010000;
      patterns[41002] = 29'b1_010000000101_010_0_100000001011;
      patterns[41003] = 29'b1_010000000101_011_1_000000010110;
      patterns[41004] = 29'b1_010000000101_100_1_101000000010;
      patterns[41005] = 29'b1_010000000101_101_0_110100000001;
      patterns[41006] = 29'b1_010000000101_110_1_010000000101;
      patterns[41007] = 29'b1_010000000101_111_1_010000000101;
      patterns[41008] = 29'b1_010000000110_000_1_010000000110;
      patterns[41009] = 29'b1_010000000110_001_1_000110010000;
      patterns[41010] = 29'b1_010000000110_010_0_100000001101;
      patterns[41011] = 29'b1_010000000110_011_1_000000011010;
      patterns[41012] = 29'b1_010000000110_100_0_101000000011;
      patterns[41013] = 29'b1_010000000110_101_1_010100000001;
      patterns[41014] = 29'b1_010000000110_110_1_010000000110;
      patterns[41015] = 29'b1_010000000110_111_1_010000000110;
      patterns[41016] = 29'b1_010000000111_000_1_010000000111;
      patterns[41017] = 29'b1_010000000111_001_1_000111010000;
      patterns[41018] = 29'b1_010000000111_010_0_100000001111;
      patterns[41019] = 29'b1_010000000111_011_1_000000011110;
      patterns[41020] = 29'b1_010000000111_100_1_101000000011;
      patterns[41021] = 29'b1_010000000111_101_1_110100000001;
      patterns[41022] = 29'b1_010000000111_110_1_010000000111;
      patterns[41023] = 29'b1_010000000111_111_1_010000000111;
      patterns[41024] = 29'b1_010000001000_000_1_010000001000;
      patterns[41025] = 29'b1_010000001000_001_1_001000010000;
      patterns[41026] = 29'b1_010000001000_010_0_100000010001;
      patterns[41027] = 29'b1_010000001000_011_1_000000100010;
      patterns[41028] = 29'b1_010000001000_100_0_101000000100;
      patterns[41029] = 29'b1_010000001000_101_0_010100000010;
      patterns[41030] = 29'b1_010000001000_110_1_010000001000;
      patterns[41031] = 29'b1_010000001000_111_1_010000001000;
      patterns[41032] = 29'b1_010000001001_000_1_010000001001;
      patterns[41033] = 29'b1_010000001001_001_1_001001010000;
      patterns[41034] = 29'b1_010000001001_010_0_100000010011;
      patterns[41035] = 29'b1_010000001001_011_1_000000100110;
      patterns[41036] = 29'b1_010000001001_100_1_101000000100;
      patterns[41037] = 29'b1_010000001001_101_0_110100000010;
      patterns[41038] = 29'b1_010000001001_110_1_010000001001;
      patterns[41039] = 29'b1_010000001001_111_1_010000001001;
      patterns[41040] = 29'b1_010000001010_000_1_010000001010;
      patterns[41041] = 29'b1_010000001010_001_1_001010010000;
      patterns[41042] = 29'b1_010000001010_010_0_100000010101;
      patterns[41043] = 29'b1_010000001010_011_1_000000101010;
      patterns[41044] = 29'b1_010000001010_100_0_101000000101;
      patterns[41045] = 29'b1_010000001010_101_1_010100000010;
      patterns[41046] = 29'b1_010000001010_110_1_010000001010;
      patterns[41047] = 29'b1_010000001010_111_1_010000001010;
      patterns[41048] = 29'b1_010000001011_000_1_010000001011;
      patterns[41049] = 29'b1_010000001011_001_1_001011010000;
      patterns[41050] = 29'b1_010000001011_010_0_100000010111;
      patterns[41051] = 29'b1_010000001011_011_1_000000101110;
      patterns[41052] = 29'b1_010000001011_100_1_101000000101;
      patterns[41053] = 29'b1_010000001011_101_1_110100000010;
      patterns[41054] = 29'b1_010000001011_110_1_010000001011;
      patterns[41055] = 29'b1_010000001011_111_1_010000001011;
      patterns[41056] = 29'b1_010000001100_000_1_010000001100;
      patterns[41057] = 29'b1_010000001100_001_1_001100010000;
      patterns[41058] = 29'b1_010000001100_010_0_100000011001;
      patterns[41059] = 29'b1_010000001100_011_1_000000110010;
      patterns[41060] = 29'b1_010000001100_100_0_101000000110;
      patterns[41061] = 29'b1_010000001100_101_0_010100000011;
      patterns[41062] = 29'b1_010000001100_110_1_010000001100;
      patterns[41063] = 29'b1_010000001100_111_1_010000001100;
      patterns[41064] = 29'b1_010000001101_000_1_010000001101;
      patterns[41065] = 29'b1_010000001101_001_1_001101010000;
      patterns[41066] = 29'b1_010000001101_010_0_100000011011;
      patterns[41067] = 29'b1_010000001101_011_1_000000110110;
      patterns[41068] = 29'b1_010000001101_100_1_101000000110;
      patterns[41069] = 29'b1_010000001101_101_0_110100000011;
      patterns[41070] = 29'b1_010000001101_110_1_010000001101;
      patterns[41071] = 29'b1_010000001101_111_1_010000001101;
      patterns[41072] = 29'b1_010000001110_000_1_010000001110;
      patterns[41073] = 29'b1_010000001110_001_1_001110010000;
      patterns[41074] = 29'b1_010000001110_010_0_100000011101;
      patterns[41075] = 29'b1_010000001110_011_1_000000111010;
      patterns[41076] = 29'b1_010000001110_100_0_101000000111;
      patterns[41077] = 29'b1_010000001110_101_1_010100000011;
      patterns[41078] = 29'b1_010000001110_110_1_010000001110;
      patterns[41079] = 29'b1_010000001110_111_1_010000001110;
      patterns[41080] = 29'b1_010000001111_000_1_010000001111;
      patterns[41081] = 29'b1_010000001111_001_1_001111010000;
      patterns[41082] = 29'b1_010000001111_010_0_100000011111;
      patterns[41083] = 29'b1_010000001111_011_1_000000111110;
      patterns[41084] = 29'b1_010000001111_100_1_101000000111;
      patterns[41085] = 29'b1_010000001111_101_1_110100000011;
      patterns[41086] = 29'b1_010000001111_110_1_010000001111;
      patterns[41087] = 29'b1_010000001111_111_1_010000001111;
      patterns[41088] = 29'b1_010000010000_000_1_010000010000;
      patterns[41089] = 29'b1_010000010000_001_1_010000010000;
      patterns[41090] = 29'b1_010000010000_010_0_100000100001;
      patterns[41091] = 29'b1_010000010000_011_1_000001000010;
      patterns[41092] = 29'b1_010000010000_100_0_101000001000;
      patterns[41093] = 29'b1_010000010000_101_0_010100000100;
      patterns[41094] = 29'b1_010000010000_110_1_010000010000;
      patterns[41095] = 29'b1_010000010000_111_1_010000010000;
      patterns[41096] = 29'b1_010000010001_000_1_010000010001;
      patterns[41097] = 29'b1_010000010001_001_1_010001010000;
      patterns[41098] = 29'b1_010000010001_010_0_100000100011;
      patterns[41099] = 29'b1_010000010001_011_1_000001000110;
      patterns[41100] = 29'b1_010000010001_100_1_101000001000;
      patterns[41101] = 29'b1_010000010001_101_0_110100000100;
      patterns[41102] = 29'b1_010000010001_110_1_010000010001;
      patterns[41103] = 29'b1_010000010001_111_1_010000010001;
      patterns[41104] = 29'b1_010000010010_000_1_010000010010;
      patterns[41105] = 29'b1_010000010010_001_1_010010010000;
      patterns[41106] = 29'b1_010000010010_010_0_100000100101;
      patterns[41107] = 29'b1_010000010010_011_1_000001001010;
      patterns[41108] = 29'b1_010000010010_100_0_101000001001;
      patterns[41109] = 29'b1_010000010010_101_1_010100000100;
      patterns[41110] = 29'b1_010000010010_110_1_010000010010;
      patterns[41111] = 29'b1_010000010010_111_1_010000010010;
      patterns[41112] = 29'b1_010000010011_000_1_010000010011;
      patterns[41113] = 29'b1_010000010011_001_1_010011010000;
      patterns[41114] = 29'b1_010000010011_010_0_100000100111;
      patterns[41115] = 29'b1_010000010011_011_1_000001001110;
      patterns[41116] = 29'b1_010000010011_100_1_101000001001;
      patterns[41117] = 29'b1_010000010011_101_1_110100000100;
      patterns[41118] = 29'b1_010000010011_110_1_010000010011;
      patterns[41119] = 29'b1_010000010011_111_1_010000010011;
      patterns[41120] = 29'b1_010000010100_000_1_010000010100;
      patterns[41121] = 29'b1_010000010100_001_1_010100010000;
      patterns[41122] = 29'b1_010000010100_010_0_100000101001;
      patterns[41123] = 29'b1_010000010100_011_1_000001010010;
      patterns[41124] = 29'b1_010000010100_100_0_101000001010;
      patterns[41125] = 29'b1_010000010100_101_0_010100000101;
      patterns[41126] = 29'b1_010000010100_110_1_010000010100;
      patterns[41127] = 29'b1_010000010100_111_1_010000010100;
      patterns[41128] = 29'b1_010000010101_000_1_010000010101;
      patterns[41129] = 29'b1_010000010101_001_1_010101010000;
      patterns[41130] = 29'b1_010000010101_010_0_100000101011;
      patterns[41131] = 29'b1_010000010101_011_1_000001010110;
      patterns[41132] = 29'b1_010000010101_100_1_101000001010;
      patterns[41133] = 29'b1_010000010101_101_0_110100000101;
      patterns[41134] = 29'b1_010000010101_110_1_010000010101;
      patterns[41135] = 29'b1_010000010101_111_1_010000010101;
      patterns[41136] = 29'b1_010000010110_000_1_010000010110;
      patterns[41137] = 29'b1_010000010110_001_1_010110010000;
      patterns[41138] = 29'b1_010000010110_010_0_100000101101;
      patterns[41139] = 29'b1_010000010110_011_1_000001011010;
      patterns[41140] = 29'b1_010000010110_100_0_101000001011;
      patterns[41141] = 29'b1_010000010110_101_1_010100000101;
      patterns[41142] = 29'b1_010000010110_110_1_010000010110;
      patterns[41143] = 29'b1_010000010110_111_1_010000010110;
      patterns[41144] = 29'b1_010000010111_000_1_010000010111;
      patterns[41145] = 29'b1_010000010111_001_1_010111010000;
      patterns[41146] = 29'b1_010000010111_010_0_100000101111;
      patterns[41147] = 29'b1_010000010111_011_1_000001011110;
      patterns[41148] = 29'b1_010000010111_100_1_101000001011;
      patterns[41149] = 29'b1_010000010111_101_1_110100000101;
      patterns[41150] = 29'b1_010000010111_110_1_010000010111;
      patterns[41151] = 29'b1_010000010111_111_1_010000010111;
      patterns[41152] = 29'b1_010000011000_000_1_010000011000;
      patterns[41153] = 29'b1_010000011000_001_1_011000010000;
      patterns[41154] = 29'b1_010000011000_010_0_100000110001;
      patterns[41155] = 29'b1_010000011000_011_1_000001100010;
      patterns[41156] = 29'b1_010000011000_100_0_101000001100;
      patterns[41157] = 29'b1_010000011000_101_0_010100000110;
      patterns[41158] = 29'b1_010000011000_110_1_010000011000;
      patterns[41159] = 29'b1_010000011000_111_1_010000011000;
      patterns[41160] = 29'b1_010000011001_000_1_010000011001;
      patterns[41161] = 29'b1_010000011001_001_1_011001010000;
      patterns[41162] = 29'b1_010000011001_010_0_100000110011;
      patterns[41163] = 29'b1_010000011001_011_1_000001100110;
      patterns[41164] = 29'b1_010000011001_100_1_101000001100;
      patterns[41165] = 29'b1_010000011001_101_0_110100000110;
      patterns[41166] = 29'b1_010000011001_110_1_010000011001;
      patterns[41167] = 29'b1_010000011001_111_1_010000011001;
      patterns[41168] = 29'b1_010000011010_000_1_010000011010;
      patterns[41169] = 29'b1_010000011010_001_1_011010010000;
      patterns[41170] = 29'b1_010000011010_010_0_100000110101;
      patterns[41171] = 29'b1_010000011010_011_1_000001101010;
      patterns[41172] = 29'b1_010000011010_100_0_101000001101;
      patterns[41173] = 29'b1_010000011010_101_1_010100000110;
      patterns[41174] = 29'b1_010000011010_110_1_010000011010;
      patterns[41175] = 29'b1_010000011010_111_1_010000011010;
      patterns[41176] = 29'b1_010000011011_000_1_010000011011;
      patterns[41177] = 29'b1_010000011011_001_1_011011010000;
      patterns[41178] = 29'b1_010000011011_010_0_100000110111;
      patterns[41179] = 29'b1_010000011011_011_1_000001101110;
      patterns[41180] = 29'b1_010000011011_100_1_101000001101;
      patterns[41181] = 29'b1_010000011011_101_1_110100000110;
      patterns[41182] = 29'b1_010000011011_110_1_010000011011;
      patterns[41183] = 29'b1_010000011011_111_1_010000011011;
      patterns[41184] = 29'b1_010000011100_000_1_010000011100;
      patterns[41185] = 29'b1_010000011100_001_1_011100010000;
      patterns[41186] = 29'b1_010000011100_010_0_100000111001;
      patterns[41187] = 29'b1_010000011100_011_1_000001110010;
      patterns[41188] = 29'b1_010000011100_100_0_101000001110;
      patterns[41189] = 29'b1_010000011100_101_0_010100000111;
      patterns[41190] = 29'b1_010000011100_110_1_010000011100;
      patterns[41191] = 29'b1_010000011100_111_1_010000011100;
      patterns[41192] = 29'b1_010000011101_000_1_010000011101;
      patterns[41193] = 29'b1_010000011101_001_1_011101010000;
      patterns[41194] = 29'b1_010000011101_010_0_100000111011;
      patterns[41195] = 29'b1_010000011101_011_1_000001110110;
      patterns[41196] = 29'b1_010000011101_100_1_101000001110;
      patterns[41197] = 29'b1_010000011101_101_0_110100000111;
      patterns[41198] = 29'b1_010000011101_110_1_010000011101;
      patterns[41199] = 29'b1_010000011101_111_1_010000011101;
      patterns[41200] = 29'b1_010000011110_000_1_010000011110;
      patterns[41201] = 29'b1_010000011110_001_1_011110010000;
      patterns[41202] = 29'b1_010000011110_010_0_100000111101;
      patterns[41203] = 29'b1_010000011110_011_1_000001111010;
      patterns[41204] = 29'b1_010000011110_100_0_101000001111;
      patterns[41205] = 29'b1_010000011110_101_1_010100000111;
      patterns[41206] = 29'b1_010000011110_110_1_010000011110;
      patterns[41207] = 29'b1_010000011110_111_1_010000011110;
      patterns[41208] = 29'b1_010000011111_000_1_010000011111;
      patterns[41209] = 29'b1_010000011111_001_1_011111010000;
      patterns[41210] = 29'b1_010000011111_010_0_100000111111;
      patterns[41211] = 29'b1_010000011111_011_1_000001111110;
      patterns[41212] = 29'b1_010000011111_100_1_101000001111;
      patterns[41213] = 29'b1_010000011111_101_1_110100000111;
      patterns[41214] = 29'b1_010000011111_110_1_010000011111;
      patterns[41215] = 29'b1_010000011111_111_1_010000011111;
      patterns[41216] = 29'b1_010000100000_000_1_010000100000;
      patterns[41217] = 29'b1_010000100000_001_1_100000010000;
      patterns[41218] = 29'b1_010000100000_010_0_100001000001;
      patterns[41219] = 29'b1_010000100000_011_1_000010000010;
      patterns[41220] = 29'b1_010000100000_100_0_101000010000;
      patterns[41221] = 29'b1_010000100000_101_0_010100001000;
      patterns[41222] = 29'b1_010000100000_110_1_010000100000;
      patterns[41223] = 29'b1_010000100000_111_1_010000100000;
      patterns[41224] = 29'b1_010000100001_000_1_010000100001;
      patterns[41225] = 29'b1_010000100001_001_1_100001010000;
      patterns[41226] = 29'b1_010000100001_010_0_100001000011;
      patterns[41227] = 29'b1_010000100001_011_1_000010000110;
      patterns[41228] = 29'b1_010000100001_100_1_101000010000;
      patterns[41229] = 29'b1_010000100001_101_0_110100001000;
      patterns[41230] = 29'b1_010000100001_110_1_010000100001;
      patterns[41231] = 29'b1_010000100001_111_1_010000100001;
      patterns[41232] = 29'b1_010000100010_000_1_010000100010;
      patterns[41233] = 29'b1_010000100010_001_1_100010010000;
      patterns[41234] = 29'b1_010000100010_010_0_100001000101;
      patterns[41235] = 29'b1_010000100010_011_1_000010001010;
      patterns[41236] = 29'b1_010000100010_100_0_101000010001;
      patterns[41237] = 29'b1_010000100010_101_1_010100001000;
      patterns[41238] = 29'b1_010000100010_110_1_010000100010;
      patterns[41239] = 29'b1_010000100010_111_1_010000100010;
      patterns[41240] = 29'b1_010000100011_000_1_010000100011;
      patterns[41241] = 29'b1_010000100011_001_1_100011010000;
      patterns[41242] = 29'b1_010000100011_010_0_100001000111;
      patterns[41243] = 29'b1_010000100011_011_1_000010001110;
      patterns[41244] = 29'b1_010000100011_100_1_101000010001;
      patterns[41245] = 29'b1_010000100011_101_1_110100001000;
      patterns[41246] = 29'b1_010000100011_110_1_010000100011;
      patterns[41247] = 29'b1_010000100011_111_1_010000100011;
      patterns[41248] = 29'b1_010000100100_000_1_010000100100;
      patterns[41249] = 29'b1_010000100100_001_1_100100010000;
      patterns[41250] = 29'b1_010000100100_010_0_100001001001;
      patterns[41251] = 29'b1_010000100100_011_1_000010010010;
      patterns[41252] = 29'b1_010000100100_100_0_101000010010;
      patterns[41253] = 29'b1_010000100100_101_0_010100001001;
      patterns[41254] = 29'b1_010000100100_110_1_010000100100;
      patterns[41255] = 29'b1_010000100100_111_1_010000100100;
      patterns[41256] = 29'b1_010000100101_000_1_010000100101;
      patterns[41257] = 29'b1_010000100101_001_1_100101010000;
      patterns[41258] = 29'b1_010000100101_010_0_100001001011;
      patterns[41259] = 29'b1_010000100101_011_1_000010010110;
      patterns[41260] = 29'b1_010000100101_100_1_101000010010;
      patterns[41261] = 29'b1_010000100101_101_0_110100001001;
      patterns[41262] = 29'b1_010000100101_110_1_010000100101;
      patterns[41263] = 29'b1_010000100101_111_1_010000100101;
      patterns[41264] = 29'b1_010000100110_000_1_010000100110;
      patterns[41265] = 29'b1_010000100110_001_1_100110010000;
      patterns[41266] = 29'b1_010000100110_010_0_100001001101;
      patterns[41267] = 29'b1_010000100110_011_1_000010011010;
      patterns[41268] = 29'b1_010000100110_100_0_101000010011;
      patterns[41269] = 29'b1_010000100110_101_1_010100001001;
      patterns[41270] = 29'b1_010000100110_110_1_010000100110;
      patterns[41271] = 29'b1_010000100110_111_1_010000100110;
      patterns[41272] = 29'b1_010000100111_000_1_010000100111;
      patterns[41273] = 29'b1_010000100111_001_1_100111010000;
      patterns[41274] = 29'b1_010000100111_010_0_100001001111;
      patterns[41275] = 29'b1_010000100111_011_1_000010011110;
      patterns[41276] = 29'b1_010000100111_100_1_101000010011;
      patterns[41277] = 29'b1_010000100111_101_1_110100001001;
      patterns[41278] = 29'b1_010000100111_110_1_010000100111;
      patterns[41279] = 29'b1_010000100111_111_1_010000100111;
      patterns[41280] = 29'b1_010000101000_000_1_010000101000;
      patterns[41281] = 29'b1_010000101000_001_1_101000010000;
      patterns[41282] = 29'b1_010000101000_010_0_100001010001;
      patterns[41283] = 29'b1_010000101000_011_1_000010100010;
      patterns[41284] = 29'b1_010000101000_100_0_101000010100;
      patterns[41285] = 29'b1_010000101000_101_0_010100001010;
      patterns[41286] = 29'b1_010000101000_110_1_010000101000;
      patterns[41287] = 29'b1_010000101000_111_1_010000101000;
      patterns[41288] = 29'b1_010000101001_000_1_010000101001;
      patterns[41289] = 29'b1_010000101001_001_1_101001010000;
      patterns[41290] = 29'b1_010000101001_010_0_100001010011;
      patterns[41291] = 29'b1_010000101001_011_1_000010100110;
      patterns[41292] = 29'b1_010000101001_100_1_101000010100;
      patterns[41293] = 29'b1_010000101001_101_0_110100001010;
      patterns[41294] = 29'b1_010000101001_110_1_010000101001;
      patterns[41295] = 29'b1_010000101001_111_1_010000101001;
      patterns[41296] = 29'b1_010000101010_000_1_010000101010;
      patterns[41297] = 29'b1_010000101010_001_1_101010010000;
      patterns[41298] = 29'b1_010000101010_010_0_100001010101;
      patterns[41299] = 29'b1_010000101010_011_1_000010101010;
      patterns[41300] = 29'b1_010000101010_100_0_101000010101;
      patterns[41301] = 29'b1_010000101010_101_1_010100001010;
      patterns[41302] = 29'b1_010000101010_110_1_010000101010;
      patterns[41303] = 29'b1_010000101010_111_1_010000101010;
      patterns[41304] = 29'b1_010000101011_000_1_010000101011;
      patterns[41305] = 29'b1_010000101011_001_1_101011010000;
      patterns[41306] = 29'b1_010000101011_010_0_100001010111;
      patterns[41307] = 29'b1_010000101011_011_1_000010101110;
      patterns[41308] = 29'b1_010000101011_100_1_101000010101;
      patterns[41309] = 29'b1_010000101011_101_1_110100001010;
      patterns[41310] = 29'b1_010000101011_110_1_010000101011;
      patterns[41311] = 29'b1_010000101011_111_1_010000101011;
      patterns[41312] = 29'b1_010000101100_000_1_010000101100;
      patterns[41313] = 29'b1_010000101100_001_1_101100010000;
      patterns[41314] = 29'b1_010000101100_010_0_100001011001;
      patterns[41315] = 29'b1_010000101100_011_1_000010110010;
      patterns[41316] = 29'b1_010000101100_100_0_101000010110;
      patterns[41317] = 29'b1_010000101100_101_0_010100001011;
      patterns[41318] = 29'b1_010000101100_110_1_010000101100;
      patterns[41319] = 29'b1_010000101100_111_1_010000101100;
      patterns[41320] = 29'b1_010000101101_000_1_010000101101;
      patterns[41321] = 29'b1_010000101101_001_1_101101010000;
      patterns[41322] = 29'b1_010000101101_010_0_100001011011;
      patterns[41323] = 29'b1_010000101101_011_1_000010110110;
      patterns[41324] = 29'b1_010000101101_100_1_101000010110;
      patterns[41325] = 29'b1_010000101101_101_0_110100001011;
      patterns[41326] = 29'b1_010000101101_110_1_010000101101;
      patterns[41327] = 29'b1_010000101101_111_1_010000101101;
      patterns[41328] = 29'b1_010000101110_000_1_010000101110;
      patterns[41329] = 29'b1_010000101110_001_1_101110010000;
      patterns[41330] = 29'b1_010000101110_010_0_100001011101;
      patterns[41331] = 29'b1_010000101110_011_1_000010111010;
      patterns[41332] = 29'b1_010000101110_100_0_101000010111;
      patterns[41333] = 29'b1_010000101110_101_1_010100001011;
      patterns[41334] = 29'b1_010000101110_110_1_010000101110;
      patterns[41335] = 29'b1_010000101110_111_1_010000101110;
      patterns[41336] = 29'b1_010000101111_000_1_010000101111;
      patterns[41337] = 29'b1_010000101111_001_1_101111010000;
      patterns[41338] = 29'b1_010000101111_010_0_100001011111;
      patterns[41339] = 29'b1_010000101111_011_1_000010111110;
      patterns[41340] = 29'b1_010000101111_100_1_101000010111;
      patterns[41341] = 29'b1_010000101111_101_1_110100001011;
      patterns[41342] = 29'b1_010000101111_110_1_010000101111;
      patterns[41343] = 29'b1_010000101111_111_1_010000101111;
      patterns[41344] = 29'b1_010000110000_000_1_010000110000;
      patterns[41345] = 29'b1_010000110000_001_1_110000010000;
      patterns[41346] = 29'b1_010000110000_010_0_100001100001;
      patterns[41347] = 29'b1_010000110000_011_1_000011000010;
      patterns[41348] = 29'b1_010000110000_100_0_101000011000;
      patterns[41349] = 29'b1_010000110000_101_0_010100001100;
      patterns[41350] = 29'b1_010000110000_110_1_010000110000;
      patterns[41351] = 29'b1_010000110000_111_1_010000110000;
      patterns[41352] = 29'b1_010000110001_000_1_010000110001;
      patterns[41353] = 29'b1_010000110001_001_1_110001010000;
      patterns[41354] = 29'b1_010000110001_010_0_100001100011;
      patterns[41355] = 29'b1_010000110001_011_1_000011000110;
      patterns[41356] = 29'b1_010000110001_100_1_101000011000;
      patterns[41357] = 29'b1_010000110001_101_0_110100001100;
      patterns[41358] = 29'b1_010000110001_110_1_010000110001;
      patterns[41359] = 29'b1_010000110001_111_1_010000110001;
      patterns[41360] = 29'b1_010000110010_000_1_010000110010;
      patterns[41361] = 29'b1_010000110010_001_1_110010010000;
      patterns[41362] = 29'b1_010000110010_010_0_100001100101;
      patterns[41363] = 29'b1_010000110010_011_1_000011001010;
      patterns[41364] = 29'b1_010000110010_100_0_101000011001;
      patterns[41365] = 29'b1_010000110010_101_1_010100001100;
      patterns[41366] = 29'b1_010000110010_110_1_010000110010;
      patterns[41367] = 29'b1_010000110010_111_1_010000110010;
      patterns[41368] = 29'b1_010000110011_000_1_010000110011;
      patterns[41369] = 29'b1_010000110011_001_1_110011010000;
      patterns[41370] = 29'b1_010000110011_010_0_100001100111;
      patterns[41371] = 29'b1_010000110011_011_1_000011001110;
      patterns[41372] = 29'b1_010000110011_100_1_101000011001;
      patterns[41373] = 29'b1_010000110011_101_1_110100001100;
      patterns[41374] = 29'b1_010000110011_110_1_010000110011;
      patterns[41375] = 29'b1_010000110011_111_1_010000110011;
      patterns[41376] = 29'b1_010000110100_000_1_010000110100;
      patterns[41377] = 29'b1_010000110100_001_1_110100010000;
      patterns[41378] = 29'b1_010000110100_010_0_100001101001;
      patterns[41379] = 29'b1_010000110100_011_1_000011010010;
      patterns[41380] = 29'b1_010000110100_100_0_101000011010;
      patterns[41381] = 29'b1_010000110100_101_0_010100001101;
      patterns[41382] = 29'b1_010000110100_110_1_010000110100;
      patterns[41383] = 29'b1_010000110100_111_1_010000110100;
      patterns[41384] = 29'b1_010000110101_000_1_010000110101;
      patterns[41385] = 29'b1_010000110101_001_1_110101010000;
      patterns[41386] = 29'b1_010000110101_010_0_100001101011;
      patterns[41387] = 29'b1_010000110101_011_1_000011010110;
      patterns[41388] = 29'b1_010000110101_100_1_101000011010;
      patterns[41389] = 29'b1_010000110101_101_0_110100001101;
      patterns[41390] = 29'b1_010000110101_110_1_010000110101;
      patterns[41391] = 29'b1_010000110101_111_1_010000110101;
      patterns[41392] = 29'b1_010000110110_000_1_010000110110;
      patterns[41393] = 29'b1_010000110110_001_1_110110010000;
      patterns[41394] = 29'b1_010000110110_010_0_100001101101;
      patterns[41395] = 29'b1_010000110110_011_1_000011011010;
      patterns[41396] = 29'b1_010000110110_100_0_101000011011;
      patterns[41397] = 29'b1_010000110110_101_1_010100001101;
      patterns[41398] = 29'b1_010000110110_110_1_010000110110;
      patterns[41399] = 29'b1_010000110110_111_1_010000110110;
      patterns[41400] = 29'b1_010000110111_000_1_010000110111;
      patterns[41401] = 29'b1_010000110111_001_1_110111010000;
      patterns[41402] = 29'b1_010000110111_010_0_100001101111;
      patterns[41403] = 29'b1_010000110111_011_1_000011011110;
      patterns[41404] = 29'b1_010000110111_100_1_101000011011;
      patterns[41405] = 29'b1_010000110111_101_1_110100001101;
      patterns[41406] = 29'b1_010000110111_110_1_010000110111;
      patterns[41407] = 29'b1_010000110111_111_1_010000110111;
      patterns[41408] = 29'b1_010000111000_000_1_010000111000;
      patterns[41409] = 29'b1_010000111000_001_1_111000010000;
      patterns[41410] = 29'b1_010000111000_010_0_100001110001;
      patterns[41411] = 29'b1_010000111000_011_1_000011100010;
      patterns[41412] = 29'b1_010000111000_100_0_101000011100;
      patterns[41413] = 29'b1_010000111000_101_0_010100001110;
      patterns[41414] = 29'b1_010000111000_110_1_010000111000;
      patterns[41415] = 29'b1_010000111000_111_1_010000111000;
      patterns[41416] = 29'b1_010000111001_000_1_010000111001;
      patterns[41417] = 29'b1_010000111001_001_1_111001010000;
      patterns[41418] = 29'b1_010000111001_010_0_100001110011;
      patterns[41419] = 29'b1_010000111001_011_1_000011100110;
      patterns[41420] = 29'b1_010000111001_100_1_101000011100;
      patterns[41421] = 29'b1_010000111001_101_0_110100001110;
      patterns[41422] = 29'b1_010000111001_110_1_010000111001;
      patterns[41423] = 29'b1_010000111001_111_1_010000111001;
      patterns[41424] = 29'b1_010000111010_000_1_010000111010;
      patterns[41425] = 29'b1_010000111010_001_1_111010010000;
      patterns[41426] = 29'b1_010000111010_010_0_100001110101;
      patterns[41427] = 29'b1_010000111010_011_1_000011101010;
      patterns[41428] = 29'b1_010000111010_100_0_101000011101;
      patterns[41429] = 29'b1_010000111010_101_1_010100001110;
      patterns[41430] = 29'b1_010000111010_110_1_010000111010;
      patterns[41431] = 29'b1_010000111010_111_1_010000111010;
      patterns[41432] = 29'b1_010000111011_000_1_010000111011;
      patterns[41433] = 29'b1_010000111011_001_1_111011010000;
      patterns[41434] = 29'b1_010000111011_010_0_100001110111;
      patterns[41435] = 29'b1_010000111011_011_1_000011101110;
      patterns[41436] = 29'b1_010000111011_100_1_101000011101;
      patterns[41437] = 29'b1_010000111011_101_1_110100001110;
      patterns[41438] = 29'b1_010000111011_110_1_010000111011;
      patterns[41439] = 29'b1_010000111011_111_1_010000111011;
      patterns[41440] = 29'b1_010000111100_000_1_010000111100;
      patterns[41441] = 29'b1_010000111100_001_1_111100010000;
      patterns[41442] = 29'b1_010000111100_010_0_100001111001;
      patterns[41443] = 29'b1_010000111100_011_1_000011110010;
      patterns[41444] = 29'b1_010000111100_100_0_101000011110;
      patterns[41445] = 29'b1_010000111100_101_0_010100001111;
      patterns[41446] = 29'b1_010000111100_110_1_010000111100;
      patterns[41447] = 29'b1_010000111100_111_1_010000111100;
      patterns[41448] = 29'b1_010000111101_000_1_010000111101;
      patterns[41449] = 29'b1_010000111101_001_1_111101010000;
      patterns[41450] = 29'b1_010000111101_010_0_100001111011;
      patterns[41451] = 29'b1_010000111101_011_1_000011110110;
      patterns[41452] = 29'b1_010000111101_100_1_101000011110;
      patterns[41453] = 29'b1_010000111101_101_0_110100001111;
      patterns[41454] = 29'b1_010000111101_110_1_010000111101;
      patterns[41455] = 29'b1_010000111101_111_1_010000111101;
      patterns[41456] = 29'b1_010000111110_000_1_010000111110;
      patterns[41457] = 29'b1_010000111110_001_1_111110010000;
      patterns[41458] = 29'b1_010000111110_010_0_100001111101;
      patterns[41459] = 29'b1_010000111110_011_1_000011111010;
      patterns[41460] = 29'b1_010000111110_100_0_101000011111;
      patterns[41461] = 29'b1_010000111110_101_1_010100001111;
      patterns[41462] = 29'b1_010000111110_110_1_010000111110;
      patterns[41463] = 29'b1_010000111110_111_1_010000111110;
      patterns[41464] = 29'b1_010000111111_000_1_010000111111;
      patterns[41465] = 29'b1_010000111111_001_1_111111010000;
      patterns[41466] = 29'b1_010000111111_010_0_100001111111;
      patterns[41467] = 29'b1_010000111111_011_1_000011111110;
      patterns[41468] = 29'b1_010000111111_100_1_101000011111;
      patterns[41469] = 29'b1_010000111111_101_1_110100001111;
      patterns[41470] = 29'b1_010000111111_110_1_010000111111;
      patterns[41471] = 29'b1_010000111111_111_1_010000111111;
      patterns[41472] = 29'b1_010001000000_000_1_010001000000;
      patterns[41473] = 29'b1_010001000000_001_1_000000010001;
      patterns[41474] = 29'b1_010001000000_010_0_100010000001;
      patterns[41475] = 29'b1_010001000000_011_1_000100000010;
      patterns[41476] = 29'b1_010001000000_100_0_101000100000;
      patterns[41477] = 29'b1_010001000000_101_0_010100010000;
      patterns[41478] = 29'b1_010001000000_110_1_010001000000;
      patterns[41479] = 29'b1_010001000000_111_1_010001000000;
      patterns[41480] = 29'b1_010001000001_000_1_010001000001;
      patterns[41481] = 29'b1_010001000001_001_1_000001010001;
      patterns[41482] = 29'b1_010001000001_010_0_100010000011;
      patterns[41483] = 29'b1_010001000001_011_1_000100000110;
      patterns[41484] = 29'b1_010001000001_100_1_101000100000;
      patterns[41485] = 29'b1_010001000001_101_0_110100010000;
      patterns[41486] = 29'b1_010001000001_110_1_010001000001;
      patterns[41487] = 29'b1_010001000001_111_1_010001000001;
      patterns[41488] = 29'b1_010001000010_000_1_010001000010;
      patterns[41489] = 29'b1_010001000010_001_1_000010010001;
      patterns[41490] = 29'b1_010001000010_010_0_100010000101;
      patterns[41491] = 29'b1_010001000010_011_1_000100001010;
      patterns[41492] = 29'b1_010001000010_100_0_101000100001;
      patterns[41493] = 29'b1_010001000010_101_1_010100010000;
      patterns[41494] = 29'b1_010001000010_110_1_010001000010;
      patterns[41495] = 29'b1_010001000010_111_1_010001000010;
      patterns[41496] = 29'b1_010001000011_000_1_010001000011;
      patterns[41497] = 29'b1_010001000011_001_1_000011010001;
      patterns[41498] = 29'b1_010001000011_010_0_100010000111;
      patterns[41499] = 29'b1_010001000011_011_1_000100001110;
      patterns[41500] = 29'b1_010001000011_100_1_101000100001;
      patterns[41501] = 29'b1_010001000011_101_1_110100010000;
      patterns[41502] = 29'b1_010001000011_110_1_010001000011;
      patterns[41503] = 29'b1_010001000011_111_1_010001000011;
      patterns[41504] = 29'b1_010001000100_000_1_010001000100;
      patterns[41505] = 29'b1_010001000100_001_1_000100010001;
      patterns[41506] = 29'b1_010001000100_010_0_100010001001;
      patterns[41507] = 29'b1_010001000100_011_1_000100010010;
      patterns[41508] = 29'b1_010001000100_100_0_101000100010;
      patterns[41509] = 29'b1_010001000100_101_0_010100010001;
      patterns[41510] = 29'b1_010001000100_110_1_010001000100;
      patterns[41511] = 29'b1_010001000100_111_1_010001000100;
      patterns[41512] = 29'b1_010001000101_000_1_010001000101;
      patterns[41513] = 29'b1_010001000101_001_1_000101010001;
      patterns[41514] = 29'b1_010001000101_010_0_100010001011;
      patterns[41515] = 29'b1_010001000101_011_1_000100010110;
      patterns[41516] = 29'b1_010001000101_100_1_101000100010;
      patterns[41517] = 29'b1_010001000101_101_0_110100010001;
      patterns[41518] = 29'b1_010001000101_110_1_010001000101;
      patterns[41519] = 29'b1_010001000101_111_1_010001000101;
      patterns[41520] = 29'b1_010001000110_000_1_010001000110;
      patterns[41521] = 29'b1_010001000110_001_1_000110010001;
      patterns[41522] = 29'b1_010001000110_010_0_100010001101;
      patterns[41523] = 29'b1_010001000110_011_1_000100011010;
      patterns[41524] = 29'b1_010001000110_100_0_101000100011;
      patterns[41525] = 29'b1_010001000110_101_1_010100010001;
      patterns[41526] = 29'b1_010001000110_110_1_010001000110;
      patterns[41527] = 29'b1_010001000110_111_1_010001000110;
      patterns[41528] = 29'b1_010001000111_000_1_010001000111;
      patterns[41529] = 29'b1_010001000111_001_1_000111010001;
      patterns[41530] = 29'b1_010001000111_010_0_100010001111;
      patterns[41531] = 29'b1_010001000111_011_1_000100011110;
      patterns[41532] = 29'b1_010001000111_100_1_101000100011;
      patterns[41533] = 29'b1_010001000111_101_1_110100010001;
      patterns[41534] = 29'b1_010001000111_110_1_010001000111;
      patterns[41535] = 29'b1_010001000111_111_1_010001000111;
      patterns[41536] = 29'b1_010001001000_000_1_010001001000;
      patterns[41537] = 29'b1_010001001000_001_1_001000010001;
      patterns[41538] = 29'b1_010001001000_010_0_100010010001;
      patterns[41539] = 29'b1_010001001000_011_1_000100100010;
      patterns[41540] = 29'b1_010001001000_100_0_101000100100;
      patterns[41541] = 29'b1_010001001000_101_0_010100010010;
      patterns[41542] = 29'b1_010001001000_110_1_010001001000;
      patterns[41543] = 29'b1_010001001000_111_1_010001001000;
      patterns[41544] = 29'b1_010001001001_000_1_010001001001;
      patterns[41545] = 29'b1_010001001001_001_1_001001010001;
      patterns[41546] = 29'b1_010001001001_010_0_100010010011;
      patterns[41547] = 29'b1_010001001001_011_1_000100100110;
      patterns[41548] = 29'b1_010001001001_100_1_101000100100;
      patterns[41549] = 29'b1_010001001001_101_0_110100010010;
      patterns[41550] = 29'b1_010001001001_110_1_010001001001;
      patterns[41551] = 29'b1_010001001001_111_1_010001001001;
      patterns[41552] = 29'b1_010001001010_000_1_010001001010;
      patterns[41553] = 29'b1_010001001010_001_1_001010010001;
      patterns[41554] = 29'b1_010001001010_010_0_100010010101;
      patterns[41555] = 29'b1_010001001010_011_1_000100101010;
      patterns[41556] = 29'b1_010001001010_100_0_101000100101;
      patterns[41557] = 29'b1_010001001010_101_1_010100010010;
      patterns[41558] = 29'b1_010001001010_110_1_010001001010;
      patterns[41559] = 29'b1_010001001010_111_1_010001001010;
      patterns[41560] = 29'b1_010001001011_000_1_010001001011;
      patterns[41561] = 29'b1_010001001011_001_1_001011010001;
      patterns[41562] = 29'b1_010001001011_010_0_100010010111;
      patterns[41563] = 29'b1_010001001011_011_1_000100101110;
      patterns[41564] = 29'b1_010001001011_100_1_101000100101;
      patterns[41565] = 29'b1_010001001011_101_1_110100010010;
      patterns[41566] = 29'b1_010001001011_110_1_010001001011;
      patterns[41567] = 29'b1_010001001011_111_1_010001001011;
      patterns[41568] = 29'b1_010001001100_000_1_010001001100;
      patterns[41569] = 29'b1_010001001100_001_1_001100010001;
      patterns[41570] = 29'b1_010001001100_010_0_100010011001;
      patterns[41571] = 29'b1_010001001100_011_1_000100110010;
      patterns[41572] = 29'b1_010001001100_100_0_101000100110;
      patterns[41573] = 29'b1_010001001100_101_0_010100010011;
      patterns[41574] = 29'b1_010001001100_110_1_010001001100;
      patterns[41575] = 29'b1_010001001100_111_1_010001001100;
      patterns[41576] = 29'b1_010001001101_000_1_010001001101;
      patterns[41577] = 29'b1_010001001101_001_1_001101010001;
      patterns[41578] = 29'b1_010001001101_010_0_100010011011;
      patterns[41579] = 29'b1_010001001101_011_1_000100110110;
      patterns[41580] = 29'b1_010001001101_100_1_101000100110;
      patterns[41581] = 29'b1_010001001101_101_0_110100010011;
      patterns[41582] = 29'b1_010001001101_110_1_010001001101;
      patterns[41583] = 29'b1_010001001101_111_1_010001001101;
      patterns[41584] = 29'b1_010001001110_000_1_010001001110;
      patterns[41585] = 29'b1_010001001110_001_1_001110010001;
      patterns[41586] = 29'b1_010001001110_010_0_100010011101;
      patterns[41587] = 29'b1_010001001110_011_1_000100111010;
      patterns[41588] = 29'b1_010001001110_100_0_101000100111;
      patterns[41589] = 29'b1_010001001110_101_1_010100010011;
      patterns[41590] = 29'b1_010001001110_110_1_010001001110;
      patterns[41591] = 29'b1_010001001110_111_1_010001001110;
      patterns[41592] = 29'b1_010001001111_000_1_010001001111;
      patterns[41593] = 29'b1_010001001111_001_1_001111010001;
      patterns[41594] = 29'b1_010001001111_010_0_100010011111;
      patterns[41595] = 29'b1_010001001111_011_1_000100111110;
      patterns[41596] = 29'b1_010001001111_100_1_101000100111;
      patterns[41597] = 29'b1_010001001111_101_1_110100010011;
      patterns[41598] = 29'b1_010001001111_110_1_010001001111;
      patterns[41599] = 29'b1_010001001111_111_1_010001001111;
      patterns[41600] = 29'b1_010001010000_000_1_010001010000;
      patterns[41601] = 29'b1_010001010000_001_1_010000010001;
      patterns[41602] = 29'b1_010001010000_010_0_100010100001;
      patterns[41603] = 29'b1_010001010000_011_1_000101000010;
      patterns[41604] = 29'b1_010001010000_100_0_101000101000;
      patterns[41605] = 29'b1_010001010000_101_0_010100010100;
      patterns[41606] = 29'b1_010001010000_110_1_010001010000;
      patterns[41607] = 29'b1_010001010000_111_1_010001010000;
      patterns[41608] = 29'b1_010001010001_000_1_010001010001;
      patterns[41609] = 29'b1_010001010001_001_1_010001010001;
      patterns[41610] = 29'b1_010001010001_010_0_100010100011;
      patterns[41611] = 29'b1_010001010001_011_1_000101000110;
      patterns[41612] = 29'b1_010001010001_100_1_101000101000;
      patterns[41613] = 29'b1_010001010001_101_0_110100010100;
      patterns[41614] = 29'b1_010001010001_110_1_010001010001;
      patterns[41615] = 29'b1_010001010001_111_1_010001010001;
      patterns[41616] = 29'b1_010001010010_000_1_010001010010;
      patterns[41617] = 29'b1_010001010010_001_1_010010010001;
      patterns[41618] = 29'b1_010001010010_010_0_100010100101;
      patterns[41619] = 29'b1_010001010010_011_1_000101001010;
      patterns[41620] = 29'b1_010001010010_100_0_101000101001;
      patterns[41621] = 29'b1_010001010010_101_1_010100010100;
      patterns[41622] = 29'b1_010001010010_110_1_010001010010;
      patterns[41623] = 29'b1_010001010010_111_1_010001010010;
      patterns[41624] = 29'b1_010001010011_000_1_010001010011;
      patterns[41625] = 29'b1_010001010011_001_1_010011010001;
      patterns[41626] = 29'b1_010001010011_010_0_100010100111;
      patterns[41627] = 29'b1_010001010011_011_1_000101001110;
      patterns[41628] = 29'b1_010001010011_100_1_101000101001;
      patterns[41629] = 29'b1_010001010011_101_1_110100010100;
      patterns[41630] = 29'b1_010001010011_110_1_010001010011;
      patterns[41631] = 29'b1_010001010011_111_1_010001010011;
      patterns[41632] = 29'b1_010001010100_000_1_010001010100;
      patterns[41633] = 29'b1_010001010100_001_1_010100010001;
      patterns[41634] = 29'b1_010001010100_010_0_100010101001;
      patterns[41635] = 29'b1_010001010100_011_1_000101010010;
      patterns[41636] = 29'b1_010001010100_100_0_101000101010;
      patterns[41637] = 29'b1_010001010100_101_0_010100010101;
      patterns[41638] = 29'b1_010001010100_110_1_010001010100;
      patterns[41639] = 29'b1_010001010100_111_1_010001010100;
      patterns[41640] = 29'b1_010001010101_000_1_010001010101;
      patterns[41641] = 29'b1_010001010101_001_1_010101010001;
      patterns[41642] = 29'b1_010001010101_010_0_100010101011;
      patterns[41643] = 29'b1_010001010101_011_1_000101010110;
      patterns[41644] = 29'b1_010001010101_100_1_101000101010;
      patterns[41645] = 29'b1_010001010101_101_0_110100010101;
      patterns[41646] = 29'b1_010001010101_110_1_010001010101;
      patterns[41647] = 29'b1_010001010101_111_1_010001010101;
      patterns[41648] = 29'b1_010001010110_000_1_010001010110;
      patterns[41649] = 29'b1_010001010110_001_1_010110010001;
      patterns[41650] = 29'b1_010001010110_010_0_100010101101;
      patterns[41651] = 29'b1_010001010110_011_1_000101011010;
      patterns[41652] = 29'b1_010001010110_100_0_101000101011;
      patterns[41653] = 29'b1_010001010110_101_1_010100010101;
      patterns[41654] = 29'b1_010001010110_110_1_010001010110;
      patterns[41655] = 29'b1_010001010110_111_1_010001010110;
      patterns[41656] = 29'b1_010001010111_000_1_010001010111;
      patterns[41657] = 29'b1_010001010111_001_1_010111010001;
      patterns[41658] = 29'b1_010001010111_010_0_100010101111;
      patterns[41659] = 29'b1_010001010111_011_1_000101011110;
      patterns[41660] = 29'b1_010001010111_100_1_101000101011;
      patterns[41661] = 29'b1_010001010111_101_1_110100010101;
      patterns[41662] = 29'b1_010001010111_110_1_010001010111;
      patterns[41663] = 29'b1_010001010111_111_1_010001010111;
      patterns[41664] = 29'b1_010001011000_000_1_010001011000;
      patterns[41665] = 29'b1_010001011000_001_1_011000010001;
      patterns[41666] = 29'b1_010001011000_010_0_100010110001;
      patterns[41667] = 29'b1_010001011000_011_1_000101100010;
      patterns[41668] = 29'b1_010001011000_100_0_101000101100;
      patterns[41669] = 29'b1_010001011000_101_0_010100010110;
      patterns[41670] = 29'b1_010001011000_110_1_010001011000;
      patterns[41671] = 29'b1_010001011000_111_1_010001011000;
      patterns[41672] = 29'b1_010001011001_000_1_010001011001;
      patterns[41673] = 29'b1_010001011001_001_1_011001010001;
      patterns[41674] = 29'b1_010001011001_010_0_100010110011;
      patterns[41675] = 29'b1_010001011001_011_1_000101100110;
      patterns[41676] = 29'b1_010001011001_100_1_101000101100;
      patterns[41677] = 29'b1_010001011001_101_0_110100010110;
      patterns[41678] = 29'b1_010001011001_110_1_010001011001;
      patterns[41679] = 29'b1_010001011001_111_1_010001011001;
      patterns[41680] = 29'b1_010001011010_000_1_010001011010;
      patterns[41681] = 29'b1_010001011010_001_1_011010010001;
      patterns[41682] = 29'b1_010001011010_010_0_100010110101;
      patterns[41683] = 29'b1_010001011010_011_1_000101101010;
      patterns[41684] = 29'b1_010001011010_100_0_101000101101;
      patterns[41685] = 29'b1_010001011010_101_1_010100010110;
      patterns[41686] = 29'b1_010001011010_110_1_010001011010;
      patterns[41687] = 29'b1_010001011010_111_1_010001011010;
      patterns[41688] = 29'b1_010001011011_000_1_010001011011;
      patterns[41689] = 29'b1_010001011011_001_1_011011010001;
      patterns[41690] = 29'b1_010001011011_010_0_100010110111;
      patterns[41691] = 29'b1_010001011011_011_1_000101101110;
      patterns[41692] = 29'b1_010001011011_100_1_101000101101;
      patterns[41693] = 29'b1_010001011011_101_1_110100010110;
      patterns[41694] = 29'b1_010001011011_110_1_010001011011;
      patterns[41695] = 29'b1_010001011011_111_1_010001011011;
      patterns[41696] = 29'b1_010001011100_000_1_010001011100;
      patterns[41697] = 29'b1_010001011100_001_1_011100010001;
      patterns[41698] = 29'b1_010001011100_010_0_100010111001;
      patterns[41699] = 29'b1_010001011100_011_1_000101110010;
      patterns[41700] = 29'b1_010001011100_100_0_101000101110;
      patterns[41701] = 29'b1_010001011100_101_0_010100010111;
      patterns[41702] = 29'b1_010001011100_110_1_010001011100;
      patterns[41703] = 29'b1_010001011100_111_1_010001011100;
      patterns[41704] = 29'b1_010001011101_000_1_010001011101;
      patterns[41705] = 29'b1_010001011101_001_1_011101010001;
      patterns[41706] = 29'b1_010001011101_010_0_100010111011;
      patterns[41707] = 29'b1_010001011101_011_1_000101110110;
      patterns[41708] = 29'b1_010001011101_100_1_101000101110;
      patterns[41709] = 29'b1_010001011101_101_0_110100010111;
      patterns[41710] = 29'b1_010001011101_110_1_010001011101;
      patterns[41711] = 29'b1_010001011101_111_1_010001011101;
      patterns[41712] = 29'b1_010001011110_000_1_010001011110;
      patterns[41713] = 29'b1_010001011110_001_1_011110010001;
      patterns[41714] = 29'b1_010001011110_010_0_100010111101;
      patterns[41715] = 29'b1_010001011110_011_1_000101111010;
      patterns[41716] = 29'b1_010001011110_100_0_101000101111;
      patterns[41717] = 29'b1_010001011110_101_1_010100010111;
      patterns[41718] = 29'b1_010001011110_110_1_010001011110;
      patterns[41719] = 29'b1_010001011110_111_1_010001011110;
      patterns[41720] = 29'b1_010001011111_000_1_010001011111;
      patterns[41721] = 29'b1_010001011111_001_1_011111010001;
      patterns[41722] = 29'b1_010001011111_010_0_100010111111;
      patterns[41723] = 29'b1_010001011111_011_1_000101111110;
      patterns[41724] = 29'b1_010001011111_100_1_101000101111;
      patterns[41725] = 29'b1_010001011111_101_1_110100010111;
      patterns[41726] = 29'b1_010001011111_110_1_010001011111;
      patterns[41727] = 29'b1_010001011111_111_1_010001011111;
      patterns[41728] = 29'b1_010001100000_000_1_010001100000;
      patterns[41729] = 29'b1_010001100000_001_1_100000010001;
      patterns[41730] = 29'b1_010001100000_010_0_100011000001;
      patterns[41731] = 29'b1_010001100000_011_1_000110000010;
      patterns[41732] = 29'b1_010001100000_100_0_101000110000;
      patterns[41733] = 29'b1_010001100000_101_0_010100011000;
      patterns[41734] = 29'b1_010001100000_110_1_010001100000;
      patterns[41735] = 29'b1_010001100000_111_1_010001100000;
      patterns[41736] = 29'b1_010001100001_000_1_010001100001;
      patterns[41737] = 29'b1_010001100001_001_1_100001010001;
      patterns[41738] = 29'b1_010001100001_010_0_100011000011;
      patterns[41739] = 29'b1_010001100001_011_1_000110000110;
      patterns[41740] = 29'b1_010001100001_100_1_101000110000;
      patterns[41741] = 29'b1_010001100001_101_0_110100011000;
      patterns[41742] = 29'b1_010001100001_110_1_010001100001;
      patterns[41743] = 29'b1_010001100001_111_1_010001100001;
      patterns[41744] = 29'b1_010001100010_000_1_010001100010;
      patterns[41745] = 29'b1_010001100010_001_1_100010010001;
      patterns[41746] = 29'b1_010001100010_010_0_100011000101;
      patterns[41747] = 29'b1_010001100010_011_1_000110001010;
      patterns[41748] = 29'b1_010001100010_100_0_101000110001;
      patterns[41749] = 29'b1_010001100010_101_1_010100011000;
      patterns[41750] = 29'b1_010001100010_110_1_010001100010;
      patterns[41751] = 29'b1_010001100010_111_1_010001100010;
      patterns[41752] = 29'b1_010001100011_000_1_010001100011;
      patterns[41753] = 29'b1_010001100011_001_1_100011010001;
      patterns[41754] = 29'b1_010001100011_010_0_100011000111;
      patterns[41755] = 29'b1_010001100011_011_1_000110001110;
      patterns[41756] = 29'b1_010001100011_100_1_101000110001;
      patterns[41757] = 29'b1_010001100011_101_1_110100011000;
      patterns[41758] = 29'b1_010001100011_110_1_010001100011;
      patterns[41759] = 29'b1_010001100011_111_1_010001100011;
      patterns[41760] = 29'b1_010001100100_000_1_010001100100;
      patterns[41761] = 29'b1_010001100100_001_1_100100010001;
      patterns[41762] = 29'b1_010001100100_010_0_100011001001;
      patterns[41763] = 29'b1_010001100100_011_1_000110010010;
      patterns[41764] = 29'b1_010001100100_100_0_101000110010;
      patterns[41765] = 29'b1_010001100100_101_0_010100011001;
      patterns[41766] = 29'b1_010001100100_110_1_010001100100;
      patterns[41767] = 29'b1_010001100100_111_1_010001100100;
      patterns[41768] = 29'b1_010001100101_000_1_010001100101;
      patterns[41769] = 29'b1_010001100101_001_1_100101010001;
      patterns[41770] = 29'b1_010001100101_010_0_100011001011;
      patterns[41771] = 29'b1_010001100101_011_1_000110010110;
      patterns[41772] = 29'b1_010001100101_100_1_101000110010;
      patterns[41773] = 29'b1_010001100101_101_0_110100011001;
      patterns[41774] = 29'b1_010001100101_110_1_010001100101;
      patterns[41775] = 29'b1_010001100101_111_1_010001100101;
      patterns[41776] = 29'b1_010001100110_000_1_010001100110;
      patterns[41777] = 29'b1_010001100110_001_1_100110010001;
      patterns[41778] = 29'b1_010001100110_010_0_100011001101;
      patterns[41779] = 29'b1_010001100110_011_1_000110011010;
      patterns[41780] = 29'b1_010001100110_100_0_101000110011;
      patterns[41781] = 29'b1_010001100110_101_1_010100011001;
      patterns[41782] = 29'b1_010001100110_110_1_010001100110;
      patterns[41783] = 29'b1_010001100110_111_1_010001100110;
      patterns[41784] = 29'b1_010001100111_000_1_010001100111;
      patterns[41785] = 29'b1_010001100111_001_1_100111010001;
      patterns[41786] = 29'b1_010001100111_010_0_100011001111;
      patterns[41787] = 29'b1_010001100111_011_1_000110011110;
      patterns[41788] = 29'b1_010001100111_100_1_101000110011;
      patterns[41789] = 29'b1_010001100111_101_1_110100011001;
      patterns[41790] = 29'b1_010001100111_110_1_010001100111;
      patterns[41791] = 29'b1_010001100111_111_1_010001100111;
      patterns[41792] = 29'b1_010001101000_000_1_010001101000;
      patterns[41793] = 29'b1_010001101000_001_1_101000010001;
      patterns[41794] = 29'b1_010001101000_010_0_100011010001;
      patterns[41795] = 29'b1_010001101000_011_1_000110100010;
      patterns[41796] = 29'b1_010001101000_100_0_101000110100;
      patterns[41797] = 29'b1_010001101000_101_0_010100011010;
      patterns[41798] = 29'b1_010001101000_110_1_010001101000;
      patterns[41799] = 29'b1_010001101000_111_1_010001101000;
      patterns[41800] = 29'b1_010001101001_000_1_010001101001;
      patterns[41801] = 29'b1_010001101001_001_1_101001010001;
      patterns[41802] = 29'b1_010001101001_010_0_100011010011;
      patterns[41803] = 29'b1_010001101001_011_1_000110100110;
      patterns[41804] = 29'b1_010001101001_100_1_101000110100;
      patterns[41805] = 29'b1_010001101001_101_0_110100011010;
      patterns[41806] = 29'b1_010001101001_110_1_010001101001;
      patterns[41807] = 29'b1_010001101001_111_1_010001101001;
      patterns[41808] = 29'b1_010001101010_000_1_010001101010;
      patterns[41809] = 29'b1_010001101010_001_1_101010010001;
      patterns[41810] = 29'b1_010001101010_010_0_100011010101;
      patterns[41811] = 29'b1_010001101010_011_1_000110101010;
      patterns[41812] = 29'b1_010001101010_100_0_101000110101;
      patterns[41813] = 29'b1_010001101010_101_1_010100011010;
      patterns[41814] = 29'b1_010001101010_110_1_010001101010;
      patterns[41815] = 29'b1_010001101010_111_1_010001101010;
      patterns[41816] = 29'b1_010001101011_000_1_010001101011;
      patterns[41817] = 29'b1_010001101011_001_1_101011010001;
      patterns[41818] = 29'b1_010001101011_010_0_100011010111;
      patterns[41819] = 29'b1_010001101011_011_1_000110101110;
      patterns[41820] = 29'b1_010001101011_100_1_101000110101;
      patterns[41821] = 29'b1_010001101011_101_1_110100011010;
      patterns[41822] = 29'b1_010001101011_110_1_010001101011;
      patterns[41823] = 29'b1_010001101011_111_1_010001101011;
      patterns[41824] = 29'b1_010001101100_000_1_010001101100;
      patterns[41825] = 29'b1_010001101100_001_1_101100010001;
      patterns[41826] = 29'b1_010001101100_010_0_100011011001;
      patterns[41827] = 29'b1_010001101100_011_1_000110110010;
      patterns[41828] = 29'b1_010001101100_100_0_101000110110;
      patterns[41829] = 29'b1_010001101100_101_0_010100011011;
      patterns[41830] = 29'b1_010001101100_110_1_010001101100;
      patterns[41831] = 29'b1_010001101100_111_1_010001101100;
      patterns[41832] = 29'b1_010001101101_000_1_010001101101;
      patterns[41833] = 29'b1_010001101101_001_1_101101010001;
      patterns[41834] = 29'b1_010001101101_010_0_100011011011;
      patterns[41835] = 29'b1_010001101101_011_1_000110110110;
      patterns[41836] = 29'b1_010001101101_100_1_101000110110;
      patterns[41837] = 29'b1_010001101101_101_0_110100011011;
      patterns[41838] = 29'b1_010001101101_110_1_010001101101;
      patterns[41839] = 29'b1_010001101101_111_1_010001101101;
      patterns[41840] = 29'b1_010001101110_000_1_010001101110;
      patterns[41841] = 29'b1_010001101110_001_1_101110010001;
      patterns[41842] = 29'b1_010001101110_010_0_100011011101;
      patterns[41843] = 29'b1_010001101110_011_1_000110111010;
      patterns[41844] = 29'b1_010001101110_100_0_101000110111;
      patterns[41845] = 29'b1_010001101110_101_1_010100011011;
      patterns[41846] = 29'b1_010001101110_110_1_010001101110;
      patterns[41847] = 29'b1_010001101110_111_1_010001101110;
      patterns[41848] = 29'b1_010001101111_000_1_010001101111;
      patterns[41849] = 29'b1_010001101111_001_1_101111010001;
      patterns[41850] = 29'b1_010001101111_010_0_100011011111;
      patterns[41851] = 29'b1_010001101111_011_1_000110111110;
      patterns[41852] = 29'b1_010001101111_100_1_101000110111;
      patterns[41853] = 29'b1_010001101111_101_1_110100011011;
      patterns[41854] = 29'b1_010001101111_110_1_010001101111;
      patterns[41855] = 29'b1_010001101111_111_1_010001101111;
      patterns[41856] = 29'b1_010001110000_000_1_010001110000;
      patterns[41857] = 29'b1_010001110000_001_1_110000010001;
      patterns[41858] = 29'b1_010001110000_010_0_100011100001;
      patterns[41859] = 29'b1_010001110000_011_1_000111000010;
      patterns[41860] = 29'b1_010001110000_100_0_101000111000;
      patterns[41861] = 29'b1_010001110000_101_0_010100011100;
      patterns[41862] = 29'b1_010001110000_110_1_010001110000;
      patterns[41863] = 29'b1_010001110000_111_1_010001110000;
      patterns[41864] = 29'b1_010001110001_000_1_010001110001;
      patterns[41865] = 29'b1_010001110001_001_1_110001010001;
      patterns[41866] = 29'b1_010001110001_010_0_100011100011;
      patterns[41867] = 29'b1_010001110001_011_1_000111000110;
      patterns[41868] = 29'b1_010001110001_100_1_101000111000;
      patterns[41869] = 29'b1_010001110001_101_0_110100011100;
      patterns[41870] = 29'b1_010001110001_110_1_010001110001;
      patterns[41871] = 29'b1_010001110001_111_1_010001110001;
      patterns[41872] = 29'b1_010001110010_000_1_010001110010;
      patterns[41873] = 29'b1_010001110010_001_1_110010010001;
      patterns[41874] = 29'b1_010001110010_010_0_100011100101;
      patterns[41875] = 29'b1_010001110010_011_1_000111001010;
      patterns[41876] = 29'b1_010001110010_100_0_101000111001;
      patterns[41877] = 29'b1_010001110010_101_1_010100011100;
      patterns[41878] = 29'b1_010001110010_110_1_010001110010;
      patterns[41879] = 29'b1_010001110010_111_1_010001110010;
      patterns[41880] = 29'b1_010001110011_000_1_010001110011;
      patterns[41881] = 29'b1_010001110011_001_1_110011010001;
      patterns[41882] = 29'b1_010001110011_010_0_100011100111;
      patterns[41883] = 29'b1_010001110011_011_1_000111001110;
      patterns[41884] = 29'b1_010001110011_100_1_101000111001;
      patterns[41885] = 29'b1_010001110011_101_1_110100011100;
      patterns[41886] = 29'b1_010001110011_110_1_010001110011;
      patterns[41887] = 29'b1_010001110011_111_1_010001110011;
      patterns[41888] = 29'b1_010001110100_000_1_010001110100;
      patterns[41889] = 29'b1_010001110100_001_1_110100010001;
      patterns[41890] = 29'b1_010001110100_010_0_100011101001;
      patterns[41891] = 29'b1_010001110100_011_1_000111010010;
      patterns[41892] = 29'b1_010001110100_100_0_101000111010;
      patterns[41893] = 29'b1_010001110100_101_0_010100011101;
      patterns[41894] = 29'b1_010001110100_110_1_010001110100;
      patterns[41895] = 29'b1_010001110100_111_1_010001110100;
      patterns[41896] = 29'b1_010001110101_000_1_010001110101;
      patterns[41897] = 29'b1_010001110101_001_1_110101010001;
      patterns[41898] = 29'b1_010001110101_010_0_100011101011;
      patterns[41899] = 29'b1_010001110101_011_1_000111010110;
      patterns[41900] = 29'b1_010001110101_100_1_101000111010;
      patterns[41901] = 29'b1_010001110101_101_0_110100011101;
      patterns[41902] = 29'b1_010001110101_110_1_010001110101;
      patterns[41903] = 29'b1_010001110101_111_1_010001110101;
      patterns[41904] = 29'b1_010001110110_000_1_010001110110;
      patterns[41905] = 29'b1_010001110110_001_1_110110010001;
      patterns[41906] = 29'b1_010001110110_010_0_100011101101;
      patterns[41907] = 29'b1_010001110110_011_1_000111011010;
      patterns[41908] = 29'b1_010001110110_100_0_101000111011;
      patterns[41909] = 29'b1_010001110110_101_1_010100011101;
      patterns[41910] = 29'b1_010001110110_110_1_010001110110;
      patterns[41911] = 29'b1_010001110110_111_1_010001110110;
      patterns[41912] = 29'b1_010001110111_000_1_010001110111;
      patterns[41913] = 29'b1_010001110111_001_1_110111010001;
      patterns[41914] = 29'b1_010001110111_010_0_100011101111;
      patterns[41915] = 29'b1_010001110111_011_1_000111011110;
      patterns[41916] = 29'b1_010001110111_100_1_101000111011;
      patterns[41917] = 29'b1_010001110111_101_1_110100011101;
      patterns[41918] = 29'b1_010001110111_110_1_010001110111;
      patterns[41919] = 29'b1_010001110111_111_1_010001110111;
      patterns[41920] = 29'b1_010001111000_000_1_010001111000;
      patterns[41921] = 29'b1_010001111000_001_1_111000010001;
      patterns[41922] = 29'b1_010001111000_010_0_100011110001;
      patterns[41923] = 29'b1_010001111000_011_1_000111100010;
      patterns[41924] = 29'b1_010001111000_100_0_101000111100;
      patterns[41925] = 29'b1_010001111000_101_0_010100011110;
      patterns[41926] = 29'b1_010001111000_110_1_010001111000;
      patterns[41927] = 29'b1_010001111000_111_1_010001111000;
      patterns[41928] = 29'b1_010001111001_000_1_010001111001;
      patterns[41929] = 29'b1_010001111001_001_1_111001010001;
      patterns[41930] = 29'b1_010001111001_010_0_100011110011;
      patterns[41931] = 29'b1_010001111001_011_1_000111100110;
      patterns[41932] = 29'b1_010001111001_100_1_101000111100;
      patterns[41933] = 29'b1_010001111001_101_0_110100011110;
      patterns[41934] = 29'b1_010001111001_110_1_010001111001;
      patterns[41935] = 29'b1_010001111001_111_1_010001111001;
      patterns[41936] = 29'b1_010001111010_000_1_010001111010;
      patterns[41937] = 29'b1_010001111010_001_1_111010010001;
      patterns[41938] = 29'b1_010001111010_010_0_100011110101;
      patterns[41939] = 29'b1_010001111010_011_1_000111101010;
      patterns[41940] = 29'b1_010001111010_100_0_101000111101;
      patterns[41941] = 29'b1_010001111010_101_1_010100011110;
      patterns[41942] = 29'b1_010001111010_110_1_010001111010;
      patterns[41943] = 29'b1_010001111010_111_1_010001111010;
      patterns[41944] = 29'b1_010001111011_000_1_010001111011;
      patterns[41945] = 29'b1_010001111011_001_1_111011010001;
      patterns[41946] = 29'b1_010001111011_010_0_100011110111;
      patterns[41947] = 29'b1_010001111011_011_1_000111101110;
      patterns[41948] = 29'b1_010001111011_100_1_101000111101;
      patterns[41949] = 29'b1_010001111011_101_1_110100011110;
      patterns[41950] = 29'b1_010001111011_110_1_010001111011;
      patterns[41951] = 29'b1_010001111011_111_1_010001111011;
      patterns[41952] = 29'b1_010001111100_000_1_010001111100;
      patterns[41953] = 29'b1_010001111100_001_1_111100010001;
      patterns[41954] = 29'b1_010001111100_010_0_100011111001;
      patterns[41955] = 29'b1_010001111100_011_1_000111110010;
      patterns[41956] = 29'b1_010001111100_100_0_101000111110;
      patterns[41957] = 29'b1_010001111100_101_0_010100011111;
      patterns[41958] = 29'b1_010001111100_110_1_010001111100;
      patterns[41959] = 29'b1_010001111100_111_1_010001111100;
      patterns[41960] = 29'b1_010001111101_000_1_010001111101;
      patterns[41961] = 29'b1_010001111101_001_1_111101010001;
      patterns[41962] = 29'b1_010001111101_010_0_100011111011;
      patterns[41963] = 29'b1_010001111101_011_1_000111110110;
      patterns[41964] = 29'b1_010001111101_100_1_101000111110;
      patterns[41965] = 29'b1_010001111101_101_0_110100011111;
      patterns[41966] = 29'b1_010001111101_110_1_010001111101;
      patterns[41967] = 29'b1_010001111101_111_1_010001111101;
      patterns[41968] = 29'b1_010001111110_000_1_010001111110;
      patterns[41969] = 29'b1_010001111110_001_1_111110010001;
      patterns[41970] = 29'b1_010001111110_010_0_100011111101;
      patterns[41971] = 29'b1_010001111110_011_1_000111111010;
      patterns[41972] = 29'b1_010001111110_100_0_101000111111;
      patterns[41973] = 29'b1_010001111110_101_1_010100011111;
      patterns[41974] = 29'b1_010001111110_110_1_010001111110;
      patterns[41975] = 29'b1_010001111110_111_1_010001111110;
      patterns[41976] = 29'b1_010001111111_000_1_010001111111;
      patterns[41977] = 29'b1_010001111111_001_1_111111010001;
      patterns[41978] = 29'b1_010001111111_010_0_100011111111;
      patterns[41979] = 29'b1_010001111111_011_1_000111111110;
      patterns[41980] = 29'b1_010001111111_100_1_101000111111;
      patterns[41981] = 29'b1_010001111111_101_1_110100011111;
      patterns[41982] = 29'b1_010001111111_110_1_010001111111;
      patterns[41983] = 29'b1_010001111111_111_1_010001111111;
      patterns[41984] = 29'b1_010010000000_000_1_010010000000;
      patterns[41985] = 29'b1_010010000000_001_1_000000010010;
      patterns[41986] = 29'b1_010010000000_010_0_100100000001;
      patterns[41987] = 29'b1_010010000000_011_1_001000000010;
      patterns[41988] = 29'b1_010010000000_100_0_101001000000;
      patterns[41989] = 29'b1_010010000000_101_0_010100100000;
      patterns[41990] = 29'b1_010010000000_110_1_010010000000;
      patterns[41991] = 29'b1_010010000000_111_1_010010000000;
      patterns[41992] = 29'b1_010010000001_000_1_010010000001;
      patterns[41993] = 29'b1_010010000001_001_1_000001010010;
      patterns[41994] = 29'b1_010010000001_010_0_100100000011;
      patterns[41995] = 29'b1_010010000001_011_1_001000000110;
      patterns[41996] = 29'b1_010010000001_100_1_101001000000;
      patterns[41997] = 29'b1_010010000001_101_0_110100100000;
      patterns[41998] = 29'b1_010010000001_110_1_010010000001;
      patterns[41999] = 29'b1_010010000001_111_1_010010000001;
      patterns[42000] = 29'b1_010010000010_000_1_010010000010;
      patterns[42001] = 29'b1_010010000010_001_1_000010010010;
      patterns[42002] = 29'b1_010010000010_010_0_100100000101;
      patterns[42003] = 29'b1_010010000010_011_1_001000001010;
      patterns[42004] = 29'b1_010010000010_100_0_101001000001;
      patterns[42005] = 29'b1_010010000010_101_1_010100100000;
      patterns[42006] = 29'b1_010010000010_110_1_010010000010;
      patterns[42007] = 29'b1_010010000010_111_1_010010000010;
      patterns[42008] = 29'b1_010010000011_000_1_010010000011;
      patterns[42009] = 29'b1_010010000011_001_1_000011010010;
      patterns[42010] = 29'b1_010010000011_010_0_100100000111;
      patterns[42011] = 29'b1_010010000011_011_1_001000001110;
      patterns[42012] = 29'b1_010010000011_100_1_101001000001;
      patterns[42013] = 29'b1_010010000011_101_1_110100100000;
      patterns[42014] = 29'b1_010010000011_110_1_010010000011;
      patterns[42015] = 29'b1_010010000011_111_1_010010000011;
      patterns[42016] = 29'b1_010010000100_000_1_010010000100;
      patterns[42017] = 29'b1_010010000100_001_1_000100010010;
      patterns[42018] = 29'b1_010010000100_010_0_100100001001;
      patterns[42019] = 29'b1_010010000100_011_1_001000010010;
      patterns[42020] = 29'b1_010010000100_100_0_101001000010;
      patterns[42021] = 29'b1_010010000100_101_0_010100100001;
      patterns[42022] = 29'b1_010010000100_110_1_010010000100;
      patterns[42023] = 29'b1_010010000100_111_1_010010000100;
      patterns[42024] = 29'b1_010010000101_000_1_010010000101;
      patterns[42025] = 29'b1_010010000101_001_1_000101010010;
      patterns[42026] = 29'b1_010010000101_010_0_100100001011;
      patterns[42027] = 29'b1_010010000101_011_1_001000010110;
      patterns[42028] = 29'b1_010010000101_100_1_101001000010;
      patterns[42029] = 29'b1_010010000101_101_0_110100100001;
      patterns[42030] = 29'b1_010010000101_110_1_010010000101;
      patterns[42031] = 29'b1_010010000101_111_1_010010000101;
      patterns[42032] = 29'b1_010010000110_000_1_010010000110;
      patterns[42033] = 29'b1_010010000110_001_1_000110010010;
      patterns[42034] = 29'b1_010010000110_010_0_100100001101;
      patterns[42035] = 29'b1_010010000110_011_1_001000011010;
      patterns[42036] = 29'b1_010010000110_100_0_101001000011;
      patterns[42037] = 29'b1_010010000110_101_1_010100100001;
      patterns[42038] = 29'b1_010010000110_110_1_010010000110;
      patterns[42039] = 29'b1_010010000110_111_1_010010000110;
      patterns[42040] = 29'b1_010010000111_000_1_010010000111;
      patterns[42041] = 29'b1_010010000111_001_1_000111010010;
      patterns[42042] = 29'b1_010010000111_010_0_100100001111;
      patterns[42043] = 29'b1_010010000111_011_1_001000011110;
      patterns[42044] = 29'b1_010010000111_100_1_101001000011;
      patterns[42045] = 29'b1_010010000111_101_1_110100100001;
      patterns[42046] = 29'b1_010010000111_110_1_010010000111;
      patterns[42047] = 29'b1_010010000111_111_1_010010000111;
      patterns[42048] = 29'b1_010010001000_000_1_010010001000;
      patterns[42049] = 29'b1_010010001000_001_1_001000010010;
      patterns[42050] = 29'b1_010010001000_010_0_100100010001;
      patterns[42051] = 29'b1_010010001000_011_1_001000100010;
      patterns[42052] = 29'b1_010010001000_100_0_101001000100;
      patterns[42053] = 29'b1_010010001000_101_0_010100100010;
      patterns[42054] = 29'b1_010010001000_110_1_010010001000;
      patterns[42055] = 29'b1_010010001000_111_1_010010001000;
      patterns[42056] = 29'b1_010010001001_000_1_010010001001;
      patterns[42057] = 29'b1_010010001001_001_1_001001010010;
      patterns[42058] = 29'b1_010010001001_010_0_100100010011;
      patterns[42059] = 29'b1_010010001001_011_1_001000100110;
      patterns[42060] = 29'b1_010010001001_100_1_101001000100;
      patterns[42061] = 29'b1_010010001001_101_0_110100100010;
      patterns[42062] = 29'b1_010010001001_110_1_010010001001;
      patterns[42063] = 29'b1_010010001001_111_1_010010001001;
      patterns[42064] = 29'b1_010010001010_000_1_010010001010;
      patterns[42065] = 29'b1_010010001010_001_1_001010010010;
      patterns[42066] = 29'b1_010010001010_010_0_100100010101;
      patterns[42067] = 29'b1_010010001010_011_1_001000101010;
      patterns[42068] = 29'b1_010010001010_100_0_101001000101;
      patterns[42069] = 29'b1_010010001010_101_1_010100100010;
      patterns[42070] = 29'b1_010010001010_110_1_010010001010;
      patterns[42071] = 29'b1_010010001010_111_1_010010001010;
      patterns[42072] = 29'b1_010010001011_000_1_010010001011;
      patterns[42073] = 29'b1_010010001011_001_1_001011010010;
      patterns[42074] = 29'b1_010010001011_010_0_100100010111;
      patterns[42075] = 29'b1_010010001011_011_1_001000101110;
      patterns[42076] = 29'b1_010010001011_100_1_101001000101;
      patterns[42077] = 29'b1_010010001011_101_1_110100100010;
      patterns[42078] = 29'b1_010010001011_110_1_010010001011;
      patterns[42079] = 29'b1_010010001011_111_1_010010001011;
      patterns[42080] = 29'b1_010010001100_000_1_010010001100;
      patterns[42081] = 29'b1_010010001100_001_1_001100010010;
      patterns[42082] = 29'b1_010010001100_010_0_100100011001;
      patterns[42083] = 29'b1_010010001100_011_1_001000110010;
      patterns[42084] = 29'b1_010010001100_100_0_101001000110;
      patterns[42085] = 29'b1_010010001100_101_0_010100100011;
      patterns[42086] = 29'b1_010010001100_110_1_010010001100;
      patterns[42087] = 29'b1_010010001100_111_1_010010001100;
      patterns[42088] = 29'b1_010010001101_000_1_010010001101;
      patterns[42089] = 29'b1_010010001101_001_1_001101010010;
      patterns[42090] = 29'b1_010010001101_010_0_100100011011;
      patterns[42091] = 29'b1_010010001101_011_1_001000110110;
      patterns[42092] = 29'b1_010010001101_100_1_101001000110;
      patterns[42093] = 29'b1_010010001101_101_0_110100100011;
      patterns[42094] = 29'b1_010010001101_110_1_010010001101;
      patterns[42095] = 29'b1_010010001101_111_1_010010001101;
      patterns[42096] = 29'b1_010010001110_000_1_010010001110;
      patterns[42097] = 29'b1_010010001110_001_1_001110010010;
      patterns[42098] = 29'b1_010010001110_010_0_100100011101;
      patterns[42099] = 29'b1_010010001110_011_1_001000111010;
      patterns[42100] = 29'b1_010010001110_100_0_101001000111;
      patterns[42101] = 29'b1_010010001110_101_1_010100100011;
      patterns[42102] = 29'b1_010010001110_110_1_010010001110;
      patterns[42103] = 29'b1_010010001110_111_1_010010001110;
      patterns[42104] = 29'b1_010010001111_000_1_010010001111;
      patterns[42105] = 29'b1_010010001111_001_1_001111010010;
      patterns[42106] = 29'b1_010010001111_010_0_100100011111;
      patterns[42107] = 29'b1_010010001111_011_1_001000111110;
      patterns[42108] = 29'b1_010010001111_100_1_101001000111;
      patterns[42109] = 29'b1_010010001111_101_1_110100100011;
      patterns[42110] = 29'b1_010010001111_110_1_010010001111;
      patterns[42111] = 29'b1_010010001111_111_1_010010001111;
      patterns[42112] = 29'b1_010010010000_000_1_010010010000;
      patterns[42113] = 29'b1_010010010000_001_1_010000010010;
      patterns[42114] = 29'b1_010010010000_010_0_100100100001;
      patterns[42115] = 29'b1_010010010000_011_1_001001000010;
      patterns[42116] = 29'b1_010010010000_100_0_101001001000;
      patterns[42117] = 29'b1_010010010000_101_0_010100100100;
      patterns[42118] = 29'b1_010010010000_110_1_010010010000;
      patterns[42119] = 29'b1_010010010000_111_1_010010010000;
      patterns[42120] = 29'b1_010010010001_000_1_010010010001;
      patterns[42121] = 29'b1_010010010001_001_1_010001010010;
      patterns[42122] = 29'b1_010010010001_010_0_100100100011;
      patterns[42123] = 29'b1_010010010001_011_1_001001000110;
      patterns[42124] = 29'b1_010010010001_100_1_101001001000;
      patterns[42125] = 29'b1_010010010001_101_0_110100100100;
      patterns[42126] = 29'b1_010010010001_110_1_010010010001;
      patterns[42127] = 29'b1_010010010001_111_1_010010010001;
      patterns[42128] = 29'b1_010010010010_000_1_010010010010;
      patterns[42129] = 29'b1_010010010010_001_1_010010010010;
      patterns[42130] = 29'b1_010010010010_010_0_100100100101;
      patterns[42131] = 29'b1_010010010010_011_1_001001001010;
      patterns[42132] = 29'b1_010010010010_100_0_101001001001;
      patterns[42133] = 29'b1_010010010010_101_1_010100100100;
      patterns[42134] = 29'b1_010010010010_110_1_010010010010;
      patterns[42135] = 29'b1_010010010010_111_1_010010010010;
      patterns[42136] = 29'b1_010010010011_000_1_010010010011;
      patterns[42137] = 29'b1_010010010011_001_1_010011010010;
      patterns[42138] = 29'b1_010010010011_010_0_100100100111;
      patterns[42139] = 29'b1_010010010011_011_1_001001001110;
      patterns[42140] = 29'b1_010010010011_100_1_101001001001;
      patterns[42141] = 29'b1_010010010011_101_1_110100100100;
      patterns[42142] = 29'b1_010010010011_110_1_010010010011;
      patterns[42143] = 29'b1_010010010011_111_1_010010010011;
      patterns[42144] = 29'b1_010010010100_000_1_010010010100;
      patterns[42145] = 29'b1_010010010100_001_1_010100010010;
      patterns[42146] = 29'b1_010010010100_010_0_100100101001;
      patterns[42147] = 29'b1_010010010100_011_1_001001010010;
      patterns[42148] = 29'b1_010010010100_100_0_101001001010;
      patterns[42149] = 29'b1_010010010100_101_0_010100100101;
      patterns[42150] = 29'b1_010010010100_110_1_010010010100;
      patterns[42151] = 29'b1_010010010100_111_1_010010010100;
      patterns[42152] = 29'b1_010010010101_000_1_010010010101;
      patterns[42153] = 29'b1_010010010101_001_1_010101010010;
      patterns[42154] = 29'b1_010010010101_010_0_100100101011;
      patterns[42155] = 29'b1_010010010101_011_1_001001010110;
      patterns[42156] = 29'b1_010010010101_100_1_101001001010;
      patterns[42157] = 29'b1_010010010101_101_0_110100100101;
      patterns[42158] = 29'b1_010010010101_110_1_010010010101;
      patterns[42159] = 29'b1_010010010101_111_1_010010010101;
      patterns[42160] = 29'b1_010010010110_000_1_010010010110;
      patterns[42161] = 29'b1_010010010110_001_1_010110010010;
      patterns[42162] = 29'b1_010010010110_010_0_100100101101;
      patterns[42163] = 29'b1_010010010110_011_1_001001011010;
      patterns[42164] = 29'b1_010010010110_100_0_101001001011;
      patterns[42165] = 29'b1_010010010110_101_1_010100100101;
      patterns[42166] = 29'b1_010010010110_110_1_010010010110;
      patterns[42167] = 29'b1_010010010110_111_1_010010010110;
      patterns[42168] = 29'b1_010010010111_000_1_010010010111;
      patterns[42169] = 29'b1_010010010111_001_1_010111010010;
      patterns[42170] = 29'b1_010010010111_010_0_100100101111;
      patterns[42171] = 29'b1_010010010111_011_1_001001011110;
      patterns[42172] = 29'b1_010010010111_100_1_101001001011;
      patterns[42173] = 29'b1_010010010111_101_1_110100100101;
      patterns[42174] = 29'b1_010010010111_110_1_010010010111;
      patterns[42175] = 29'b1_010010010111_111_1_010010010111;
      patterns[42176] = 29'b1_010010011000_000_1_010010011000;
      patterns[42177] = 29'b1_010010011000_001_1_011000010010;
      patterns[42178] = 29'b1_010010011000_010_0_100100110001;
      patterns[42179] = 29'b1_010010011000_011_1_001001100010;
      patterns[42180] = 29'b1_010010011000_100_0_101001001100;
      patterns[42181] = 29'b1_010010011000_101_0_010100100110;
      patterns[42182] = 29'b1_010010011000_110_1_010010011000;
      patterns[42183] = 29'b1_010010011000_111_1_010010011000;
      patterns[42184] = 29'b1_010010011001_000_1_010010011001;
      patterns[42185] = 29'b1_010010011001_001_1_011001010010;
      patterns[42186] = 29'b1_010010011001_010_0_100100110011;
      patterns[42187] = 29'b1_010010011001_011_1_001001100110;
      patterns[42188] = 29'b1_010010011001_100_1_101001001100;
      patterns[42189] = 29'b1_010010011001_101_0_110100100110;
      patterns[42190] = 29'b1_010010011001_110_1_010010011001;
      patterns[42191] = 29'b1_010010011001_111_1_010010011001;
      patterns[42192] = 29'b1_010010011010_000_1_010010011010;
      patterns[42193] = 29'b1_010010011010_001_1_011010010010;
      patterns[42194] = 29'b1_010010011010_010_0_100100110101;
      patterns[42195] = 29'b1_010010011010_011_1_001001101010;
      patterns[42196] = 29'b1_010010011010_100_0_101001001101;
      patterns[42197] = 29'b1_010010011010_101_1_010100100110;
      patterns[42198] = 29'b1_010010011010_110_1_010010011010;
      patterns[42199] = 29'b1_010010011010_111_1_010010011010;
      patterns[42200] = 29'b1_010010011011_000_1_010010011011;
      patterns[42201] = 29'b1_010010011011_001_1_011011010010;
      patterns[42202] = 29'b1_010010011011_010_0_100100110111;
      patterns[42203] = 29'b1_010010011011_011_1_001001101110;
      patterns[42204] = 29'b1_010010011011_100_1_101001001101;
      patterns[42205] = 29'b1_010010011011_101_1_110100100110;
      patterns[42206] = 29'b1_010010011011_110_1_010010011011;
      patterns[42207] = 29'b1_010010011011_111_1_010010011011;
      patterns[42208] = 29'b1_010010011100_000_1_010010011100;
      patterns[42209] = 29'b1_010010011100_001_1_011100010010;
      patterns[42210] = 29'b1_010010011100_010_0_100100111001;
      patterns[42211] = 29'b1_010010011100_011_1_001001110010;
      patterns[42212] = 29'b1_010010011100_100_0_101001001110;
      patterns[42213] = 29'b1_010010011100_101_0_010100100111;
      patterns[42214] = 29'b1_010010011100_110_1_010010011100;
      patterns[42215] = 29'b1_010010011100_111_1_010010011100;
      patterns[42216] = 29'b1_010010011101_000_1_010010011101;
      patterns[42217] = 29'b1_010010011101_001_1_011101010010;
      patterns[42218] = 29'b1_010010011101_010_0_100100111011;
      patterns[42219] = 29'b1_010010011101_011_1_001001110110;
      patterns[42220] = 29'b1_010010011101_100_1_101001001110;
      patterns[42221] = 29'b1_010010011101_101_0_110100100111;
      patterns[42222] = 29'b1_010010011101_110_1_010010011101;
      patterns[42223] = 29'b1_010010011101_111_1_010010011101;
      patterns[42224] = 29'b1_010010011110_000_1_010010011110;
      patterns[42225] = 29'b1_010010011110_001_1_011110010010;
      patterns[42226] = 29'b1_010010011110_010_0_100100111101;
      patterns[42227] = 29'b1_010010011110_011_1_001001111010;
      patterns[42228] = 29'b1_010010011110_100_0_101001001111;
      patterns[42229] = 29'b1_010010011110_101_1_010100100111;
      patterns[42230] = 29'b1_010010011110_110_1_010010011110;
      patterns[42231] = 29'b1_010010011110_111_1_010010011110;
      patterns[42232] = 29'b1_010010011111_000_1_010010011111;
      patterns[42233] = 29'b1_010010011111_001_1_011111010010;
      patterns[42234] = 29'b1_010010011111_010_0_100100111111;
      patterns[42235] = 29'b1_010010011111_011_1_001001111110;
      patterns[42236] = 29'b1_010010011111_100_1_101001001111;
      patterns[42237] = 29'b1_010010011111_101_1_110100100111;
      patterns[42238] = 29'b1_010010011111_110_1_010010011111;
      patterns[42239] = 29'b1_010010011111_111_1_010010011111;
      patterns[42240] = 29'b1_010010100000_000_1_010010100000;
      patterns[42241] = 29'b1_010010100000_001_1_100000010010;
      patterns[42242] = 29'b1_010010100000_010_0_100101000001;
      patterns[42243] = 29'b1_010010100000_011_1_001010000010;
      patterns[42244] = 29'b1_010010100000_100_0_101001010000;
      patterns[42245] = 29'b1_010010100000_101_0_010100101000;
      patterns[42246] = 29'b1_010010100000_110_1_010010100000;
      patterns[42247] = 29'b1_010010100000_111_1_010010100000;
      patterns[42248] = 29'b1_010010100001_000_1_010010100001;
      patterns[42249] = 29'b1_010010100001_001_1_100001010010;
      patterns[42250] = 29'b1_010010100001_010_0_100101000011;
      patterns[42251] = 29'b1_010010100001_011_1_001010000110;
      patterns[42252] = 29'b1_010010100001_100_1_101001010000;
      patterns[42253] = 29'b1_010010100001_101_0_110100101000;
      patterns[42254] = 29'b1_010010100001_110_1_010010100001;
      patterns[42255] = 29'b1_010010100001_111_1_010010100001;
      patterns[42256] = 29'b1_010010100010_000_1_010010100010;
      patterns[42257] = 29'b1_010010100010_001_1_100010010010;
      patterns[42258] = 29'b1_010010100010_010_0_100101000101;
      patterns[42259] = 29'b1_010010100010_011_1_001010001010;
      patterns[42260] = 29'b1_010010100010_100_0_101001010001;
      patterns[42261] = 29'b1_010010100010_101_1_010100101000;
      patterns[42262] = 29'b1_010010100010_110_1_010010100010;
      patterns[42263] = 29'b1_010010100010_111_1_010010100010;
      patterns[42264] = 29'b1_010010100011_000_1_010010100011;
      patterns[42265] = 29'b1_010010100011_001_1_100011010010;
      patterns[42266] = 29'b1_010010100011_010_0_100101000111;
      patterns[42267] = 29'b1_010010100011_011_1_001010001110;
      patterns[42268] = 29'b1_010010100011_100_1_101001010001;
      patterns[42269] = 29'b1_010010100011_101_1_110100101000;
      patterns[42270] = 29'b1_010010100011_110_1_010010100011;
      patterns[42271] = 29'b1_010010100011_111_1_010010100011;
      patterns[42272] = 29'b1_010010100100_000_1_010010100100;
      patterns[42273] = 29'b1_010010100100_001_1_100100010010;
      patterns[42274] = 29'b1_010010100100_010_0_100101001001;
      patterns[42275] = 29'b1_010010100100_011_1_001010010010;
      patterns[42276] = 29'b1_010010100100_100_0_101001010010;
      patterns[42277] = 29'b1_010010100100_101_0_010100101001;
      patterns[42278] = 29'b1_010010100100_110_1_010010100100;
      patterns[42279] = 29'b1_010010100100_111_1_010010100100;
      patterns[42280] = 29'b1_010010100101_000_1_010010100101;
      patterns[42281] = 29'b1_010010100101_001_1_100101010010;
      patterns[42282] = 29'b1_010010100101_010_0_100101001011;
      patterns[42283] = 29'b1_010010100101_011_1_001010010110;
      patterns[42284] = 29'b1_010010100101_100_1_101001010010;
      patterns[42285] = 29'b1_010010100101_101_0_110100101001;
      patterns[42286] = 29'b1_010010100101_110_1_010010100101;
      patterns[42287] = 29'b1_010010100101_111_1_010010100101;
      patterns[42288] = 29'b1_010010100110_000_1_010010100110;
      patterns[42289] = 29'b1_010010100110_001_1_100110010010;
      patterns[42290] = 29'b1_010010100110_010_0_100101001101;
      patterns[42291] = 29'b1_010010100110_011_1_001010011010;
      patterns[42292] = 29'b1_010010100110_100_0_101001010011;
      patterns[42293] = 29'b1_010010100110_101_1_010100101001;
      patterns[42294] = 29'b1_010010100110_110_1_010010100110;
      patterns[42295] = 29'b1_010010100110_111_1_010010100110;
      patterns[42296] = 29'b1_010010100111_000_1_010010100111;
      patterns[42297] = 29'b1_010010100111_001_1_100111010010;
      patterns[42298] = 29'b1_010010100111_010_0_100101001111;
      patterns[42299] = 29'b1_010010100111_011_1_001010011110;
      patterns[42300] = 29'b1_010010100111_100_1_101001010011;
      patterns[42301] = 29'b1_010010100111_101_1_110100101001;
      patterns[42302] = 29'b1_010010100111_110_1_010010100111;
      patterns[42303] = 29'b1_010010100111_111_1_010010100111;
      patterns[42304] = 29'b1_010010101000_000_1_010010101000;
      patterns[42305] = 29'b1_010010101000_001_1_101000010010;
      patterns[42306] = 29'b1_010010101000_010_0_100101010001;
      patterns[42307] = 29'b1_010010101000_011_1_001010100010;
      patterns[42308] = 29'b1_010010101000_100_0_101001010100;
      patterns[42309] = 29'b1_010010101000_101_0_010100101010;
      patterns[42310] = 29'b1_010010101000_110_1_010010101000;
      patterns[42311] = 29'b1_010010101000_111_1_010010101000;
      patterns[42312] = 29'b1_010010101001_000_1_010010101001;
      patterns[42313] = 29'b1_010010101001_001_1_101001010010;
      patterns[42314] = 29'b1_010010101001_010_0_100101010011;
      patterns[42315] = 29'b1_010010101001_011_1_001010100110;
      patterns[42316] = 29'b1_010010101001_100_1_101001010100;
      patterns[42317] = 29'b1_010010101001_101_0_110100101010;
      patterns[42318] = 29'b1_010010101001_110_1_010010101001;
      patterns[42319] = 29'b1_010010101001_111_1_010010101001;
      patterns[42320] = 29'b1_010010101010_000_1_010010101010;
      patterns[42321] = 29'b1_010010101010_001_1_101010010010;
      patterns[42322] = 29'b1_010010101010_010_0_100101010101;
      patterns[42323] = 29'b1_010010101010_011_1_001010101010;
      patterns[42324] = 29'b1_010010101010_100_0_101001010101;
      patterns[42325] = 29'b1_010010101010_101_1_010100101010;
      patterns[42326] = 29'b1_010010101010_110_1_010010101010;
      patterns[42327] = 29'b1_010010101010_111_1_010010101010;
      patterns[42328] = 29'b1_010010101011_000_1_010010101011;
      patterns[42329] = 29'b1_010010101011_001_1_101011010010;
      patterns[42330] = 29'b1_010010101011_010_0_100101010111;
      patterns[42331] = 29'b1_010010101011_011_1_001010101110;
      patterns[42332] = 29'b1_010010101011_100_1_101001010101;
      patterns[42333] = 29'b1_010010101011_101_1_110100101010;
      patterns[42334] = 29'b1_010010101011_110_1_010010101011;
      patterns[42335] = 29'b1_010010101011_111_1_010010101011;
      patterns[42336] = 29'b1_010010101100_000_1_010010101100;
      patterns[42337] = 29'b1_010010101100_001_1_101100010010;
      patterns[42338] = 29'b1_010010101100_010_0_100101011001;
      patterns[42339] = 29'b1_010010101100_011_1_001010110010;
      patterns[42340] = 29'b1_010010101100_100_0_101001010110;
      patterns[42341] = 29'b1_010010101100_101_0_010100101011;
      patterns[42342] = 29'b1_010010101100_110_1_010010101100;
      patterns[42343] = 29'b1_010010101100_111_1_010010101100;
      patterns[42344] = 29'b1_010010101101_000_1_010010101101;
      patterns[42345] = 29'b1_010010101101_001_1_101101010010;
      patterns[42346] = 29'b1_010010101101_010_0_100101011011;
      patterns[42347] = 29'b1_010010101101_011_1_001010110110;
      patterns[42348] = 29'b1_010010101101_100_1_101001010110;
      patterns[42349] = 29'b1_010010101101_101_0_110100101011;
      patterns[42350] = 29'b1_010010101101_110_1_010010101101;
      patterns[42351] = 29'b1_010010101101_111_1_010010101101;
      patterns[42352] = 29'b1_010010101110_000_1_010010101110;
      patterns[42353] = 29'b1_010010101110_001_1_101110010010;
      patterns[42354] = 29'b1_010010101110_010_0_100101011101;
      patterns[42355] = 29'b1_010010101110_011_1_001010111010;
      patterns[42356] = 29'b1_010010101110_100_0_101001010111;
      patterns[42357] = 29'b1_010010101110_101_1_010100101011;
      patterns[42358] = 29'b1_010010101110_110_1_010010101110;
      patterns[42359] = 29'b1_010010101110_111_1_010010101110;
      patterns[42360] = 29'b1_010010101111_000_1_010010101111;
      patterns[42361] = 29'b1_010010101111_001_1_101111010010;
      patterns[42362] = 29'b1_010010101111_010_0_100101011111;
      patterns[42363] = 29'b1_010010101111_011_1_001010111110;
      patterns[42364] = 29'b1_010010101111_100_1_101001010111;
      patterns[42365] = 29'b1_010010101111_101_1_110100101011;
      patterns[42366] = 29'b1_010010101111_110_1_010010101111;
      patterns[42367] = 29'b1_010010101111_111_1_010010101111;
      patterns[42368] = 29'b1_010010110000_000_1_010010110000;
      patterns[42369] = 29'b1_010010110000_001_1_110000010010;
      patterns[42370] = 29'b1_010010110000_010_0_100101100001;
      patterns[42371] = 29'b1_010010110000_011_1_001011000010;
      patterns[42372] = 29'b1_010010110000_100_0_101001011000;
      patterns[42373] = 29'b1_010010110000_101_0_010100101100;
      patterns[42374] = 29'b1_010010110000_110_1_010010110000;
      patterns[42375] = 29'b1_010010110000_111_1_010010110000;
      patterns[42376] = 29'b1_010010110001_000_1_010010110001;
      patterns[42377] = 29'b1_010010110001_001_1_110001010010;
      patterns[42378] = 29'b1_010010110001_010_0_100101100011;
      patterns[42379] = 29'b1_010010110001_011_1_001011000110;
      patterns[42380] = 29'b1_010010110001_100_1_101001011000;
      patterns[42381] = 29'b1_010010110001_101_0_110100101100;
      patterns[42382] = 29'b1_010010110001_110_1_010010110001;
      patterns[42383] = 29'b1_010010110001_111_1_010010110001;
      patterns[42384] = 29'b1_010010110010_000_1_010010110010;
      patterns[42385] = 29'b1_010010110010_001_1_110010010010;
      patterns[42386] = 29'b1_010010110010_010_0_100101100101;
      patterns[42387] = 29'b1_010010110010_011_1_001011001010;
      patterns[42388] = 29'b1_010010110010_100_0_101001011001;
      patterns[42389] = 29'b1_010010110010_101_1_010100101100;
      patterns[42390] = 29'b1_010010110010_110_1_010010110010;
      patterns[42391] = 29'b1_010010110010_111_1_010010110010;
      patterns[42392] = 29'b1_010010110011_000_1_010010110011;
      patterns[42393] = 29'b1_010010110011_001_1_110011010010;
      patterns[42394] = 29'b1_010010110011_010_0_100101100111;
      patterns[42395] = 29'b1_010010110011_011_1_001011001110;
      patterns[42396] = 29'b1_010010110011_100_1_101001011001;
      patterns[42397] = 29'b1_010010110011_101_1_110100101100;
      patterns[42398] = 29'b1_010010110011_110_1_010010110011;
      patterns[42399] = 29'b1_010010110011_111_1_010010110011;
      patterns[42400] = 29'b1_010010110100_000_1_010010110100;
      patterns[42401] = 29'b1_010010110100_001_1_110100010010;
      patterns[42402] = 29'b1_010010110100_010_0_100101101001;
      patterns[42403] = 29'b1_010010110100_011_1_001011010010;
      patterns[42404] = 29'b1_010010110100_100_0_101001011010;
      patterns[42405] = 29'b1_010010110100_101_0_010100101101;
      patterns[42406] = 29'b1_010010110100_110_1_010010110100;
      patterns[42407] = 29'b1_010010110100_111_1_010010110100;
      patterns[42408] = 29'b1_010010110101_000_1_010010110101;
      patterns[42409] = 29'b1_010010110101_001_1_110101010010;
      patterns[42410] = 29'b1_010010110101_010_0_100101101011;
      patterns[42411] = 29'b1_010010110101_011_1_001011010110;
      patterns[42412] = 29'b1_010010110101_100_1_101001011010;
      patterns[42413] = 29'b1_010010110101_101_0_110100101101;
      patterns[42414] = 29'b1_010010110101_110_1_010010110101;
      patterns[42415] = 29'b1_010010110101_111_1_010010110101;
      patterns[42416] = 29'b1_010010110110_000_1_010010110110;
      patterns[42417] = 29'b1_010010110110_001_1_110110010010;
      patterns[42418] = 29'b1_010010110110_010_0_100101101101;
      patterns[42419] = 29'b1_010010110110_011_1_001011011010;
      patterns[42420] = 29'b1_010010110110_100_0_101001011011;
      patterns[42421] = 29'b1_010010110110_101_1_010100101101;
      patterns[42422] = 29'b1_010010110110_110_1_010010110110;
      patterns[42423] = 29'b1_010010110110_111_1_010010110110;
      patterns[42424] = 29'b1_010010110111_000_1_010010110111;
      patterns[42425] = 29'b1_010010110111_001_1_110111010010;
      patterns[42426] = 29'b1_010010110111_010_0_100101101111;
      patterns[42427] = 29'b1_010010110111_011_1_001011011110;
      patterns[42428] = 29'b1_010010110111_100_1_101001011011;
      patterns[42429] = 29'b1_010010110111_101_1_110100101101;
      patterns[42430] = 29'b1_010010110111_110_1_010010110111;
      patterns[42431] = 29'b1_010010110111_111_1_010010110111;
      patterns[42432] = 29'b1_010010111000_000_1_010010111000;
      patterns[42433] = 29'b1_010010111000_001_1_111000010010;
      patterns[42434] = 29'b1_010010111000_010_0_100101110001;
      patterns[42435] = 29'b1_010010111000_011_1_001011100010;
      patterns[42436] = 29'b1_010010111000_100_0_101001011100;
      patterns[42437] = 29'b1_010010111000_101_0_010100101110;
      patterns[42438] = 29'b1_010010111000_110_1_010010111000;
      patterns[42439] = 29'b1_010010111000_111_1_010010111000;
      patterns[42440] = 29'b1_010010111001_000_1_010010111001;
      patterns[42441] = 29'b1_010010111001_001_1_111001010010;
      patterns[42442] = 29'b1_010010111001_010_0_100101110011;
      patterns[42443] = 29'b1_010010111001_011_1_001011100110;
      patterns[42444] = 29'b1_010010111001_100_1_101001011100;
      patterns[42445] = 29'b1_010010111001_101_0_110100101110;
      patterns[42446] = 29'b1_010010111001_110_1_010010111001;
      patterns[42447] = 29'b1_010010111001_111_1_010010111001;
      patterns[42448] = 29'b1_010010111010_000_1_010010111010;
      patterns[42449] = 29'b1_010010111010_001_1_111010010010;
      patterns[42450] = 29'b1_010010111010_010_0_100101110101;
      patterns[42451] = 29'b1_010010111010_011_1_001011101010;
      patterns[42452] = 29'b1_010010111010_100_0_101001011101;
      patterns[42453] = 29'b1_010010111010_101_1_010100101110;
      patterns[42454] = 29'b1_010010111010_110_1_010010111010;
      patterns[42455] = 29'b1_010010111010_111_1_010010111010;
      patterns[42456] = 29'b1_010010111011_000_1_010010111011;
      patterns[42457] = 29'b1_010010111011_001_1_111011010010;
      patterns[42458] = 29'b1_010010111011_010_0_100101110111;
      patterns[42459] = 29'b1_010010111011_011_1_001011101110;
      patterns[42460] = 29'b1_010010111011_100_1_101001011101;
      patterns[42461] = 29'b1_010010111011_101_1_110100101110;
      patterns[42462] = 29'b1_010010111011_110_1_010010111011;
      patterns[42463] = 29'b1_010010111011_111_1_010010111011;
      patterns[42464] = 29'b1_010010111100_000_1_010010111100;
      patterns[42465] = 29'b1_010010111100_001_1_111100010010;
      patterns[42466] = 29'b1_010010111100_010_0_100101111001;
      patterns[42467] = 29'b1_010010111100_011_1_001011110010;
      patterns[42468] = 29'b1_010010111100_100_0_101001011110;
      patterns[42469] = 29'b1_010010111100_101_0_010100101111;
      patterns[42470] = 29'b1_010010111100_110_1_010010111100;
      patterns[42471] = 29'b1_010010111100_111_1_010010111100;
      patterns[42472] = 29'b1_010010111101_000_1_010010111101;
      patterns[42473] = 29'b1_010010111101_001_1_111101010010;
      patterns[42474] = 29'b1_010010111101_010_0_100101111011;
      patterns[42475] = 29'b1_010010111101_011_1_001011110110;
      patterns[42476] = 29'b1_010010111101_100_1_101001011110;
      patterns[42477] = 29'b1_010010111101_101_0_110100101111;
      patterns[42478] = 29'b1_010010111101_110_1_010010111101;
      patterns[42479] = 29'b1_010010111101_111_1_010010111101;
      patterns[42480] = 29'b1_010010111110_000_1_010010111110;
      patterns[42481] = 29'b1_010010111110_001_1_111110010010;
      patterns[42482] = 29'b1_010010111110_010_0_100101111101;
      patterns[42483] = 29'b1_010010111110_011_1_001011111010;
      patterns[42484] = 29'b1_010010111110_100_0_101001011111;
      patterns[42485] = 29'b1_010010111110_101_1_010100101111;
      patterns[42486] = 29'b1_010010111110_110_1_010010111110;
      patterns[42487] = 29'b1_010010111110_111_1_010010111110;
      patterns[42488] = 29'b1_010010111111_000_1_010010111111;
      patterns[42489] = 29'b1_010010111111_001_1_111111010010;
      patterns[42490] = 29'b1_010010111111_010_0_100101111111;
      patterns[42491] = 29'b1_010010111111_011_1_001011111110;
      patterns[42492] = 29'b1_010010111111_100_1_101001011111;
      patterns[42493] = 29'b1_010010111111_101_1_110100101111;
      patterns[42494] = 29'b1_010010111111_110_1_010010111111;
      patterns[42495] = 29'b1_010010111111_111_1_010010111111;
      patterns[42496] = 29'b1_010011000000_000_1_010011000000;
      patterns[42497] = 29'b1_010011000000_001_1_000000010011;
      patterns[42498] = 29'b1_010011000000_010_0_100110000001;
      patterns[42499] = 29'b1_010011000000_011_1_001100000010;
      patterns[42500] = 29'b1_010011000000_100_0_101001100000;
      patterns[42501] = 29'b1_010011000000_101_0_010100110000;
      patterns[42502] = 29'b1_010011000000_110_1_010011000000;
      patterns[42503] = 29'b1_010011000000_111_1_010011000000;
      patterns[42504] = 29'b1_010011000001_000_1_010011000001;
      patterns[42505] = 29'b1_010011000001_001_1_000001010011;
      patterns[42506] = 29'b1_010011000001_010_0_100110000011;
      patterns[42507] = 29'b1_010011000001_011_1_001100000110;
      patterns[42508] = 29'b1_010011000001_100_1_101001100000;
      patterns[42509] = 29'b1_010011000001_101_0_110100110000;
      patterns[42510] = 29'b1_010011000001_110_1_010011000001;
      patterns[42511] = 29'b1_010011000001_111_1_010011000001;
      patterns[42512] = 29'b1_010011000010_000_1_010011000010;
      patterns[42513] = 29'b1_010011000010_001_1_000010010011;
      patterns[42514] = 29'b1_010011000010_010_0_100110000101;
      patterns[42515] = 29'b1_010011000010_011_1_001100001010;
      patterns[42516] = 29'b1_010011000010_100_0_101001100001;
      patterns[42517] = 29'b1_010011000010_101_1_010100110000;
      patterns[42518] = 29'b1_010011000010_110_1_010011000010;
      patterns[42519] = 29'b1_010011000010_111_1_010011000010;
      patterns[42520] = 29'b1_010011000011_000_1_010011000011;
      patterns[42521] = 29'b1_010011000011_001_1_000011010011;
      patterns[42522] = 29'b1_010011000011_010_0_100110000111;
      patterns[42523] = 29'b1_010011000011_011_1_001100001110;
      patterns[42524] = 29'b1_010011000011_100_1_101001100001;
      patterns[42525] = 29'b1_010011000011_101_1_110100110000;
      patterns[42526] = 29'b1_010011000011_110_1_010011000011;
      patterns[42527] = 29'b1_010011000011_111_1_010011000011;
      patterns[42528] = 29'b1_010011000100_000_1_010011000100;
      patterns[42529] = 29'b1_010011000100_001_1_000100010011;
      patterns[42530] = 29'b1_010011000100_010_0_100110001001;
      patterns[42531] = 29'b1_010011000100_011_1_001100010010;
      patterns[42532] = 29'b1_010011000100_100_0_101001100010;
      patterns[42533] = 29'b1_010011000100_101_0_010100110001;
      patterns[42534] = 29'b1_010011000100_110_1_010011000100;
      patterns[42535] = 29'b1_010011000100_111_1_010011000100;
      patterns[42536] = 29'b1_010011000101_000_1_010011000101;
      patterns[42537] = 29'b1_010011000101_001_1_000101010011;
      patterns[42538] = 29'b1_010011000101_010_0_100110001011;
      patterns[42539] = 29'b1_010011000101_011_1_001100010110;
      patterns[42540] = 29'b1_010011000101_100_1_101001100010;
      patterns[42541] = 29'b1_010011000101_101_0_110100110001;
      patterns[42542] = 29'b1_010011000101_110_1_010011000101;
      patterns[42543] = 29'b1_010011000101_111_1_010011000101;
      patterns[42544] = 29'b1_010011000110_000_1_010011000110;
      patterns[42545] = 29'b1_010011000110_001_1_000110010011;
      patterns[42546] = 29'b1_010011000110_010_0_100110001101;
      patterns[42547] = 29'b1_010011000110_011_1_001100011010;
      patterns[42548] = 29'b1_010011000110_100_0_101001100011;
      patterns[42549] = 29'b1_010011000110_101_1_010100110001;
      patterns[42550] = 29'b1_010011000110_110_1_010011000110;
      patterns[42551] = 29'b1_010011000110_111_1_010011000110;
      patterns[42552] = 29'b1_010011000111_000_1_010011000111;
      patterns[42553] = 29'b1_010011000111_001_1_000111010011;
      patterns[42554] = 29'b1_010011000111_010_0_100110001111;
      patterns[42555] = 29'b1_010011000111_011_1_001100011110;
      patterns[42556] = 29'b1_010011000111_100_1_101001100011;
      patterns[42557] = 29'b1_010011000111_101_1_110100110001;
      patterns[42558] = 29'b1_010011000111_110_1_010011000111;
      patterns[42559] = 29'b1_010011000111_111_1_010011000111;
      patterns[42560] = 29'b1_010011001000_000_1_010011001000;
      patterns[42561] = 29'b1_010011001000_001_1_001000010011;
      patterns[42562] = 29'b1_010011001000_010_0_100110010001;
      patterns[42563] = 29'b1_010011001000_011_1_001100100010;
      patterns[42564] = 29'b1_010011001000_100_0_101001100100;
      patterns[42565] = 29'b1_010011001000_101_0_010100110010;
      patterns[42566] = 29'b1_010011001000_110_1_010011001000;
      patterns[42567] = 29'b1_010011001000_111_1_010011001000;
      patterns[42568] = 29'b1_010011001001_000_1_010011001001;
      patterns[42569] = 29'b1_010011001001_001_1_001001010011;
      patterns[42570] = 29'b1_010011001001_010_0_100110010011;
      patterns[42571] = 29'b1_010011001001_011_1_001100100110;
      patterns[42572] = 29'b1_010011001001_100_1_101001100100;
      patterns[42573] = 29'b1_010011001001_101_0_110100110010;
      patterns[42574] = 29'b1_010011001001_110_1_010011001001;
      patterns[42575] = 29'b1_010011001001_111_1_010011001001;
      patterns[42576] = 29'b1_010011001010_000_1_010011001010;
      patterns[42577] = 29'b1_010011001010_001_1_001010010011;
      patterns[42578] = 29'b1_010011001010_010_0_100110010101;
      patterns[42579] = 29'b1_010011001010_011_1_001100101010;
      patterns[42580] = 29'b1_010011001010_100_0_101001100101;
      patterns[42581] = 29'b1_010011001010_101_1_010100110010;
      patterns[42582] = 29'b1_010011001010_110_1_010011001010;
      patterns[42583] = 29'b1_010011001010_111_1_010011001010;
      patterns[42584] = 29'b1_010011001011_000_1_010011001011;
      patterns[42585] = 29'b1_010011001011_001_1_001011010011;
      patterns[42586] = 29'b1_010011001011_010_0_100110010111;
      patterns[42587] = 29'b1_010011001011_011_1_001100101110;
      patterns[42588] = 29'b1_010011001011_100_1_101001100101;
      patterns[42589] = 29'b1_010011001011_101_1_110100110010;
      patterns[42590] = 29'b1_010011001011_110_1_010011001011;
      patterns[42591] = 29'b1_010011001011_111_1_010011001011;
      patterns[42592] = 29'b1_010011001100_000_1_010011001100;
      patterns[42593] = 29'b1_010011001100_001_1_001100010011;
      patterns[42594] = 29'b1_010011001100_010_0_100110011001;
      patterns[42595] = 29'b1_010011001100_011_1_001100110010;
      patterns[42596] = 29'b1_010011001100_100_0_101001100110;
      patterns[42597] = 29'b1_010011001100_101_0_010100110011;
      patterns[42598] = 29'b1_010011001100_110_1_010011001100;
      patterns[42599] = 29'b1_010011001100_111_1_010011001100;
      patterns[42600] = 29'b1_010011001101_000_1_010011001101;
      patterns[42601] = 29'b1_010011001101_001_1_001101010011;
      patterns[42602] = 29'b1_010011001101_010_0_100110011011;
      patterns[42603] = 29'b1_010011001101_011_1_001100110110;
      patterns[42604] = 29'b1_010011001101_100_1_101001100110;
      patterns[42605] = 29'b1_010011001101_101_0_110100110011;
      patterns[42606] = 29'b1_010011001101_110_1_010011001101;
      patterns[42607] = 29'b1_010011001101_111_1_010011001101;
      patterns[42608] = 29'b1_010011001110_000_1_010011001110;
      patterns[42609] = 29'b1_010011001110_001_1_001110010011;
      patterns[42610] = 29'b1_010011001110_010_0_100110011101;
      patterns[42611] = 29'b1_010011001110_011_1_001100111010;
      patterns[42612] = 29'b1_010011001110_100_0_101001100111;
      patterns[42613] = 29'b1_010011001110_101_1_010100110011;
      patterns[42614] = 29'b1_010011001110_110_1_010011001110;
      patterns[42615] = 29'b1_010011001110_111_1_010011001110;
      patterns[42616] = 29'b1_010011001111_000_1_010011001111;
      patterns[42617] = 29'b1_010011001111_001_1_001111010011;
      patterns[42618] = 29'b1_010011001111_010_0_100110011111;
      patterns[42619] = 29'b1_010011001111_011_1_001100111110;
      patterns[42620] = 29'b1_010011001111_100_1_101001100111;
      patterns[42621] = 29'b1_010011001111_101_1_110100110011;
      patterns[42622] = 29'b1_010011001111_110_1_010011001111;
      patterns[42623] = 29'b1_010011001111_111_1_010011001111;
      patterns[42624] = 29'b1_010011010000_000_1_010011010000;
      patterns[42625] = 29'b1_010011010000_001_1_010000010011;
      patterns[42626] = 29'b1_010011010000_010_0_100110100001;
      patterns[42627] = 29'b1_010011010000_011_1_001101000010;
      patterns[42628] = 29'b1_010011010000_100_0_101001101000;
      patterns[42629] = 29'b1_010011010000_101_0_010100110100;
      patterns[42630] = 29'b1_010011010000_110_1_010011010000;
      patterns[42631] = 29'b1_010011010000_111_1_010011010000;
      patterns[42632] = 29'b1_010011010001_000_1_010011010001;
      patterns[42633] = 29'b1_010011010001_001_1_010001010011;
      patterns[42634] = 29'b1_010011010001_010_0_100110100011;
      patterns[42635] = 29'b1_010011010001_011_1_001101000110;
      patterns[42636] = 29'b1_010011010001_100_1_101001101000;
      patterns[42637] = 29'b1_010011010001_101_0_110100110100;
      patterns[42638] = 29'b1_010011010001_110_1_010011010001;
      patterns[42639] = 29'b1_010011010001_111_1_010011010001;
      patterns[42640] = 29'b1_010011010010_000_1_010011010010;
      patterns[42641] = 29'b1_010011010010_001_1_010010010011;
      patterns[42642] = 29'b1_010011010010_010_0_100110100101;
      patterns[42643] = 29'b1_010011010010_011_1_001101001010;
      patterns[42644] = 29'b1_010011010010_100_0_101001101001;
      patterns[42645] = 29'b1_010011010010_101_1_010100110100;
      patterns[42646] = 29'b1_010011010010_110_1_010011010010;
      patterns[42647] = 29'b1_010011010010_111_1_010011010010;
      patterns[42648] = 29'b1_010011010011_000_1_010011010011;
      patterns[42649] = 29'b1_010011010011_001_1_010011010011;
      patterns[42650] = 29'b1_010011010011_010_0_100110100111;
      patterns[42651] = 29'b1_010011010011_011_1_001101001110;
      patterns[42652] = 29'b1_010011010011_100_1_101001101001;
      patterns[42653] = 29'b1_010011010011_101_1_110100110100;
      patterns[42654] = 29'b1_010011010011_110_1_010011010011;
      patterns[42655] = 29'b1_010011010011_111_1_010011010011;
      patterns[42656] = 29'b1_010011010100_000_1_010011010100;
      patterns[42657] = 29'b1_010011010100_001_1_010100010011;
      patterns[42658] = 29'b1_010011010100_010_0_100110101001;
      patterns[42659] = 29'b1_010011010100_011_1_001101010010;
      patterns[42660] = 29'b1_010011010100_100_0_101001101010;
      patterns[42661] = 29'b1_010011010100_101_0_010100110101;
      patterns[42662] = 29'b1_010011010100_110_1_010011010100;
      patterns[42663] = 29'b1_010011010100_111_1_010011010100;
      patterns[42664] = 29'b1_010011010101_000_1_010011010101;
      patterns[42665] = 29'b1_010011010101_001_1_010101010011;
      patterns[42666] = 29'b1_010011010101_010_0_100110101011;
      patterns[42667] = 29'b1_010011010101_011_1_001101010110;
      patterns[42668] = 29'b1_010011010101_100_1_101001101010;
      patterns[42669] = 29'b1_010011010101_101_0_110100110101;
      patterns[42670] = 29'b1_010011010101_110_1_010011010101;
      patterns[42671] = 29'b1_010011010101_111_1_010011010101;
      patterns[42672] = 29'b1_010011010110_000_1_010011010110;
      patterns[42673] = 29'b1_010011010110_001_1_010110010011;
      patterns[42674] = 29'b1_010011010110_010_0_100110101101;
      patterns[42675] = 29'b1_010011010110_011_1_001101011010;
      patterns[42676] = 29'b1_010011010110_100_0_101001101011;
      patterns[42677] = 29'b1_010011010110_101_1_010100110101;
      patterns[42678] = 29'b1_010011010110_110_1_010011010110;
      patterns[42679] = 29'b1_010011010110_111_1_010011010110;
      patterns[42680] = 29'b1_010011010111_000_1_010011010111;
      patterns[42681] = 29'b1_010011010111_001_1_010111010011;
      patterns[42682] = 29'b1_010011010111_010_0_100110101111;
      patterns[42683] = 29'b1_010011010111_011_1_001101011110;
      patterns[42684] = 29'b1_010011010111_100_1_101001101011;
      patterns[42685] = 29'b1_010011010111_101_1_110100110101;
      patterns[42686] = 29'b1_010011010111_110_1_010011010111;
      patterns[42687] = 29'b1_010011010111_111_1_010011010111;
      patterns[42688] = 29'b1_010011011000_000_1_010011011000;
      patterns[42689] = 29'b1_010011011000_001_1_011000010011;
      patterns[42690] = 29'b1_010011011000_010_0_100110110001;
      patterns[42691] = 29'b1_010011011000_011_1_001101100010;
      patterns[42692] = 29'b1_010011011000_100_0_101001101100;
      patterns[42693] = 29'b1_010011011000_101_0_010100110110;
      patterns[42694] = 29'b1_010011011000_110_1_010011011000;
      patterns[42695] = 29'b1_010011011000_111_1_010011011000;
      patterns[42696] = 29'b1_010011011001_000_1_010011011001;
      patterns[42697] = 29'b1_010011011001_001_1_011001010011;
      patterns[42698] = 29'b1_010011011001_010_0_100110110011;
      patterns[42699] = 29'b1_010011011001_011_1_001101100110;
      patterns[42700] = 29'b1_010011011001_100_1_101001101100;
      patterns[42701] = 29'b1_010011011001_101_0_110100110110;
      patterns[42702] = 29'b1_010011011001_110_1_010011011001;
      patterns[42703] = 29'b1_010011011001_111_1_010011011001;
      patterns[42704] = 29'b1_010011011010_000_1_010011011010;
      patterns[42705] = 29'b1_010011011010_001_1_011010010011;
      patterns[42706] = 29'b1_010011011010_010_0_100110110101;
      patterns[42707] = 29'b1_010011011010_011_1_001101101010;
      patterns[42708] = 29'b1_010011011010_100_0_101001101101;
      patterns[42709] = 29'b1_010011011010_101_1_010100110110;
      patterns[42710] = 29'b1_010011011010_110_1_010011011010;
      patterns[42711] = 29'b1_010011011010_111_1_010011011010;
      patterns[42712] = 29'b1_010011011011_000_1_010011011011;
      patterns[42713] = 29'b1_010011011011_001_1_011011010011;
      patterns[42714] = 29'b1_010011011011_010_0_100110110111;
      patterns[42715] = 29'b1_010011011011_011_1_001101101110;
      patterns[42716] = 29'b1_010011011011_100_1_101001101101;
      patterns[42717] = 29'b1_010011011011_101_1_110100110110;
      patterns[42718] = 29'b1_010011011011_110_1_010011011011;
      patterns[42719] = 29'b1_010011011011_111_1_010011011011;
      patterns[42720] = 29'b1_010011011100_000_1_010011011100;
      patterns[42721] = 29'b1_010011011100_001_1_011100010011;
      patterns[42722] = 29'b1_010011011100_010_0_100110111001;
      patterns[42723] = 29'b1_010011011100_011_1_001101110010;
      patterns[42724] = 29'b1_010011011100_100_0_101001101110;
      patterns[42725] = 29'b1_010011011100_101_0_010100110111;
      patterns[42726] = 29'b1_010011011100_110_1_010011011100;
      patterns[42727] = 29'b1_010011011100_111_1_010011011100;
      patterns[42728] = 29'b1_010011011101_000_1_010011011101;
      patterns[42729] = 29'b1_010011011101_001_1_011101010011;
      patterns[42730] = 29'b1_010011011101_010_0_100110111011;
      patterns[42731] = 29'b1_010011011101_011_1_001101110110;
      patterns[42732] = 29'b1_010011011101_100_1_101001101110;
      patterns[42733] = 29'b1_010011011101_101_0_110100110111;
      patterns[42734] = 29'b1_010011011101_110_1_010011011101;
      patterns[42735] = 29'b1_010011011101_111_1_010011011101;
      patterns[42736] = 29'b1_010011011110_000_1_010011011110;
      patterns[42737] = 29'b1_010011011110_001_1_011110010011;
      patterns[42738] = 29'b1_010011011110_010_0_100110111101;
      patterns[42739] = 29'b1_010011011110_011_1_001101111010;
      patterns[42740] = 29'b1_010011011110_100_0_101001101111;
      patterns[42741] = 29'b1_010011011110_101_1_010100110111;
      patterns[42742] = 29'b1_010011011110_110_1_010011011110;
      patterns[42743] = 29'b1_010011011110_111_1_010011011110;
      patterns[42744] = 29'b1_010011011111_000_1_010011011111;
      patterns[42745] = 29'b1_010011011111_001_1_011111010011;
      patterns[42746] = 29'b1_010011011111_010_0_100110111111;
      patterns[42747] = 29'b1_010011011111_011_1_001101111110;
      patterns[42748] = 29'b1_010011011111_100_1_101001101111;
      patterns[42749] = 29'b1_010011011111_101_1_110100110111;
      patterns[42750] = 29'b1_010011011111_110_1_010011011111;
      patterns[42751] = 29'b1_010011011111_111_1_010011011111;
      patterns[42752] = 29'b1_010011100000_000_1_010011100000;
      patterns[42753] = 29'b1_010011100000_001_1_100000010011;
      patterns[42754] = 29'b1_010011100000_010_0_100111000001;
      patterns[42755] = 29'b1_010011100000_011_1_001110000010;
      patterns[42756] = 29'b1_010011100000_100_0_101001110000;
      patterns[42757] = 29'b1_010011100000_101_0_010100111000;
      patterns[42758] = 29'b1_010011100000_110_1_010011100000;
      patterns[42759] = 29'b1_010011100000_111_1_010011100000;
      patterns[42760] = 29'b1_010011100001_000_1_010011100001;
      patterns[42761] = 29'b1_010011100001_001_1_100001010011;
      patterns[42762] = 29'b1_010011100001_010_0_100111000011;
      patterns[42763] = 29'b1_010011100001_011_1_001110000110;
      patterns[42764] = 29'b1_010011100001_100_1_101001110000;
      patterns[42765] = 29'b1_010011100001_101_0_110100111000;
      patterns[42766] = 29'b1_010011100001_110_1_010011100001;
      patterns[42767] = 29'b1_010011100001_111_1_010011100001;
      patterns[42768] = 29'b1_010011100010_000_1_010011100010;
      patterns[42769] = 29'b1_010011100010_001_1_100010010011;
      patterns[42770] = 29'b1_010011100010_010_0_100111000101;
      patterns[42771] = 29'b1_010011100010_011_1_001110001010;
      patterns[42772] = 29'b1_010011100010_100_0_101001110001;
      patterns[42773] = 29'b1_010011100010_101_1_010100111000;
      patterns[42774] = 29'b1_010011100010_110_1_010011100010;
      patterns[42775] = 29'b1_010011100010_111_1_010011100010;
      patterns[42776] = 29'b1_010011100011_000_1_010011100011;
      patterns[42777] = 29'b1_010011100011_001_1_100011010011;
      patterns[42778] = 29'b1_010011100011_010_0_100111000111;
      patterns[42779] = 29'b1_010011100011_011_1_001110001110;
      patterns[42780] = 29'b1_010011100011_100_1_101001110001;
      patterns[42781] = 29'b1_010011100011_101_1_110100111000;
      patterns[42782] = 29'b1_010011100011_110_1_010011100011;
      patterns[42783] = 29'b1_010011100011_111_1_010011100011;
      patterns[42784] = 29'b1_010011100100_000_1_010011100100;
      patterns[42785] = 29'b1_010011100100_001_1_100100010011;
      patterns[42786] = 29'b1_010011100100_010_0_100111001001;
      patterns[42787] = 29'b1_010011100100_011_1_001110010010;
      patterns[42788] = 29'b1_010011100100_100_0_101001110010;
      patterns[42789] = 29'b1_010011100100_101_0_010100111001;
      patterns[42790] = 29'b1_010011100100_110_1_010011100100;
      patterns[42791] = 29'b1_010011100100_111_1_010011100100;
      patterns[42792] = 29'b1_010011100101_000_1_010011100101;
      patterns[42793] = 29'b1_010011100101_001_1_100101010011;
      patterns[42794] = 29'b1_010011100101_010_0_100111001011;
      patterns[42795] = 29'b1_010011100101_011_1_001110010110;
      patterns[42796] = 29'b1_010011100101_100_1_101001110010;
      patterns[42797] = 29'b1_010011100101_101_0_110100111001;
      patterns[42798] = 29'b1_010011100101_110_1_010011100101;
      patterns[42799] = 29'b1_010011100101_111_1_010011100101;
      patterns[42800] = 29'b1_010011100110_000_1_010011100110;
      patterns[42801] = 29'b1_010011100110_001_1_100110010011;
      patterns[42802] = 29'b1_010011100110_010_0_100111001101;
      patterns[42803] = 29'b1_010011100110_011_1_001110011010;
      patterns[42804] = 29'b1_010011100110_100_0_101001110011;
      patterns[42805] = 29'b1_010011100110_101_1_010100111001;
      patterns[42806] = 29'b1_010011100110_110_1_010011100110;
      patterns[42807] = 29'b1_010011100110_111_1_010011100110;
      patterns[42808] = 29'b1_010011100111_000_1_010011100111;
      patterns[42809] = 29'b1_010011100111_001_1_100111010011;
      patterns[42810] = 29'b1_010011100111_010_0_100111001111;
      patterns[42811] = 29'b1_010011100111_011_1_001110011110;
      patterns[42812] = 29'b1_010011100111_100_1_101001110011;
      patterns[42813] = 29'b1_010011100111_101_1_110100111001;
      patterns[42814] = 29'b1_010011100111_110_1_010011100111;
      patterns[42815] = 29'b1_010011100111_111_1_010011100111;
      patterns[42816] = 29'b1_010011101000_000_1_010011101000;
      patterns[42817] = 29'b1_010011101000_001_1_101000010011;
      patterns[42818] = 29'b1_010011101000_010_0_100111010001;
      patterns[42819] = 29'b1_010011101000_011_1_001110100010;
      patterns[42820] = 29'b1_010011101000_100_0_101001110100;
      patterns[42821] = 29'b1_010011101000_101_0_010100111010;
      patterns[42822] = 29'b1_010011101000_110_1_010011101000;
      patterns[42823] = 29'b1_010011101000_111_1_010011101000;
      patterns[42824] = 29'b1_010011101001_000_1_010011101001;
      patterns[42825] = 29'b1_010011101001_001_1_101001010011;
      patterns[42826] = 29'b1_010011101001_010_0_100111010011;
      patterns[42827] = 29'b1_010011101001_011_1_001110100110;
      patterns[42828] = 29'b1_010011101001_100_1_101001110100;
      patterns[42829] = 29'b1_010011101001_101_0_110100111010;
      patterns[42830] = 29'b1_010011101001_110_1_010011101001;
      patterns[42831] = 29'b1_010011101001_111_1_010011101001;
      patterns[42832] = 29'b1_010011101010_000_1_010011101010;
      patterns[42833] = 29'b1_010011101010_001_1_101010010011;
      patterns[42834] = 29'b1_010011101010_010_0_100111010101;
      patterns[42835] = 29'b1_010011101010_011_1_001110101010;
      patterns[42836] = 29'b1_010011101010_100_0_101001110101;
      patterns[42837] = 29'b1_010011101010_101_1_010100111010;
      patterns[42838] = 29'b1_010011101010_110_1_010011101010;
      patterns[42839] = 29'b1_010011101010_111_1_010011101010;
      patterns[42840] = 29'b1_010011101011_000_1_010011101011;
      patterns[42841] = 29'b1_010011101011_001_1_101011010011;
      patterns[42842] = 29'b1_010011101011_010_0_100111010111;
      patterns[42843] = 29'b1_010011101011_011_1_001110101110;
      patterns[42844] = 29'b1_010011101011_100_1_101001110101;
      patterns[42845] = 29'b1_010011101011_101_1_110100111010;
      patterns[42846] = 29'b1_010011101011_110_1_010011101011;
      patterns[42847] = 29'b1_010011101011_111_1_010011101011;
      patterns[42848] = 29'b1_010011101100_000_1_010011101100;
      patterns[42849] = 29'b1_010011101100_001_1_101100010011;
      patterns[42850] = 29'b1_010011101100_010_0_100111011001;
      patterns[42851] = 29'b1_010011101100_011_1_001110110010;
      patterns[42852] = 29'b1_010011101100_100_0_101001110110;
      patterns[42853] = 29'b1_010011101100_101_0_010100111011;
      patterns[42854] = 29'b1_010011101100_110_1_010011101100;
      patterns[42855] = 29'b1_010011101100_111_1_010011101100;
      patterns[42856] = 29'b1_010011101101_000_1_010011101101;
      patterns[42857] = 29'b1_010011101101_001_1_101101010011;
      patterns[42858] = 29'b1_010011101101_010_0_100111011011;
      patterns[42859] = 29'b1_010011101101_011_1_001110110110;
      patterns[42860] = 29'b1_010011101101_100_1_101001110110;
      patterns[42861] = 29'b1_010011101101_101_0_110100111011;
      patterns[42862] = 29'b1_010011101101_110_1_010011101101;
      patterns[42863] = 29'b1_010011101101_111_1_010011101101;
      patterns[42864] = 29'b1_010011101110_000_1_010011101110;
      patterns[42865] = 29'b1_010011101110_001_1_101110010011;
      patterns[42866] = 29'b1_010011101110_010_0_100111011101;
      patterns[42867] = 29'b1_010011101110_011_1_001110111010;
      patterns[42868] = 29'b1_010011101110_100_0_101001110111;
      patterns[42869] = 29'b1_010011101110_101_1_010100111011;
      patterns[42870] = 29'b1_010011101110_110_1_010011101110;
      patterns[42871] = 29'b1_010011101110_111_1_010011101110;
      patterns[42872] = 29'b1_010011101111_000_1_010011101111;
      patterns[42873] = 29'b1_010011101111_001_1_101111010011;
      patterns[42874] = 29'b1_010011101111_010_0_100111011111;
      patterns[42875] = 29'b1_010011101111_011_1_001110111110;
      patterns[42876] = 29'b1_010011101111_100_1_101001110111;
      patterns[42877] = 29'b1_010011101111_101_1_110100111011;
      patterns[42878] = 29'b1_010011101111_110_1_010011101111;
      patterns[42879] = 29'b1_010011101111_111_1_010011101111;
      patterns[42880] = 29'b1_010011110000_000_1_010011110000;
      patterns[42881] = 29'b1_010011110000_001_1_110000010011;
      patterns[42882] = 29'b1_010011110000_010_0_100111100001;
      patterns[42883] = 29'b1_010011110000_011_1_001111000010;
      patterns[42884] = 29'b1_010011110000_100_0_101001111000;
      patterns[42885] = 29'b1_010011110000_101_0_010100111100;
      patterns[42886] = 29'b1_010011110000_110_1_010011110000;
      patterns[42887] = 29'b1_010011110000_111_1_010011110000;
      patterns[42888] = 29'b1_010011110001_000_1_010011110001;
      patterns[42889] = 29'b1_010011110001_001_1_110001010011;
      patterns[42890] = 29'b1_010011110001_010_0_100111100011;
      patterns[42891] = 29'b1_010011110001_011_1_001111000110;
      patterns[42892] = 29'b1_010011110001_100_1_101001111000;
      patterns[42893] = 29'b1_010011110001_101_0_110100111100;
      patterns[42894] = 29'b1_010011110001_110_1_010011110001;
      patterns[42895] = 29'b1_010011110001_111_1_010011110001;
      patterns[42896] = 29'b1_010011110010_000_1_010011110010;
      patterns[42897] = 29'b1_010011110010_001_1_110010010011;
      patterns[42898] = 29'b1_010011110010_010_0_100111100101;
      patterns[42899] = 29'b1_010011110010_011_1_001111001010;
      patterns[42900] = 29'b1_010011110010_100_0_101001111001;
      patterns[42901] = 29'b1_010011110010_101_1_010100111100;
      patterns[42902] = 29'b1_010011110010_110_1_010011110010;
      patterns[42903] = 29'b1_010011110010_111_1_010011110010;
      patterns[42904] = 29'b1_010011110011_000_1_010011110011;
      patterns[42905] = 29'b1_010011110011_001_1_110011010011;
      patterns[42906] = 29'b1_010011110011_010_0_100111100111;
      patterns[42907] = 29'b1_010011110011_011_1_001111001110;
      patterns[42908] = 29'b1_010011110011_100_1_101001111001;
      patterns[42909] = 29'b1_010011110011_101_1_110100111100;
      patterns[42910] = 29'b1_010011110011_110_1_010011110011;
      patterns[42911] = 29'b1_010011110011_111_1_010011110011;
      patterns[42912] = 29'b1_010011110100_000_1_010011110100;
      patterns[42913] = 29'b1_010011110100_001_1_110100010011;
      patterns[42914] = 29'b1_010011110100_010_0_100111101001;
      patterns[42915] = 29'b1_010011110100_011_1_001111010010;
      patterns[42916] = 29'b1_010011110100_100_0_101001111010;
      patterns[42917] = 29'b1_010011110100_101_0_010100111101;
      patterns[42918] = 29'b1_010011110100_110_1_010011110100;
      patterns[42919] = 29'b1_010011110100_111_1_010011110100;
      patterns[42920] = 29'b1_010011110101_000_1_010011110101;
      patterns[42921] = 29'b1_010011110101_001_1_110101010011;
      patterns[42922] = 29'b1_010011110101_010_0_100111101011;
      patterns[42923] = 29'b1_010011110101_011_1_001111010110;
      patterns[42924] = 29'b1_010011110101_100_1_101001111010;
      patterns[42925] = 29'b1_010011110101_101_0_110100111101;
      patterns[42926] = 29'b1_010011110101_110_1_010011110101;
      patterns[42927] = 29'b1_010011110101_111_1_010011110101;
      patterns[42928] = 29'b1_010011110110_000_1_010011110110;
      patterns[42929] = 29'b1_010011110110_001_1_110110010011;
      patterns[42930] = 29'b1_010011110110_010_0_100111101101;
      patterns[42931] = 29'b1_010011110110_011_1_001111011010;
      patterns[42932] = 29'b1_010011110110_100_0_101001111011;
      patterns[42933] = 29'b1_010011110110_101_1_010100111101;
      patterns[42934] = 29'b1_010011110110_110_1_010011110110;
      patterns[42935] = 29'b1_010011110110_111_1_010011110110;
      patterns[42936] = 29'b1_010011110111_000_1_010011110111;
      patterns[42937] = 29'b1_010011110111_001_1_110111010011;
      patterns[42938] = 29'b1_010011110111_010_0_100111101111;
      patterns[42939] = 29'b1_010011110111_011_1_001111011110;
      patterns[42940] = 29'b1_010011110111_100_1_101001111011;
      patterns[42941] = 29'b1_010011110111_101_1_110100111101;
      patterns[42942] = 29'b1_010011110111_110_1_010011110111;
      patterns[42943] = 29'b1_010011110111_111_1_010011110111;
      patterns[42944] = 29'b1_010011111000_000_1_010011111000;
      patterns[42945] = 29'b1_010011111000_001_1_111000010011;
      patterns[42946] = 29'b1_010011111000_010_0_100111110001;
      patterns[42947] = 29'b1_010011111000_011_1_001111100010;
      patterns[42948] = 29'b1_010011111000_100_0_101001111100;
      patterns[42949] = 29'b1_010011111000_101_0_010100111110;
      patterns[42950] = 29'b1_010011111000_110_1_010011111000;
      patterns[42951] = 29'b1_010011111000_111_1_010011111000;
      patterns[42952] = 29'b1_010011111001_000_1_010011111001;
      patterns[42953] = 29'b1_010011111001_001_1_111001010011;
      patterns[42954] = 29'b1_010011111001_010_0_100111110011;
      patterns[42955] = 29'b1_010011111001_011_1_001111100110;
      patterns[42956] = 29'b1_010011111001_100_1_101001111100;
      patterns[42957] = 29'b1_010011111001_101_0_110100111110;
      patterns[42958] = 29'b1_010011111001_110_1_010011111001;
      patterns[42959] = 29'b1_010011111001_111_1_010011111001;
      patterns[42960] = 29'b1_010011111010_000_1_010011111010;
      patterns[42961] = 29'b1_010011111010_001_1_111010010011;
      patterns[42962] = 29'b1_010011111010_010_0_100111110101;
      patterns[42963] = 29'b1_010011111010_011_1_001111101010;
      patterns[42964] = 29'b1_010011111010_100_0_101001111101;
      patterns[42965] = 29'b1_010011111010_101_1_010100111110;
      patterns[42966] = 29'b1_010011111010_110_1_010011111010;
      patterns[42967] = 29'b1_010011111010_111_1_010011111010;
      patterns[42968] = 29'b1_010011111011_000_1_010011111011;
      patterns[42969] = 29'b1_010011111011_001_1_111011010011;
      patterns[42970] = 29'b1_010011111011_010_0_100111110111;
      patterns[42971] = 29'b1_010011111011_011_1_001111101110;
      patterns[42972] = 29'b1_010011111011_100_1_101001111101;
      patterns[42973] = 29'b1_010011111011_101_1_110100111110;
      patterns[42974] = 29'b1_010011111011_110_1_010011111011;
      patterns[42975] = 29'b1_010011111011_111_1_010011111011;
      patterns[42976] = 29'b1_010011111100_000_1_010011111100;
      patterns[42977] = 29'b1_010011111100_001_1_111100010011;
      patterns[42978] = 29'b1_010011111100_010_0_100111111001;
      patterns[42979] = 29'b1_010011111100_011_1_001111110010;
      patterns[42980] = 29'b1_010011111100_100_0_101001111110;
      patterns[42981] = 29'b1_010011111100_101_0_010100111111;
      patterns[42982] = 29'b1_010011111100_110_1_010011111100;
      patterns[42983] = 29'b1_010011111100_111_1_010011111100;
      patterns[42984] = 29'b1_010011111101_000_1_010011111101;
      patterns[42985] = 29'b1_010011111101_001_1_111101010011;
      patterns[42986] = 29'b1_010011111101_010_0_100111111011;
      patterns[42987] = 29'b1_010011111101_011_1_001111110110;
      patterns[42988] = 29'b1_010011111101_100_1_101001111110;
      patterns[42989] = 29'b1_010011111101_101_0_110100111111;
      patterns[42990] = 29'b1_010011111101_110_1_010011111101;
      patterns[42991] = 29'b1_010011111101_111_1_010011111101;
      patterns[42992] = 29'b1_010011111110_000_1_010011111110;
      patterns[42993] = 29'b1_010011111110_001_1_111110010011;
      patterns[42994] = 29'b1_010011111110_010_0_100111111101;
      patterns[42995] = 29'b1_010011111110_011_1_001111111010;
      patterns[42996] = 29'b1_010011111110_100_0_101001111111;
      patterns[42997] = 29'b1_010011111110_101_1_010100111111;
      patterns[42998] = 29'b1_010011111110_110_1_010011111110;
      patterns[42999] = 29'b1_010011111110_111_1_010011111110;
      patterns[43000] = 29'b1_010011111111_000_1_010011111111;
      patterns[43001] = 29'b1_010011111111_001_1_111111010011;
      patterns[43002] = 29'b1_010011111111_010_0_100111111111;
      patterns[43003] = 29'b1_010011111111_011_1_001111111110;
      patterns[43004] = 29'b1_010011111111_100_1_101001111111;
      patterns[43005] = 29'b1_010011111111_101_1_110100111111;
      patterns[43006] = 29'b1_010011111111_110_1_010011111111;
      patterns[43007] = 29'b1_010011111111_111_1_010011111111;
      patterns[43008] = 29'b1_010100000000_000_1_010100000000;
      patterns[43009] = 29'b1_010100000000_001_1_000000010100;
      patterns[43010] = 29'b1_010100000000_010_0_101000000001;
      patterns[43011] = 29'b1_010100000000_011_1_010000000010;
      patterns[43012] = 29'b1_010100000000_100_0_101010000000;
      patterns[43013] = 29'b1_010100000000_101_0_010101000000;
      patterns[43014] = 29'b1_010100000000_110_1_010100000000;
      patterns[43015] = 29'b1_010100000000_111_1_010100000000;
      patterns[43016] = 29'b1_010100000001_000_1_010100000001;
      patterns[43017] = 29'b1_010100000001_001_1_000001010100;
      patterns[43018] = 29'b1_010100000001_010_0_101000000011;
      patterns[43019] = 29'b1_010100000001_011_1_010000000110;
      patterns[43020] = 29'b1_010100000001_100_1_101010000000;
      patterns[43021] = 29'b1_010100000001_101_0_110101000000;
      patterns[43022] = 29'b1_010100000001_110_1_010100000001;
      patterns[43023] = 29'b1_010100000001_111_1_010100000001;
      patterns[43024] = 29'b1_010100000010_000_1_010100000010;
      patterns[43025] = 29'b1_010100000010_001_1_000010010100;
      patterns[43026] = 29'b1_010100000010_010_0_101000000101;
      patterns[43027] = 29'b1_010100000010_011_1_010000001010;
      patterns[43028] = 29'b1_010100000010_100_0_101010000001;
      patterns[43029] = 29'b1_010100000010_101_1_010101000000;
      patterns[43030] = 29'b1_010100000010_110_1_010100000010;
      patterns[43031] = 29'b1_010100000010_111_1_010100000010;
      patterns[43032] = 29'b1_010100000011_000_1_010100000011;
      patterns[43033] = 29'b1_010100000011_001_1_000011010100;
      patterns[43034] = 29'b1_010100000011_010_0_101000000111;
      patterns[43035] = 29'b1_010100000011_011_1_010000001110;
      patterns[43036] = 29'b1_010100000011_100_1_101010000001;
      patterns[43037] = 29'b1_010100000011_101_1_110101000000;
      patterns[43038] = 29'b1_010100000011_110_1_010100000011;
      patterns[43039] = 29'b1_010100000011_111_1_010100000011;
      patterns[43040] = 29'b1_010100000100_000_1_010100000100;
      patterns[43041] = 29'b1_010100000100_001_1_000100010100;
      patterns[43042] = 29'b1_010100000100_010_0_101000001001;
      patterns[43043] = 29'b1_010100000100_011_1_010000010010;
      patterns[43044] = 29'b1_010100000100_100_0_101010000010;
      patterns[43045] = 29'b1_010100000100_101_0_010101000001;
      patterns[43046] = 29'b1_010100000100_110_1_010100000100;
      patterns[43047] = 29'b1_010100000100_111_1_010100000100;
      patterns[43048] = 29'b1_010100000101_000_1_010100000101;
      patterns[43049] = 29'b1_010100000101_001_1_000101010100;
      patterns[43050] = 29'b1_010100000101_010_0_101000001011;
      patterns[43051] = 29'b1_010100000101_011_1_010000010110;
      patterns[43052] = 29'b1_010100000101_100_1_101010000010;
      patterns[43053] = 29'b1_010100000101_101_0_110101000001;
      patterns[43054] = 29'b1_010100000101_110_1_010100000101;
      patterns[43055] = 29'b1_010100000101_111_1_010100000101;
      patterns[43056] = 29'b1_010100000110_000_1_010100000110;
      patterns[43057] = 29'b1_010100000110_001_1_000110010100;
      patterns[43058] = 29'b1_010100000110_010_0_101000001101;
      patterns[43059] = 29'b1_010100000110_011_1_010000011010;
      patterns[43060] = 29'b1_010100000110_100_0_101010000011;
      patterns[43061] = 29'b1_010100000110_101_1_010101000001;
      patterns[43062] = 29'b1_010100000110_110_1_010100000110;
      patterns[43063] = 29'b1_010100000110_111_1_010100000110;
      patterns[43064] = 29'b1_010100000111_000_1_010100000111;
      patterns[43065] = 29'b1_010100000111_001_1_000111010100;
      patterns[43066] = 29'b1_010100000111_010_0_101000001111;
      patterns[43067] = 29'b1_010100000111_011_1_010000011110;
      patterns[43068] = 29'b1_010100000111_100_1_101010000011;
      patterns[43069] = 29'b1_010100000111_101_1_110101000001;
      patterns[43070] = 29'b1_010100000111_110_1_010100000111;
      patterns[43071] = 29'b1_010100000111_111_1_010100000111;
      patterns[43072] = 29'b1_010100001000_000_1_010100001000;
      patterns[43073] = 29'b1_010100001000_001_1_001000010100;
      patterns[43074] = 29'b1_010100001000_010_0_101000010001;
      patterns[43075] = 29'b1_010100001000_011_1_010000100010;
      patterns[43076] = 29'b1_010100001000_100_0_101010000100;
      patterns[43077] = 29'b1_010100001000_101_0_010101000010;
      patterns[43078] = 29'b1_010100001000_110_1_010100001000;
      patterns[43079] = 29'b1_010100001000_111_1_010100001000;
      patterns[43080] = 29'b1_010100001001_000_1_010100001001;
      patterns[43081] = 29'b1_010100001001_001_1_001001010100;
      patterns[43082] = 29'b1_010100001001_010_0_101000010011;
      patterns[43083] = 29'b1_010100001001_011_1_010000100110;
      patterns[43084] = 29'b1_010100001001_100_1_101010000100;
      patterns[43085] = 29'b1_010100001001_101_0_110101000010;
      patterns[43086] = 29'b1_010100001001_110_1_010100001001;
      patterns[43087] = 29'b1_010100001001_111_1_010100001001;
      patterns[43088] = 29'b1_010100001010_000_1_010100001010;
      patterns[43089] = 29'b1_010100001010_001_1_001010010100;
      patterns[43090] = 29'b1_010100001010_010_0_101000010101;
      patterns[43091] = 29'b1_010100001010_011_1_010000101010;
      patterns[43092] = 29'b1_010100001010_100_0_101010000101;
      patterns[43093] = 29'b1_010100001010_101_1_010101000010;
      patterns[43094] = 29'b1_010100001010_110_1_010100001010;
      patterns[43095] = 29'b1_010100001010_111_1_010100001010;
      patterns[43096] = 29'b1_010100001011_000_1_010100001011;
      patterns[43097] = 29'b1_010100001011_001_1_001011010100;
      patterns[43098] = 29'b1_010100001011_010_0_101000010111;
      patterns[43099] = 29'b1_010100001011_011_1_010000101110;
      patterns[43100] = 29'b1_010100001011_100_1_101010000101;
      patterns[43101] = 29'b1_010100001011_101_1_110101000010;
      patterns[43102] = 29'b1_010100001011_110_1_010100001011;
      patterns[43103] = 29'b1_010100001011_111_1_010100001011;
      patterns[43104] = 29'b1_010100001100_000_1_010100001100;
      patterns[43105] = 29'b1_010100001100_001_1_001100010100;
      patterns[43106] = 29'b1_010100001100_010_0_101000011001;
      patterns[43107] = 29'b1_010100001100_011_1_010000110010;
      patterns[43108] = 29'b1_010100001100_100_0_101010000110;
      patterns[43109] = 29'b1_010100001100_101_0_010101000011;
      patterns[43110] = 29'b1_010100001100_110_1_010100001100;
      patterns[43111] = 29'b1_010100001100_111_1_010100001100;
      patterns[43112] = 29'b1_010100001101_000_1_010100001101;
      patterns[43113] = 29'b1_010100001101_001_1_001101010100;
      patterns[43114] = 29'b1_010100001101_010_0_101000011011;
      patterns[43115] = 29'b1_010100001101_011_1_010000110110;
      patterns[43116] = 29'b1_010100001101_100_1_101010000110;
      patterns[43117] = 29'b1_010100001101_101_0_110101000011;
      patterns[43118] = 29'b1_010100001101_110_1_010100001101;
      patterns[43119] = 29'b1_010100001101_111_1_010100001101;
      patterns[43120] = 29'b1_010100001110_000_1_010100001110;
      patterns[43121] = 29'b1_010100001110_001_1_001110010100;
      patterns[43122] = 29'b1_010100001110_010_0_101000011101;
      patterns[43123] = 29'b1_010100001110_011_1_010000111010;
      patterns[43124] = 29'b1_010100001110_100_0_101010000111;
      patterns[43125] = 29'b1_010100001110_101_1_010101000011;
      patterns[43126] = 29'b1_010100001110_110_1_010100001110;
      patterns[43127] = 29'b1_010100001110_111_1_010100001110;
      patterns[43128] = 29'b1_010100001111_000_1_010100001111;
      patterns[43129] = 29'b1_010100001111_001_1_001111010100;
      patterns[43130] = 29'b1_010100001111_010_0_101000011111;
      patterns[43131] = 29'b1_010100001111_011_1_010000111110;
      patterns[43132] = 29'b1_010100001111_100_1_101010000111;
      patterns[43133] = 29'b1_010100001111_101_1_110101000011;
      patterns[43134] = 29'b1_010100001111_110_1_010100001111;
      patterns[43135] = 29'b1_010100001111_111_1_010100001111;
      patterns[43136] = 29'b1_010100010000_000_1_010100010000;
      patterns[43137] = 29'b1_010100010000_001_1_010000010100;
      patterns[43138] = 29'b1_010100010000_010_0_101000100001;
      patterns[43139] = 29'b1_010100010000_011_1_010001000010;
      patterns[43140] = 29'b1_010100010000_100_0_101010001000;
      patterns[43141] = 29'b1_010100010000_101_0_010101000100;
      patterns[43142] = 29'b1_010100010000_110_1_010100010000;
      patterns[43143] = 29'b1_010100010000_111_1_010100010000;
      patterns[43144] = 29'b1_010100010001_000_1_010100010001;
      patterns[43145] = 29'b1_010100010001_001_1_010001010100;
      patterns[43146] = 29'b1_010100010001_010_0_101000100011;
      patterns[43147] = 29'b1_010100010001_011_1_010001000110;
      patterns[43148] = 29'b1_010100010001_100_1_101010001000;
      patterns[43149] = 29'b1_010100010001_101_0_110101000100;
      patterns[43150] = 29'b1_010100010001_110_1_010100010001;
      patterns[43151] = 29'b1_010100010001_111_1_010100010001;
      patterns[43152] = 29'b1_010100010010_000_1_010100010010;
      patterns[43153] = 29'b1_010100010010_001_1_010010010100;
      patterns[43154] = 29'b1_010100010010_010_0_101000100101;
      patterns[43155] = 29'b1_010100010010_011_1_010001001010;
      patterns[43156] = 29'b1_010100010010_100_0_101010001001;
      patterns[43157] = 29'b1_010100010010_101_1_010101000100;
      patterns[43158] = 29'b1_010100010010_110_1_010100010010;
      patterns[43159] = 29'b1_010100010010_111_1_010100010010;
      patterns[43160] = 29'b1_010100010011_000_1_010100010011;
      patterns[43161] = 29'b1_010100010011_001_1_010011010100;
      patterns[43162] = 29'b1_010100010011_010_0_101000100111;
      patterns[43163] = 29'b1_010100010011_011_1_010001001110;
      patterns[43164] = 29'b1_010100010011_100_1_101010001001;
      patterns[43165] = 29'b1_010100010011_101_1_110101000100;
      patterns[43166] = 29'b1_010100010011_110_1_010100010011;
      patterns[43167] = 29'b1_010100010011_111_1_010100010011;
      patterns[43168] = 29'b1_010100010100_000_1_010100010100;
      patterns[43169] = 29'b1_010100010100_001_1_010100010100;
      patterns[43170] = 29'b1_010100010100_010_0_101000101001;
      patterns[43171] = 29'b1_010100010100_011_1_010001010010;
      patterns[43172] = 29'b1_010100010100_100_0_101010001010;
      patterns[43173] = 29'b1_010100010100_101_0_010101000101;
      patterns[43174] = 29'b1_010100010100_110_1_010100010100;
      patterns[43175] = 29'b1_010100010100_111_1_010100010100;
      patterns[43176] = 29'b1_010100010101_000_1_010100010101;
      patterns[43177] = 29'b1_010100010101_001_1_010101010100;
      patterns[43178] = 29'b1_010100010101_010_0_101000101011;
      patterns[43179] = 29'b1_010100010101_011_1_010001010110;
      patterns[43180] = 29'b1_010100010101_100_1_101010001010;
      patterns[43181] = 29'b1_010100010101_101_0_110101000101;
      patterns[43182] = 29'b1_010100010101_110_1_010100010101;
      patterns[43183] = 29'b1_010100010101_111_1_010100010101;
      patterns[43184] = 29'b1_010100010110_000_1_010100010110;
      patterns[43185] = 29'b1_010100010110_001_1_010110010100;
      patterns[43186] = 29'b1_010100010110_010_0_101000101101;
      patterns[43187] = 29'b1_010100010110_011_1_010001011010;
      patterns[43188] = 29'b1_010100010110_100_0_101010001011;
      patterns[43189] = 29'b1_010100010110_101_1_010101000101;
      patterns[43190] = 29'b1_010100010110_110_1_010100010110;
      patterns[43191] = 29'b1_010100010110_111_1_010100010110;
      patterns[43192] = 29'b1_010100010111_000_1_010100010111;
      patterns[43193] = 29'b1_010100010111_001_1_010111010100;
      patterns[43194] = 29'b1_010100010111_010_0_101000101111;
      patterns[43195] = 29'b1_010100010111_011_1_010001011110;
      patterns[43196] = 29'b1_010100010111_100_1_101010001011;
      patterns[43197] = 29'b1_010100010111_101_1_110101000101;
      patterns[43198] = 29'b1_010100010111_110_1_010100010111;
      patterns[43199] = 29'b1_010100010111_111_1_010100010111;
      patterns[43200] = 29'b1_010100011000_000_1_010100011000;
      patterns[43201] = 29'b1_010100011000_001_1_011000010100;
      patterns[43202] = 29'b1_010100011000_010_0_101000110001;
      patterns[43203] = 29'b1_010100011000_011_1_010001100010;
      patterns[43204] = 29'b1_010100011000_100_0_101010001100;
      patterns[43205] = 29'b1_010100011000_101_0_010101000110;
      patterns[43206] = 29'b1_010100011000_110_1_010100011000;
      patterns[43207] = 29'b1_010100011000_111_1_010100011000;
      patterns[43208] = 29'b1_010100011001_000_1_010100011001;
      patterns[43209] = 29'b1_010100011001_001_1_011001010100;
      patterns[43210] = 29'b1_010100011001_010_0_101000110011;
      patterns[43211] = 29'b1_010100011001_011_1_010001100110;
      patterns[43212] = 29'b1_010100011001_100_1_101010001100;
      patterns[43213] = 29'b1_010100011001_101_0_110101000110;
      patterns[43214] = 29'b1_010100011001_110_1_010100011001;
      patterns[43215] = 29'b1_010100011001_111_1_010100011001;
      patterns[43216] = 29'b1_010100011010_000_1_010100011010;
      patterns[43217] = 29'b1_010100011010_001_1_011010010100;
      patterns[43218] = 29'b1_010100011010_010_0_101000110101;
      patterns[43219] = 29'b1_010100011010_011_1_010001101010;
      patterns[43220] = 29'b1_010100011010_100_0_101010001101;
      patterns[43221] = 29'b1_010100011010_101_1_010101000110;
      patterns[43222] = 29'b1_010100011010_110_1_010100011010;
      patterns[43223] = 29'b1_010100011010_111_1_010100011010;
      patterns[43224] = 29'b1_010100011011_000_1_010100011011;
      patterns[43225] = 29'b1_010100011011_001_1_011011010100;
      patterns[43226] = 29'b1_010100011011_010_0_101000110111;
      patterns[43227] = 29'b1_010100011011_011_1_010001101110;
      patterns[43228] = 29'b1_010100011011_100_1_101010001101;
      patterns[43229] = 29'b1_010100011011_101_1_110101000110;
      patterns[43230] = 29'b1_010100011011_110_1_010100011011;
      patterns[43231] = 29'b1_010100011011_111_1_010100011011;
      patterns[43232] = 29'b1_010100011100_000_1_010100011100;
      patterns[43233] = 29'b1_010100011100_001_1_011100010100;
      patterns[43234] = 29'b1_010100011100_010_0_101000111001;
      patterns[43235] = 29'b1_010100011100_011_1_010001110010;
      patterns[43236] = 29'b1_010100011100_100_0_101010001110;
      patterns[43237] = 29'b1_010100011100_101_0_010101000111;
      patterns[43238] = 29'b1_010100011100_110_1_010100011100;
      patterns[43239] = 29'b1_010100011100_111_1_010100011100;
      patterns[43240] = 29'b1_010100011101_000_1_010100011101;
      patterns[43241] = 29'b1_010100011101_001_1_011101010100;
      patterns[43242] = 29'b1_010100011101_010_0_101000111011;
      patterns[43243] = 29'b1_010100011101_011_1_010001110110;
      patterns[43244] = 29'b1_010100011101_100_1_101010001110;
      patterns[43245] = 29'b1_010100011101_101_0_110101000111;
      patterns[43246] = 29'b1_010100011101_110_1_010100011101;
      patterns[43247] = 29'b1_010100011101_111_1_010100011101;
      patterns[43248] = 29'b1_010100011110_000_1_010100011110;
      patterns[43249] = 29'b1_010100011110_001_1_011110010100;
      patterns[43250] = 29'b1_010100011110_010_0_101000111101;
      patterns[43251] = 29'b1_010100011110_011_1_010001111010;
      patterns[43252] = 29'b1_010100011110_100_0_101010001111;
      patterns[43253] = 29'b1_010100011110_101_1_010101000111;
      patterns[43254] = 29'b1_010100011110_110_1_010100011110;
      patterns[43255] = 29'b1_010100011110_111_1_010100011110;
      patterns[43256] = 29'b1_010100011111_000_1_010100011111;
      patterns[43257] = 29'b1_010100011111_001_1_011111010100;
      patterns[43258] = 29'b1_010100011111_010_0_101000111111;
      patterns[43259] = 29'b1_010100011111_011_1_010001111110;
      patterns[43260] = 29'b1_010100011111_100_1_101010001111;
      patterns[43261] = 29'b1_010100011111_101_1_110101000111;
      patterns[43262] = 29'b1_010100011111_110_1_010100011111;
      patterns[43263] = 29'b1_010100011111_111_1_010100011111;
      patterns[43264] = 29'b1_010100100000_000_1_010100100000;
      patterns[43265] = 29'b1_010100100000_001_1_100000010100;
      patterns[43266] = 29'b1_010100100000_010_0_101001000001;
      patterns[43267] = 29'b1_010100100000_011_1_010010000010;
      patterns[43268] = 29'b1_010100100000_100_0_101010010000;
      patterns[43269] = 29'b1_010100100000_101_0_010101001000;
      patterns[43270] = 29'b1_010100100000_110_1_010100100000;
      patterns[43271] = 29'b1_010100100000_111_1_010100100000;
      patterns[43272] = 29'b1_010100100001_000_1_010100100001;
      patterns[43273] = 29'b1_010100100001_001_1_100001010100;
      patterns[43274] = 29'b1_010100100001_010_0_101001000011;
      patterns[43275] = 29'b1_010100100001_011_1_010010000110;
      patterns[43276] = 29'b1_010100100001_100_1_101010010000;
      patterns[43277] = 29'b1_010100100001_101_0_110101001000;
      patterns[43278] = 29'b1_010100100001_110_1_010100100001;
      patterns[43279] = 29'b1_010100100001_111_1_010100100001;
      patterns[43280] = 29'b1_010100100010_000_1_010100100010;
      patterns[43281] = 29'b1_010100100010_001_1_100010010100;
      patterns[43282] = 29'b1_010100100010_010_0_101001000101;
      patterns[43283] = 29'b1_010100100010_011_1_010010001010;
      patterns[43284] = 29'b1_010100100010_100_0_101010010001;
      patterns[43285] = 29'b1_010100100010_101_1_010101001000;
      patterns[43286] = 29'b1_010100100010_110_1_010100100010;
      patterns[43287] = 29'b1_010100100010_111_1_010100100010;
      patterns[43288] = 29'b1_010100100011_000_1_010100100011;
      patterns[43289] = 29'b1_010100100011_001_1_100011010100;
      patterns[43290] = 29'b1_010100100011_010_0_101001000111;
      patterns[43291] = 29'b1_010100100011_011_1_010010001110;
      patterns[43292] = 29'b1_010100100011_100_1_101010010001;
      patterns[43293] = 29'b1_010100100011_101_1_110101001000;
      patterns[43294] = 29'b1_010100100011_110_1_010100100011;
      patterns[43295] = 29'b1_010100100011_111_1_010100100011;
      patterns[43296] = 29'b1_010100100100_000_1_010100100100;
      patterns[43297] = 29'b1_010100100100_001_1_100100010100;
      patterns[43298] = 29'b1_010100100100_010_0_101001001001;
      patterns[43299] = 29'b1_010100100100_011_1_010010010010;
      patterns[43300] = 29'b1_010100100100_100_0_101010010010;
      patterns[43301] = 29'b1_010100100100_101_0_010101001001;
      patterns[43302] = 29'b1_010100100100_110_1_010100100100;
      patterns[43303] = 29'b1_010100100100_111_1_010100100100;
      patterns[43304] = 29'b1_010100100101_000_1_010100100101;
      patterns[43305] = 29'b1_010100100101_001_1_100101010100;
      patterns[43306] = 29'b1_010100100101_010_0_101001001011;
      patterns[43307] = 29'b1_010100100101_011_1_010010010110;
      patterns[43308] = 29'b1_010100100101_100_1_101010010010;
      patterns[43309] = 29'b1_010100100101_101_0_110101001001;
      patterns[43310] = 29'b1_010100100101_110_1_010100100101;
      patterns[43311] = 29'b1_010100100101_111_1_010100100101;
      patterns[43312] = 29'b1_010100100110_000_1_010100100110;
      patterns[43313] = 29'b1_010100100110_001_1_100110010100;
      patterns[43314] = 29'b1_010100100110_010_0_101001001101;
      patterns[43315] = 29'b1_010100100110_011_1_010010011010;
      patterns[43316] = 29'b1_010100100110_100_0_101010010011;
      patterns[43317] = 29'b1_010100100110_101_1_010101001001;
      patterns[43318] = 29'b1_010100100110_110_1_010100100110;
      patterns[43319] = 29'b1_010100100110_111_1_010100100110;
      patterns[43320] = 29'b1_010100100111_000_1_010100100111;
      patterns[43321] = 29'b1_010100100111_001_1_100111010100;
      patterns[43322] = 29'b1_010100100111_010_0_101001001111;
      patterns[43323] = 29'b1_010100100111_011_1_010010011110;
      patterns[43324] = 29'b1_010100100111_100_1_101010010011;
      patterns[43325] = 29'b1_010100100111_101_1_110101001001;
      patterns[43326] = 29'b1_010100100111_110_1_010100100111;
      patterns[43327] = 29'b1_010100100111_111_1_010100100111;
      patterns[43328] = 29'b1_010100101000_000_1_010100101000;
      patterns[43329] = 29'b1_010100101000_001_1_101000010100;
      patterns[43330] = 29'b1_010100101000_010_0_101001010001;
      patterns[43331] = 29'b1_010100101000_011_1_010010100010;
      patterns[43332] = 29'b1_010100101000_100_0_101010010100;
      patterns[43333] = 29'b1_010100101000_101_0_010101001010;
      patterns[43334] = 29'b1_010100101000_110_1_010100101000;
      patterns[43335] = 29'b1_010100101000_111_1_010100101000;
      patterns[43336] = 29'b1_010100101001_000_1_010100101001;
      patterns[43337] = 29'b1_010100101001_001_1_101001010100;
      patterns[43338] = 29'b1_010100101001_010_0_101001010011;
      patterns[43339] = 29'b1_010100101001_011_1_010010100110;
      patterns[43340] = 29'b1_010100101001_100_1_101010010100;
      patterns[43341] = 29'b1_010100101001_101_0_110101001010;
      patterns[43342] = 29'b1_010100101001_110_1_010100101001;
      patterns[43343] = 29'b1_010100101001_111_1_010100101001;
      patterns[43344] = 29'b1_010100101010_000_1_010100101010;
      patterns[43345] = 29'b1_010100101010_001_1_101010010100;
      patterns[43346] = 29'b1_010100101010_010_0_101001010101;
      patterns[43347] = 29'b1_010100101010_011_1_010010101010;
      patterns[43348] = 29'b1_010100101010_100_0_101010010101;
      patterns[43349] = 29'b1_010100101010_101_1_010101001010;
      patterns[43350] = 29'b1_010100101010_110_1_010100101010;
      patterns[43351] = 29'b1_010100101010_111_1_010100101010;
      patterns[43352] = 29'b1_010100101011_000_1_010100101011;
      patterns[43353] = 29'b1_010100101011_001_1_101011010100;
      patterns[43354] = 29'b1_010100101011_010_0_101001010111;
      patterns[43355] = 29'b1_010100101011_011_1_010010101110;
      patterns[43356] = 29'b1_010100101011_100_1_101010010101;
      patterns[43357] = 29'b1_010100101011_101_1_110101001010;
      patterns[43358] = 29'b1_010100101011_110_1_010100101011;
      patterns[43359] = 29'b1_010100101011_111_1_010100101011;
      patterns[43360] = 29'b1_010100101100_000_1_010100101100;
      patterns[43361] = 29'b1_010100101100_001_1_101100010100;
      patterns[43362] = 29'b1_010100101100_010_0_101001011001;
      patterns[43363] = 29'b1_010100101100_011_1_010010110010;
      patterns[43364] = 29'b1_010100101100_100_0_101010010110;
      patterns[43365] = 29'b1_010100101100_101_0_010101001011;
      patterns[43366] = 29'b1_010100101100_110_1_010100101100;
      patterns[43367] = 29'b1_010100101100_111_1_010100101100;
      patterns[43368] = 29'b1_010100101101_000_1_010100101101;
      patterns[43369] = 29'b1_010100101101_001_1_101101010100;
      patterns[43370] = 29'b1_010100101101_010_0_101001011011;
      patterns[43371] = 29'b1_010100101101_011_1_010010110110;
      patterns[43372] = 29'b1_010100101101_100_1_101010010110;
      patterns[43373] = 29'b1_010100101101_101_0_110101001011;
      patterns[43374] = 29'b1_010100101101_110_1_010100101101;
      patterns[43375] = 29'b1_010100101101_111_1_010100101101;
      patterns[43376] = 29'b1_010100101110_000_1_010100101110;
      patterns[43377] = 29'b1_010100101110_001_1_101110010100;
      patterns[43378] = 29'b1_010100101110_010_0_101001011101;
      patterns[43379] = 29'b1_010100101110_011_1_010010111010;
      patterns[43380] = 29'b1_010100101110_100_0_101010010111;
      patterns[43381] = 29'b1_010100101110_101_1_010101001011;
      patterns[43382] = 29'b1_010100101110_110_1_010100101110;
      patterns[43383] = 29'b1_010100101110_111_1_010100101110;
      patterns[43384] = 29'b1_010100101111_000_1_010100101111;
      patterns[43385] = 29'b1_010100101111_001_1_101111010100;
      patterns[43386] = 29'b1_010100101111_010_0_101001011111;
      patterns[43387] = 29'b1_010100101111_011_1_010010111110;
      patterns[43388] = 29'b1_010100101111_100_1_101010010111;
      patterns[43389] = 29'b1_010100101111_101_1_110101001011;
      patterns[43390] = 29'b1_010100101111_110_1_010100101111;
      patterns[43391] = 29'b1_010100101111_111_1_010100101111;
      patterns[43392] = 29'b1_010100110000_000_1_010100110000;
      patterns[43393] = 29'b1_010100110000_001_1_110000010100;
      patterns[43394] = 29'b1_010100110000_010_0_101001100001;
      patterns[43395] = 29'b1_010100110000_011_1_010011000010;
      patterns[43396] = 29'b1_010100110000_100_0_101010011000;
      patterns[43397] = 29'b1_010100110000_101_0_010101001100;
      patterns[43398] = 29'b1_010100110000_110_1_010100110000;
      patterns[43399] = 29'b1_010100110000_111_1_010100110000;
      patterns[43400] = 29'b1_010100110001_000_1_010100110001;
      patterns[43401] = 29'b1_010100110001_001_1_110001010100;
      patterns[43402] = 29'b1_010100110001_010_0_101001100011;
      patterns[43403] = 29'b1_010100110001_011_1_010011000110;
      patterns[43404] = 29'b1_010100110001_100_1_101010011000;
      patterns[43405] = 29'b1_010100110001_101_0_110101001100;
      patterns[43406] = 29'b1_010100110001_110_1_010100110001;
      patterns[43407] = 29'b1_010100110001_111_1_010100110001;
      patterns[43408] = 29'b1_010100110010_000_1_010100110010;
      patterns[43409] = 29'b1_010100110010_001_1_110010010100;
      patterns[43410] = 29'b1_010100110010_010_0_101001100101;
      patterns[43411] = 29'b1_010100110010_011_1_010011001010;
      patterns[43412] = 29'b1_010100110010_100_0_101010011001;
      patterns[43413] = 29'b1_010100110010_101_1_010101001100;
      patterns[43414] = 29'b1_010100110010_110_1_010100110010;
      patterns[43415] = 29'b1_010100110010_111_1_010100110010;
      patterns[43416] = 29'b1_010100110011_000_1_010100110011;
      patterns[43417] = 29'b1_010100110011_001_1_110011010100;
      patterns[43418] = 29'b1_010100110011_010_0_101001100111;
      patterns[43419] = 29'b1_010100110011_011_1_010011001110;
      patterns[43420] = 29'b1_010100110011_100_1_101010011001;
      patterns[43421] = 29'b1_010100110011_101_1_110101001100;
      patterns[43422] = 29'b1_010100110011_110_1_010100110011;
      patterns[43423] = 29'b1_010100110011_111_1_010100110011;
      patterns[43424] = 29'b1_010100110100_000_1_010100110100;
      patterns[43425] = 29'b1_010100110100_001_1_110100010100;
      patterns[43426] = 29'b1_010100110100_010_0_101001101001;
      patterns[43427] = 29'b1_010100110100_011_1_010011010010;
      patterns[43428] = 29'b1_010100110100_100_0_101010011010;
      patterns[43429] = 29'b1_010100110100_101_0_010101001101;
      patterns[43430] = 29'b1_010100110100_110_1_010100110100;
      patterns[43431] = 29'b1_010100110100_111_1_010100110100;
      patterns[43432] = 29'b1_010100110101_000_1_010100110101;
      patterns[43433] = 29'b1_010100110101_001_1_110101010100;
      patterns[43434] = 29'b1_010100110101_010_0_101001101011;
      patterns[43435] = 29'b1_010100110101_011_1_010011010110;
      patterns[43436] = 29'b1_010100110101_100_1_101010011010;
      patterns[43437] = 29'b1_010100110101_101_0_110101001101;
      patterns[43438] = 29'b1_010100110101_110_1_010100110101;
      patterns[43439] = 29'b1_010100110101_111_1_010100110101;
      patterns[43440] = 29'b1_010100110110_000_1_010100110110;
      patterns[43441] = 29'b1_010100110110_001_1_110110010100;
      patterns[43442] = 29'b1_010100110110_010_0_101001101101;
      patterns[43443] = 29'b1_010100110110_011_1_010011011010;
      patterns[43444] = 29'b1_010100110110_100_0_101010011011;
      patterns[43445] = 29'b1_010100110110_101_1_010101001101;
      patterns[43446] = 29'b1_010100110110_110_1_010100110110;
      patterns[43447] = 29'b1_010100110110_111_1_010100110110;
      patterns[43448] = 29'b1_010100110111_000_1_010100110111;
      patterns[43449] = 29'b1_010100110111_001_1_110111010100;
      patterns[43450] = 29'b1_010100110111_010_0_101001101111;
      patterns[43451] = 29'b1_010100110111_011_1_010011011110;
      patterns[43452] = 29'b1_010100110111_100_1_101010011011;
      patterns[43453] = 29'b1_010100110111_101_1_110101001101;
      patterns[43454] = 29'b1_010100110111_110_1_010100110111;
      patterns[43455] = 29'b1_010100110111_111_1_010100110111;
      patterns[43456] = 29'b1_010100111000_000_1_010100111000;
      patterns[43457] = 29'b1_010100111000_001_1_111000010100;
      patterns[43458] = 29'b1_010100111000_010_0_101001110001;
      patterns[43459] = 29'b1_010100111000_011_1_010011100010;
      patterns[43460] = 29'b1_010100111000_100_0_101010011100;
      patterns[43461] = 29'b1_010100111000_101_0_010101001110;
      patterns[43462] = 29'b1_010100111000_110_1_010100111000;
      patterns[43463] = 29'b1_010100111000_111_1_010100111000;
      patterns[43464] = 29'b1_010100111001_000_1_010100111001;
      patterns[43465] = 29'b1_010100111001_001_1_111001010100;
      patterns[43466] = 29'b1_010100111001_010_0_101001110011;
      patterns[43467] = 29'b1_010100111001_011_1_010011100110;
      patterns[43468] = 29'b1_010100111001_100_1_101010011100;
      patterns[43469] = 29'b1_010100111001_101_0_110101001110;
      patterns[43470] = 29'b1_010100111001_110_1_010100111001;
      patterns[43471] = 29'b1_010100111001_111_1_010100111001;
      patterns[43472] = 29'b1_010100111010_000_1_010100111010;
      patterns[43473] = 29'b1_010100111010_001_1_111010010100;
      patterns[43474] = 29'b1_010100111010_010_0_101001110101;
      patterns[43475] = 29'b1_010100111010_011_1_010011101010;
      patterns[43476] = 29'b1_010100111010_100_0_101010011101;
      patterns[43477] = 29'b1_010100111010_101_1_010101001110;
      patterns[43478] = 29'b1_010100111010_110_1_010100111010;
      patterns[43479] = 29'b1_010100111010_111_1_010100111010;
      patterns[43480] = 29'b1_010100111011_000_1_010100111011;
      patterns[43481] = 29'b1_010100111011_001_1_111011010100;
      patterns[43482] = 29'b1_010100111011_010_0_101001110111;
      patterns[43483] = 29'b1_010100111011_011_1_010011101110;
      patterns[43484] = 29'b1_010100111011_100_1_101010011101;
      patterns[43485] = 29'b1_010100111011_101_1_110101001110;
      patterns[43486] = 29'b1_010100111011_110_1_010100111011;
      patterns[43487] = 29'b1_010100111011_111_1_010100111011;
      patterns[43488] = 29'b1_010100111100_000_1_010100111100;
      patterns[43489] = 29'b1_010100111100_001_1_111100010100;
      patterns[43490] = 29'b1_010100111100_010_0_101001111001;
      patterns[43491] = 29'b1_010100111100_011_1_010011110010;
      patterns[43492] = 29'b1_010100111100_100_0_101010011110;
      patterns[43493] = 29'b1_010100111100_101_0_010101001111;
      patterns[43494] = 29'b1_010100111100_110_1_010100111100;
      patterns[43495] = 29'b1_010100111100_111_1_010100111100;
      patterns[43496] = 29'b1_010100111101_000_1_010100111101;
      patterns[43497] = 29'b1_010100111101_001_1_111101010100;
      patterns[43498] = 29'b1_010100111101_010_0_101001111011;
      patterns[43499] = 29'b1_010100111101_011_1_010011110110;
      patterns[43500] = 29'b1_010100111101_100_1_101010011110;
      patterns[43501] = 29'b1_010100111101_101_0_110101001111;
      patterns[43502] = 29'b1_010100111101_110_1_010100111101;
      patterns[43503] = 29'b1_010100111101_111_1_010100111101;
      patterns[43504] = 29'b1_010100111110_000_1_010100111110;
      patterns[43505] = 29'b1_010100111110_001_1_111110010100;
      patterns[43506] = 29'b1_010100111110_010_0_101001111101;
      patterns[43507] = 29'b1_010100111110_011_1_010011111010;
      patterns[43508] = 29'b1_010100111110_100_0_101010011111;
      patterns[43509] = 29'b1_010100111110_101_1_010101001111;
      patterns[43510] = 29'b1_010100111110_110_1_010100111110;
      patterns[43511] = 29'b1_010100111110_111_1_010100111110;
      patterns[43512] = 29'b1_010100111111_000_1_010100111111;
      patterns[43513] = 29'b1_010100111111_001_1_111111010100;
      patterns[43514] = 29'b1_010100111111_010_0_101001111111;
      patterns[43515] = 29'b1_010100111111_011_1_010011111110;
      patterns[43516] = 29'b1_010100111111_100_1_101010011111;
      patterns[43517] = 29'b1_010100111111_101_1_110101001111;
      patterns[43518] = 29'b1_010100111111_110_1_010100111111;
      patterns[43519] = 29'b1_010100111111_111_1_010100111111;
      patterns[43520] = 29'b1_010101000000_000_1_010101000000;
      patterns[43521] = 29'b1_010101000000_001_1_000000010101;
      patterns[43522] = 29'b1_010101000000_010_0_101010000001;
      patterns[43523] = 29'b1_010101000000_011_1_010100000010;
      patterns[43524] = 29'b1_010101000000_100_0_101010100000;
      patterns[43525] = 29'b1_010101000000_101_0_010101010000;
      patterns[43526] = 29'b1_010101000000_110_1_010101000000;
      patterns[43527] = 29'b1_010101000000_111_1_010101000000;
      patterns[43528] = 29'b1_010101000001_000_1_010101000001;
      patterns[43529] = 29'b1_010101000001_001_1_000001010101;
      patterns[43530] = 29'b1_010101000001_010_0_101010000011;
      patterns[43531] = 29'b1_010101000001_011_1_010100000110;
      patterns[43532] = 29'b1_010101000001_100_1_101010100000;
      patterns[43533] = 29'b1_010101000001_101_0_110101010000;
      patterns[43534] = 29'b1_010101000001_110_1_010101000001;
      patterns[43535] = 29'b1_010101000001_111_1_010101000001;
      patterns[43536] = 29'b1_010101000010_000_1_010101000010;
      patterns[43537] = 29'b1_010101000010_001_1_000010010101;
      patterns[43538] = 29'b1_010101000010_010_0_101010000101;
      patterns[43539] = 29'b1_010101000010_011_1_010100001010;
      patterns[43540] = 29'b1_010101000010_100_0_101010100001;
      patterns[43541] = 29'b1_010101000010_101_1_010101010000;
      patterns[43542] = 29'b1_010101000010_110_1_010101000010;
      patterns[43543] = 29'b1_010101000010_111_1_010101000010;
      patterns[43544] = 29'b1_010101000011_000_1_010101000011;
      patterns[43545] = 29'b1_010101000011_001_1_000011010101;
      patterns[43546] = 29'b1_010101000011_010_0_101010000111;
      patterns[43547] = 29'b1_010101000011_011_1_010100001110;
      patterns[43548] = 29'b1_010101000011_100_1_101010100001;
      patterns[43549] = 29'b1_010101000011_101_1_110101010000;
      patterns[43550] = 29'b1_010101000011_110_1_010101000011;
      patterns[43551] = 29'b1_010101000011_111_1_010101000011;
      patterns[43552] = 29'b1_010101000100_000_1_010101000100;
      patterns[43553] = 29'b1_010101000100_001_1_000100010101;
      patterns[43554] = 29'b1_010101000100_010_0_101010001001;
      patterns[43555] = 29'b1_010101000100_011_1_010100010010;
      patterns[43556] = 29'b1_010101000100_100_0_101010100010;
      patterns[43557] = 29'b1_010101000100_101_0_010101010001;
      patterns[43558] = 29'b1_010101000100_110_1_010101000100;
      patterns[43559] = 29'b1_010101000100_111_1_010101000100;
      patterns[43560] = 29'b1_010101000101_000_1_010101000101;
      patterns[43561] = 29'b1_010101000101_001_1_000101010101;
      patterns[43562] = 29'b1_010101000101_010_0_101010001011;
      patterns[43563] = 29'b1_010101000101_011_1_010100010110;
      patterns[43564] = 29'b1_010101000101_100_1_101010100010;
      patterns[43565] = 29'b1_010101000101_101_0_110101010001;
      patterns[43566] = 29'b1_010101000101_110_1_010101000101;
      patterns[43567] = 29'b1_010101000101_111_1_010101000101;
      patterns[43568] = 29'b1_010101000110_000_1_010101000110;
      patterns[43569] = 29'b1_010101000110_001_1_000110010101;
      patterns[43570] = 29'b1_010101000110_010_0_101010001101;
      patterns[43571] = 29'b1_010101000110_011_1_010100011010;
      patterns[43572] = 29'b1_010101000110_100_0_101010100011;
      patterns[43573] = 29'b1_010101000110_101_1_010101010001;
      patterns[43574] = 29'b1_010101000110_110_1_010101000110;
      patterns[43575] = 29'b1_010101000110_111_1_010101000110;
      patterns[43576] = 29'b1_010101000111_000_1_010101000111;
      patterns[43577] = 29'b1_010101000111_001_1_000111010101;
      patterns[43578] = 29'b1_010101000111_010_0_101010001111;
      patterns[43579] = 29'b1_010101000111_011_1_010100011110;
      patterns[43580] = 29'b1_010101000111_100_1_101010100011;
      patterns[43581] = 29'b1_010101000111_101_1_110101010001;
      patterns[43582] = 29'b1_010101000111_110_1_010101000111;
      patterns[43583] = 29'b1_010101000111_111_1_010101000111;
      patterns[43584] = 29'b1_010101001000_000_1_010101001000;
      patterns[43585] = 29'b1_010101001000_001_1_001000010101;
      patterns[43586] = 29'b1_010101001000_010_0_101010010001;
      patterns[43587] = 29'b1_010101001000_011_1_010100100010;
      patterns[43588] = 29'b1_010101001000_100_0_101010100100;
      patterns[43589] = 29'b1_010101001000_101_0_010101010010;
      patterns[43590] = 29'b1_010101001000_110_1_010101001000;
      patterns[43591] = 29'b1_010101001000_111_1_010101001000;
      patterns[43592] = 29'b1_010101001001_000_1_010101001001;
      patterns[43593] = 29'b1_010101001001_001_1_001001010101;
      patterns[43594] = 29'b1_010101001001_010_0_101010010011;
      patterns[43595] = 29'b1_010101001001_011_1_010100100110;
      patterns[43596] = 29'b1_010101001001_100_1_101010100100;
      patterns[43597] = 29'b1_010101001001_101_0_110101010010;
      patterns[43598] = 29'b1_010101001001_110_1_010101001001;
      patterns[43599] = 29'b1_010101001001_111_1_010101001001;
      patterns[43600] = 29'b1_010101001010_000_1_010101001010;
      patterns[43601] = 29'b1_010101001010_001_1_001010010101;
      patterns[43602] = 29'b1_010101001010_010_0_101010010101;
      patterns[43603] = 29'b1_010101001010_011_1_010100101010;
      patterns[43604] = 29'b1_010101001010_100_0_101010100101;
      patterns[43605] = 29'b1_010101001010_101_1_010101010010;
      patterns[43606] = 29'b1_010101001010_110_1_010101001010;
      patterns[43607] = 29'b1_010101001010_111_1_010101001010;
      patterns[43608] = 29'b1_010101001011_000_1_010101001011;
      patterns[43609] = 29'b1_010101001011_001_1_001011010101;
      patterns[43610] = 29'b1_010101001011_010_0_101010010111;
      patterns[43611] = 29'b1_010101001011_011_1_010100101110;
      patterns[43612] = 29'b1_010101001011_100_1_101010100101;
      patterns[43613] = 29'b1_010101001011_101_1_110101010010;
      patterns[43614] = 29'b1_010101001011_110_1_010101001011;
      patterns[43615] = 29'b1_010101001011_111_1_010101001011;
      patterns[43616] = 29'b1_010101001100_000_1_010101001100;
      patterns[43617] = 29'b1_010101001100_001_1_001100010101;
      patterns[43618] = 29'b1_010101001100_010_0_101010011001;
      patterns[43619] = 29'b1_010101001100_011_1_010100110010;
      patterns[43620] = 29'b1_010101001100_100_0_101010100110;
      patterns[43621] = 29'b1_010101001100_101_0_010101010011;
      patterns[43622] = 29'b1_010101001100_110_1_010101001100;
      patterns[43623] = 29'b1_010101001100_111_1_010101001100;
      patterns[43624] = 29'b1_010101001101_000_1_010101001101;
      patterns[43625] = 29'b1_010101001101_001_1_001101010101;
      patterns[43626] = 29'b1_010101001101_010_0_101010011011;
      patterns[43627] = 29'b1_010101001101_011_1_010100110110;
      patterns[43628] = 29'b1_010101001101_100_1_101010100110;
      patterns[43629] = 29'b1_010101001101_101_0_110101010011;
      patterns[43630] = 29'b1_010101001101_110_1_010101001101;
      patterns[43631] = 29'b1_010101001101_111_1_010101001101;
      patterns[43632] = 29'b1_010101001110_000_1_010101001110;
      patterns[43633] = 29'b1_010101001110_001_1_001110010101;
      patterns[43634] = 29'b1_010101001110_010_0_101010011101;
      patterns[43635] = 29'b1_010101001110_011_1_010100111010;
      patterns[43636] = 29'b1_010101001110_100_0_101010100111;
      patterns[43637] = 29'b1_010101001110_101_1_010101010011;
      patterns[43638] = 29'b1_010101001110_110_1_010101001110;
      patterns[43639] = 29'b1_010101001110_111_1_010101001110;
      patterns[43640] = 29'b1_010101001111_000_1_010101001111;
      patterns[43641] = 29'b1_010101001111_001_1_001111010101;
      patterns[43642] = 29'b1_010101001111_010_0_101010011111;
      patterns[43643] = 29'b1_010101001111_011_1_010100111110;
      patterns[43644] = 29'b1_010101001111_100_1_101010100111;
      patterns[43645] = 29'b1_010101001111_101_1_110101010011;
      patterns[43646] = 29'b1_010101001111_110_1_010101001111;
      patterns[43647] = 29'b1_010101001111_111_1_010101001111;
      patterns[43648] = 29'b1_010101010000_000_1_010101010000;
      patterns[43649] = 29'b1_010101010000_001_1_010000010101;
      patterns[43650] = 29'b1_010101010000_010_0_101010100001;
      patterns[43651] = 29'b1_010101010000_011_1_010101000010;
      patterns[43652] = 29'b1_010101010000_100_0_101010101000;
      patterns[43653] = 29'b1_010101010000_101_0_010101010100;
      patterns[43654] = 29'b1_010101010000_110_1_010101010000;
      patterns[43655] = 29'b1_010101010000_111_1_010101010000;
      patterns[43656] = 29'b1_010101010001_000_1_010101010001;
      patterns[43657] = 29'b1_010101010001_001_1_010001010101;
      patterns[43658] = 29'b1_010101010001_010_0_101010100011;
      patterns[43659] = 29'b1_010101010001_011_1_010101000110;
      patterns[43660] = 29'b1_010101010001_100_1_101010101000;
      patterns[43661] = 29'b1_010101010001_101_0_110101010100;
      patterns[43662] = 29'b1_010101010001_110_1_010101010001;
      patterns[43663] = 29'b1_010101010001_111_1_010101010001;
      patterns[43664] = 29'b1_010101010010_000_1_010101010010;
      patterns[43665] = 29'b1_010101010010_001_1_010010010101;
      patterns[43666] = 29'b1_010101010010_010_0_101010100101;
      patterns[43667] = 29'b1_010101010010_011_1_010101001010;
      patterns[43668] = 29'b1_010101010010_100_0_101010101001;
      patterns[43669] = 29'b1_010101010010_101_1_010101010100;
      patterns[43670] = 29'b1_010101010010_110_1_010101010010;
      patterns[43671] = 29'b1_010101010010_111_1_010101010010;
      patterns[43672] = 29'b1_010101010011_000_1_010101010011;
      patterns[43673] = 29'b1_010101010011_001_1_010011010101;
      patterns[43674] = 29'b1_010101010011_010_0_101010100111;
      patterns[43675] = 29'b1_010101010011_011_1_010101001110;
      patterns[43676] = 29'b1_010101010011_100_1_101010101001;
      patterns[43677] = 29'b1_010101010011_101_1_110101010100;
      patterns[43678] = 29'b1_010101010011_110_1_010101010011;
      patterns[43679] = 29'b1_010101010011_111_1_010101010011;
      patterns[43680] = 29'b1_010101010100_000_1_010101010100;
      patterns[43681] = 29'b1_010101010100_001_1_010100010101;
      patterns[43682] = 29'b1_010101010100_010_0_101010101001;
      patterns[43683] = 29'b1_010101010100_011_1_010101010010;
      patterns[43684] = 29'b1_010101010100_100_0_101010101010;
      patterns[43685] = 29'b1_010101010100_101_0_010101010101;
      patterns[43686] = 29'b1_010101010100_110_1_010101010100;
      patterns[43687] = 29'b1_010101010100_111_1_010101010100;
      patterns[43688] = 29'b1_010101010101_000_1_010101010101;
      patterns[43689] = 29'b1_010101010101_001_1_010101010101;
      patterns[43690] = 29'b1_010101010101_010_0_101010101011;
      patterns[43691] = 29'b1_010101010101_011_1_010101010110;
      patterns[43692] = 29'b1_010101010101_100_1_101010101010;
      patterns[43693] = 29'b1_010101010101_101_0_110101010101;
      patterns[43694] = 29'b1_010101010101_110_1_010101010101;
      patterns[43695] = 29'b1_010101010101_111_1_010101010101;
      patterns[43696] = 29'b1_010101010110_000_1_010101010110;
      patterns[43697] = 29'b1_010101010110_001_1_010110010101;
      patterns[43698] = 29'b1_010101010110_010_0_101010101101;
      patterns[43699] = 29'b1_010101010110_011_1_010101011010;
      patterns[43700] = 29'b1_010101010110_100_0_101010101011;
      patterns[43701] = 29'b1_010101010110_101_1_010101010101;
      patterns[43702] = 29'b1_010101010110_110_1_010101010110;
      patterns[43703] = 29'b1_010101010110_111_1_010101010110;
      patterns[43704] = 29'b1_010101010111_000_1_010101010111;
      patterns[43705] = 29'b1_010101010111_001_1_010111010101;
      patterns[43706] = 29'b1_010101010111_010_0_101010101111;
      patterns[43707] = 29'b1_010101010111_011_1_010101011110;
      patterns[43708] = 29'b1_010101010111_100_1_101010101011;
      patterns[43709] = 29'b1_010101010111_101_1_110101010101;
      patterns[43710] = 29'b1_010101010111_110_1_010101010111;
      patterns[43711] = 29'b1_010101010111_111_1_010101010111;
      patterns[43712] = 29'b1_010101011000_000_1_010101011000;
      patterns[43713] = 29'b1_010101011000_001_1_011000010101;
      patterns[43714] = 29'b1_010101011000_010_0_101010110001;
      patterns[43715] = 29'b1_010101011000_011_1_010101100010;
      patterns[43716] = 29'b1_010101011000_100_0_101010101100;
      patterns[43717] = 29'b1_010101011000_101_0_010101010110;
      patterns[43718] = 29'b1_010101011000_110_1_010101011000;
      patterns[43719] = 29'b1_010101011000_111_1_010101011000;
      patterns[43720] = 29'b1_010101011001_000_1_010101011001;
      patterns[43721] = 29'b1_010101011001_001_1_011001010101;
      patterns[43722] = 29'b1_010101011001_010_0_101010110011;
      patterns[43723] = 29'b1_010101011001_011_1_010101100110;
      patterns[43724] = 29'b1_010101011001_100_1_101010101100;
      patterns[43725] = 29'b1_010101011001_101_0_110101010110;
      patterns[43726] = 29'b1_010101011001_110_1_010101011001;
      patterns[43727] = 29'b1_010101011001_111_1_010101011001;
      patterns[43728] = 29'b1_010101011010_000_1_010101011010;
      patterns[43729] = 29'b1_010101011010_001_1_011010010101;
      patterns[43730] = 29'b1_010101011010_010_0_101010110101;
      patterns[43731] = 29'b1_010101011010_011_1_010101101010;
      patterns[43732] = 29'b1_010101011010_100_0_101010101101;
      patterns[43733] = 29'b1_010101011010_101_1_010101010110;
      patterns[43734] = 29'b1_010101011010_110_1_010101011010;
      patterns[43735] = 29'b1_010101011010_111_1_010101011010;
      patterns[43736] = 29'b1_010101011011_000_1_010101011011;
      patterns[43737] = 29'b1_010101011011_001_1_011011010101;
      patterns[43738] = 29'b1_010101011011_010_0_101010110111;
      patterns[43739] = 29'b1_010101011011_011_1_010101101110;
      patterns[43740] = 29'b1_010101011011_100_1_101010101101;
      patterns[43741] = 29'b1_010101011011_101_1_110101010110;
      patterns[43742] = 29'b1_010101011011_110_1_010101011011;
      patterns[43743] = 29'b1_010101011011_111_1_010101011011;
      patterns[43744] = 29'b1_010101011100_000_1_010101011100;
      patterns[43745] = 29'b1_010101011100_001_1_011100010101;
      patterns[43746] = 29'b1_010101011100_010_0_101010111001;
      patterns[43747] = 29'b1_010101011100_011_1_010101110010;
      patterns[43748] = 29'b1_010101011100_100_0_101010101110;
      patterns[43749] = 29'b1_010101011100_101_0_010101010111;
      patterns[43750] = 29'b1_010101011100_110_1_010101011100;
      patterns[43751] = 29'b1_010101011100_111_1_010101011100;
      patterns[43752] = 29'b1_010101011101_000_1_010101011101;
      patterns[43753] = 29'b1_010101011101_001_1_011101010101;
      patterns[43754] = 29'b1_010101011101_010_0_101010111011;
      patterns[43755] = 29'b1_010101011101_011_1_010101110110;
      patterns[43756] = 29'b1_010101011101_100_1_101010101110;
      patterns[43757] = 29'b1_010101011101_101_0_110101010111;
      patterns[43758] = 29'b1_010101011101_110_1_010101011101;
      patterns[43759] = 29'b1_010101011101_111_1_010101011101;
      patterns[43760] = 29'b1_010101011110_000_1_010101011110;
      patterns[43761] = 29'b1_010101011110_001_1_011110010101;
      patterns[43762] = 29'b1_010101011110_010_0_101010111101;
      patterns[43763] = 29'b1_010101011110_011_1_010101111010;
      patterns[43764] = 29'b1_010101011110_100_0_101010101111;
      patterns[43765] = 29'b1_010101011110_101_1_010101010111;
      patterns[43766] = 29'b1_010101011110_110_1_010101011110;
      patterns[43767] = 29'b1_010101011110_111_1_010101011110;
      patterns[43768] = 29'b1_010101011111_000_1_010101011111;
      patterns[43769] = 29'b1_010101011111_001_1_011111010101;
      patterns[43770] = 29'b1_010101011111_010_0_101010111111;
      patterns[43771] = 29'b1_010101011111_011_1_010101111110;
      patterns[43772] = 29'b1_010101011111_100_1_101010101111;
      patterns[43773] = 29'b1_010101011111_101_1_110101010111;
      patterns[43774] = 29'b1_010101011111_110_1_010101011111;
      patterns[43775] = 29'b1_010101011111_111_1_010101011111;
      patterns[43776] = 29'b1_010101100000_000_1_010101100000;
      patterns[43777] = 29'b1_010101100000_001_1_100000010101;
      patterns[43778] = 29'b1_010101100000_010_0_101011000001;
      patterns[43779] = 29'b1_010101100000_011_1_010110000010;
      patterns[43780] = 29'b1_010101100000_100_0_101010110000;
      patterns[43781] = 29'b1_010101100000_101_0_010101011000;
      patterns[43782] = 29'b1_010101100000_110_1_010101100000;
      patterns[43783] = 29'b1_010101100000_111_1_010101100000;
      patterns[43784] = 29'b1_010101100001_000_1_010101100001;
      patterns[43785] = 29'b1_010101100001_001_1_100001010101;
      patterns[43786] = 29'b1_010101100001_010_0_101011000011;
      patterns[43787] = 29'b1_010101100001_011_1_010110000110;
      patterns[43788] = 29'b1_010101100001_100_1_101010110000;
      patterns[43789] = 29'b1_010101100001_101_0_110101011000;
      patterns[43790] = 29'b1_010101100001_110_1_010101100001;
      patterns[43791] = 29'b1_010101100001_111_1_010101100001;
      patterns[43792] = 29'b1_010101100010_000_1_010101100010;
      patterns[43793] = 29'b1_010101100010_001_1_100010010101;
      patterns[43794] = 29'b1_010101100010_010_0_101011000101;
      patterns[43795] = 29'b1_010101100010_011_1_010110001010;
      patterns[43796] = 29'b1_010101100010_100_0_101010110001;
      patterns[43797] = 29'b1_010101100010_101_1_010101011000;
      patterns[43798] = 29'b1_010101100010_110_1_010101100010;
      patterns[43799] = 29'b1_010101100010_111_1_010101100010;
      patterns[43800] = 29'b1_010101100011_000_1_010101100011;
      patterns[43801] = 29'b1_010101100011_001_1_100011010101;
      patterns[43802] = 29'b1_010101100011_010_0_101011000111;
      patterns[43803] = 29'b1_010101100011_011_1_010110001110;
      patterns[43804] = 29'b1_010101100011_100_1_101010110001;
      patterns[43805] = 29'b1_010101100011_101_1_110101011000;
      patterns[43806] = 29'b1_010101100011_110_1_010101100011;
      patterns[43807] = 29'b1_010101100011_111_1_010101100011;
      patterns[43808] = 29'b1_010101100100_000_1_010101100100;
      patterns[43809] = 29'b1_010101100100_001_1_100100010101;
      patterns[43810] = 29'b1_010101100100_010_0_101011001001;
      patterns[43811] = 29'b1_010101100100_011_1_010110010010;
      patterns[43812] = 29'b1_010101100100_100_0_101010110010;
      patterns[43813] = 29'b1_010101100100_101_0_010101011001;
      patterns[43814] = 29'b1_010101100100_110_1_010101100100;
      patterns[43815] = 29'b1_010101100100_111_1_010101100100;
      patterns[43816] = 29'b1_010101100101_000_1_010101100101;
      patterns[43817] = 29'b1_010101100101_001_1_100101010101;
      patterns[43818] = 29'b1_010101100101_010_0_101011001011;
      patterns[43819] = 29'b1_010101100101_011_1_010110010110;
      patterns[43820] = 29'b1_010101100101_100_1_101010110010;
      patterns[43821] = 29'b1_010101100101_101_0_110101011001;
      patterns[43822] = 29'b1_010101100101_110_1_010101100101;
      patterns[43823] = 29'b1_010101100101_111_1_010101100101;
      patterns[43824] = 29'b1_010101100110_000_1_010101100110;
      patterns[43825] = 29'b1_010101100110_001_1_100110010101;
      patterns[43826] = 29'b1_010101100110_010_0_101011001101;
      patterns[43827] = 29'b1_010101100110_011_1_010110011010;
      patterns[43828] = 29'b1_010101100110_100_0_101010110011;
      patterns[43829] = 29'b1_010101100110_101_1_010101011001;
      patterns[43830] = 29'b1_010101100110_110_1_010101100110;
      patterns[43831] = 29'b1_010101100110_111_1_010101100110;
      patterns[43832] = 29'b1_010101100111_000_1_010101100111;
      patterns[43833] = 29'b1_010101100111_001_1_100111010101;
      patterns[43834] = 29'b1_010101100111_010_0_101011001111;
      patterns[43835] = 29'b1_010101100111_011_1_010110011110;
      patterns[43836] = 29'b1_010101100111_100_1_101010110011;
      patterns[43837] = 29'b1_010101100111_101_1_110101011001;
      patterns[43838] = 29'b1_010101100111_110_1_010101100111;
      patterns[43839] = 29'b1_010101100111_111_1_010101100111;
      patterns[43840] = 29'b1_010101101000_000_1_010101101000;
      patterns[43841] = 29'b1_010101101000_001_1_101000010101;
      patterns[43842] = 29'b1_010101101000_010_0_101011010001;
      patterns[43843] = 29'b1_010101101000_011_1_010110100010;
      patterns[43844] = 29'b1_010101101000_100_0_101010110100;
      patterns[43845] = 29'b1_010101101000_101_0_010101011010;
      patterns[43846] = 29'b1_010101101000_110_1_010101101000;
      patterns[43847] = 29'b1_010101101000_111_1_010101101000;
      patterns[43848] = 29'b1_010101101001_000_1_010101101001;
      patterns[43849] = 29'b1_010101101001_001_1_101001010101;
      patterns[43850] = 29'b1_010101101001_010_0_101011010011;
      patterns[43851] = 29'b1_010101101001_011_1_010110100110;
      patterns[43852] = 29'b1_010101101001_100_1_101010110100;
      patterns[43853] = 29'b1_010101101001_101_0_110101011010;
      patterns[43854] = 29'b1_010101101001_110_1_010101101001;
      patterns[43855] = 29'b1_010101101001_111_1_010101101001;
      patterns[43856] = 29'b1_010101101010_000_1_010101101010;
      patterns[43857] = 29'b1_010101101010_001_1_101010010101;
      patterns[43858] = 29'b1_010101101010_010_0_101011010101;
      patterns[43859] = 29'b1_010101101010_011_1_010110101010;
      patterns[43860] = 29'b1_010101101010_100_0_101010110101;
      patterns[43861] = 29'b1_010101101010_101_1_010101011010;
      patterns[43862] = 29'b1_010101101010_110_1_010101101010;
      patterns[43863] = 29'b1_010101101010_111_1_010101101010;
      patterns[43864] = 29'b1_010101101011_000_1_010101101011;
      patterns[43865] = 29'b1_010101101011_001_1_101011010101;
      patterns[43866] = 29'b1_010101101011_010_0_101011010111;
      patterns[43867] = 29'b1_010101101011_011_1_010110101110;
      patterns[43868] = 29'b1_010101101011_100_1_101010110101;
      patterns[43869] = 29'b1_010101101011_101_1_110101011010;
      patterns[43870] = 29'b1_010101101011_110_1_010101101011;
      patterns[43871] = 29'b1_010101101011_111_1_010101101011;
      patterns[43872] = 29'b1_010101101100_000_1_010101101100;
      patterns[43873] = 29'b1_010101101100_001_1_101100010101;
      patterns[43874] = 29'b1_010101101100_010_0_101011011001;
      patterns[43875] = 29'b1_010101101100_011_1_010110110010;
      patterns[43876] = 29'b1_010101101100_100_0_101010110110;
      patterns[43877] = 29'b1_010101101100_101_0_010101011011;
      patterns[43878] = 29'b1_010101101100_110_1_010101101100;
      patterns[43879] = 29'b1_010101101100_111_1_010101101100;
      patterns[43880] = 29'b1_010101101101_000_1_010101101101;
      patterns[43881] = 29'b1_010101101101_001_1_101101010101;
      patterns[43882] = 29'b1_010101101101_010_0_101011011011;
      patterns[43883] = 29'b1_010101101101_011_1_010110110110;
      patterns[43884] = 29'b1_010101101101_100_1_101010110110;
      patterns[43885] = 29'b1_010101101101_101_0_110101011011;
      patterns[43886] = 29'b1_010101101101_110_1_010101101101;
      patterns[43887] = 29'b1_010101101101_111_1_010101101101;
      patterns[43888] = 29'b1_010101101110_000_1_010101101110;
      patterns[43889] = 29'b1_010101101110_001_1_101110010101;
      patterns[43890] = 29'b1_010101101110_010_0_101011011101;
      patterns[43891] = 29'b1_010101101110_011_1_010110111010;
      patterns[43892] = 29'b1_010101101110_100_0_101010110111;
      patterns[43893] = 29'b1_010101101110_101_1_010101011011;
      patterns[43894] = 29'b1_010101101110_110_1_010101101110;
      patterns[43895] = 29'b1_010101101110_111_1_010101101110;
      patterns[43896] = 29'b1_010101101111_000_1_010101101111;
      patterns[43897] = 29'b1_010101101111_001_1_101111010101;
      patterns[43898] = 29'b1_010101101111_010_0_101011011111;
      patterns[43899] = 29'b1_010101101111_011_1_010110111110;
      patterns[43900] = 29'b1_010101101111_100_1_101010110111;
      patterns[43901] = 29'b1_010101101111_101_1_110101011011;
      patterns[43902] = 29'b1_010101101111_110_1_010101101111;
      patterns[43903] = 29'b1_010101101111_111_1_010101101111;
      patterns[43904] = 29'b1_010101110000_000_1_010101110000;
      patterns[43905] = 29'b1_010101110000_001_1_110000010101;
      patterns[43906] = 29'b1_010101110000_010_0_101011100001;
      patterns[43907] = 29'b1_010101110000_011_1_010111000010;
      patterns[43908] = 29'b1_010101110000_100_0_101010111000;
      patterns[43909] = 29'b1_010101110000_101_0_010101011100;
      patterns[43910] = 29'b1_010101110000_110_1_010101110000;
      patterns[43911] = 29'b1_010101110000_111_1_010101110000;
      patterns[43912] = 29'b1_010101110001_000_1_010101110001;
      patterns[43913] = 29'b1_010101110001_001_1_110001010101;
      patterns[43914] = 29'b1_010101110001_010_0_101011100011;
      patterns[43915] = 29'b1_010101110001_011_1_010111000110;
      patterns[43916] = 29'b1_010101110001_100_1_101010111000;
      patterns[43917] = 29'b1_010101110001_101_0_110101011100;
      patterns[43918] = 29'b1_010101110001_110_1_010101110001;
      patterns[43919] = 29'b1_010101110001_111_1_010101110001;
      patterns[43920] = 29'b1_010101110010_000_1_010101110010;
      patterns[43921] = 29'b1_010101110010_001_1_110010010101;
      patterns[43922] = 29'b1_010101110010_010_0_101011100101;
      patterns[43923] = 29'b1_010101110010_011_1_010111001010;
      patterns[43924] = 29'b1_010101110010_100_0_101010111001;
      patterns[43925] = 29'b1_010101110010_101_1_010101011100;
      patterns[43926] = 29'b1_010101110010_110_1_010101110010;
      patterns[43927] = 29'b1_010101110010_111_1_010101110010;
      patterns[43928] = 29'b1_010101110011_000_1_010101110011;
      patterns[43929] = 29'b1_010101110011_001_1_110011010101;
      patterns[43930] = 29'b1_010101110011_010_0_101011100111;
      patterns[43931] = 29'b1_010101110011_011_1_010111001110;
      patterns[43932] = 29'b1_010101110011_100_1_101010111001;
      patterns[43933] = 29'b1_010101110011_101_1_110101011100;
      patterns[43934] = 29'b1_010101110011_110_1_010101110011;
      patterns[43935] = 29'b1_010101110011_111_1_010101110011;
      patterns[43936] = 29'b1_010101110100_000_1_010101110100;
      patterns[43937] = 29'b1_010101110100_001_1_110100010101;
      patterns[43938] = 29'b1_010101110100_010_0_101011101001;
      patterns[43939] = 29'b1_010101110100_011_1_010111010010;
      patterns[43940] = 29'b1_010101110100_100_0_101010111010;
      patterns[43941] = 29'b1_010101110100_101_0_010101011101;
      patterns[43942] = 29'b1_010101110100_110_1_010101110100;
      patterns[43943] = 29'b1_010101110100_111_1_010101110100;
      patterns[43944] = 29'b1_010101110101_000_1_010101110101;
      patterns[43945] = 29'b1_010101110101_001_1_110101010101;
      patterns[43946] = 29'b1_010101110101_010_0_101011101011;
      patterns[43947] = 29'b1_010101110101_011_1_010111010110;
      patterns[43948] = 29'b1_010101110101_100_1_101010111010;
      patterns[43949] = 29'b1_010101110101_101_0_110101011101;
      patterns[43950] = 29'b1_010101110101_110_1_010101110101;
      patterns[43951] = 29'b1_010101110101_111_1_010101110101;
      patterns[43952] = 29'b1_010101110110_000_1_010101110110;
      patterns[43953] = 29'b1_010101110110_001_1_110110010101;
      patterns[43954] = 29'b1_010101110110_010_0_101011101101;
      patterns[43955] = 29'b1_010101110110_011_1_010111011010;
      patterns[43956] = 29'b1_010101110110_100_0_101010111011;
      patterns[43957] = 29'b1_010101110110_101_1_010101011101;
      patterns[43958] = 29'b1_010101110110_110_1_010101110110;
      patterns[43959] = 29'b1_010101110110_111_1_010101110110;
      patterns[43960] = 29'b1_010101110111_000_1_010101110111;
      patterns[43961] = 29'b1_010101110111_001_1_110111010101;
      patterns[43962] = 29'b1_010101110111_010_0_101011101111;
      patterns[43963] = 29'b1_010101110111_011_1_010111011110;
      patterns[43964] = 29'b1_010101110111_100_1_101010111011;
      patterns[43965] = 29'b1_010101110111_101_1_110101011101;
      patterns[43966] = 29'b1_010101110111_110_1_010101110111;
      patterns[43967] = 29'b1_010101110111_111_1_010101110111;
      patterns[43968] = 29'b1_010101111000_000_1_010101111000;
      patterns[43969] = 29'b1_010101111000_001_1_111000010101;
      patterns[43970] = 29'b1_010101111000_010_0_101011110001;
      patterns[43971] = 29'b1_010101111000_011_1_010111100010;
      patterns[43972] = 29'b1_010101111000_100_0_101010111100;
      patterns[43973] = 29'b1_010101111000_101_0_010101011110;
      patterns[43974] = 29'b1_010101111000_110_1_010101111000;
      patterns[43975] = 29'b1_010101111000_111_1_010101111000;
      patterns[43976] = 29'b1_010101111001_000_1_010101111001;
      patterns[43977] = 29'b1_010101111001_001_1_111001010101;
      patterns[43978] = 29'b1_010101111001_010_0_101011110011;
      patterns[43979] = 29'b1_010101111001_011_1_010111100110;
      patterns[43980] = 29'b1_010101111001_100_1_101010111100;
      patterns[43981] = 29'b1_010101111001_101_0_110101011110;
      patterns[43982] = 29'b1_010101111001_110_1_010101111001;
      patterns[43983] = 29'b1_010101111001_111_1_010101111001;
      patterns[43984] = 29'b1_010101111010_000_1_010101111010;
      patterns[43985] = 29'b1_010101111010_001_1_111010010101;
      patterns[43986] = 29'b1_010101111010_010_0_101011110101;
      patterns[43987] = 29'b1_010101111010_011_1_010111101010;
      patterns[43988] = 29'b1_010101111010_100_0_101010111101;
      patterns[43989] = 29'b1_010101111010_101_1_010101011110;
      patterns[43990] = 29'b1_010101111010_110_1_010101111010;
      patterns[43991] = 29'b1_010101111010_111_1_010101111010;
      patterns[43992] = 29'b1_010101111011_000_1_010101111011;
      patterns[43993] = 29'b1_010101111011_001_1_111011010101;
      patterns[43994] = 29'b1_010101111011_010_0_101011110111;
      patterns[43995] = 29'b1_010101111011_011_1_010111101110;
      patterns[43996] = 29'b1_010101111011_100_1_101010111101;
      patterns[43997] = 29'b1_010101111011_101_1_110101011110;
      patterns[43998] = 29'b1_010101111011_110_1_010101111011;
      patterns[43999] = 29'b1_010101111011_111_1_010101111011;
      patterns[44000] = 29'b1_010101111100_000_1_010101111100;
      patterns[44001] = 29'b1_010101111100_001_1_111100010101;
      patterns[44002] = 29'b1_010101111100_010_0_101011111001;
      patterns[44003] = 29'b1_010101111100_011_1_010111110010;
      patterns[44004] = 29'b1_010101111100_100_0_101010111110;
      patterns[44005] = 29'b1_010101111100_101_0_010101011111;
      patterns[44006] = 29'b1_010101111100_110_1_010101111100;
      patterns[44007] = 29'b1_010101111100_111_1_010101111100;
      patterns[44008] = 29'b1_010101111101_000_1_010101111101;
      patterns[44009] = 29'b1_010101111101_001_1_111101010101;
      patterns[44010] = 29'b1_010101111101_010_0_101011111011;
      patterns[44011] = 29'b1_010101111101_011_1_010111110110;
      patterns[44012] = 29'b1_010101111101_100_1_101010111110;
      patterns[44013] = 29'b1_010101111101_101_0_110101011111;
      patterns[44014] = 29'b1_010101111101_110_1_010101111101;
      patterns[44015] = 29'b1_010101111101_111_1_010101111101;
      patterns[44016] = 29'b1_010101111110_000_1_010101111110;
      patterns[44017] = 29'b1_010101111110_001_1_111110010101;
      patterns[44018] = 29'b1_010101111110_010_0_101011111101;
      patterns[44019] = 29'b1_010101111110_011_1_010111111010;
      patterns[44020] = 29'b1_010101111110_100_0_101010111111;
      patterns[44021] = 29'b1_010101111110_101_1_010101011111;
      patterns[44022] = 29'b1_010101111110_110_1_010101111110;
      patterns[44023] = 29'b1_010101111110_111_1_010101111110;
      patterns[44024] = 29'b1_010101111111_000_1_010101111111;
      patterns[44025] = 29'b1_010101111111_001_1_111111010101;
      patterns[44026] = 29'b1_010101111111_010_0_101011111111;
      patterns[44027] = 29'b1_010101111111_011_1_010111111110;
      patterns[44028] = 29'b1_010101111111_100_1_101010111111;
      patterns[44029] = 29'b1_010101111111_101_1_110101011111;
      patterns[44030] = 29'b1_010101111111_110_1_010101111111;
      patterns[44031] = 29'b1_010101111111_111_1_010101111111;
      patterns[44032] = 29'b1_010110000000_000_1_010110000000;
      patterns[44033] = 29'b1_010110000000_001_1_000000010110;
      patterns[44034] = 29'b1_010110000000_010_0_101100000001;
      patterns[44035] = 29'b1_010110000000_011_1_011000000010;
      patterns[44036] = 29'b1_010110000000_100_0_101011000000;
      patterns[44037] = 29'b1_010110000000_101_0_010101100000;
      patterns[44038] = 29'b1_010110000000_110_1_010110000000;
      patterns[44039] = 29'b1_010110000000_111_1_010110000000;
      patterns[44040] = 29'b1_010110000001_000_1_010110000001;
      patterns[44041] = 29'b1_010110000001_001_1_000001010110;
      patterns[44042] = 29'b1_010110000001_010_0_101100000011;
      patterns[44043] = 29'b1_010110000001_011_1_011000000110;
      patterns[44044] = 29'b1_010110000001_100_1_101011000000;
      patterns[44045] = 29'b1_010110000001_101_0_110101100000;
      patterns[44046] = 29'b1_010110000001_110_1_010110000001;
      patterns[44047] = 29'b1_010110000001_111_1_010110000001;
      patterns[44048] = 29'b1_010110000010_000_1_010110000010;
      patterns[44049] = 29'b1_010110000010_001_1_000010010110;
      patterns[44050] = 29'b1_010110000010_010_0_101100000101;
      patterns[44051] = 29'b1_010110000010_011_1_011000001010;
      patterns[44052] = 29'b1_010110000010_100_0_101011000001;
      patterns[44053] = 29'b1_010110000010_101_1_010101100000;
      patterns[44054] = 29'b1_010110000010_110_1_010110000010;
      patterns[44055] = 29'b1_010110000010_111_1_010110000010;
      patterns[44056] = 29'b1_010110000011_000_1_010110000011;
      patterns[44057] = 29'b1_010110000011_001_1_000011010110;
      patterns[44058] = 29'b1_010110000011_010_0_101100000111;
      patterns[44059] = 29'b1_010110000011_011_1_011000001110;
      patterns[44060] = 29'b1_010110000011_100_1_101011000001;
      patterns[44061] = 29'b1_010110000011_101_1_110101100000;
      patterns[44062] = 29'b1_010110000011_110_1_010110000011;
      patterns[44063] = 29'b1_010110000011_111_1_010110000011;
      patterns[44064] = 29'b1_010110000100_000_1_010110000100;
      patterns[44065] = 29'b1_010110000100_001_1_000100010110;
      patterns[44066] = 29'b1_010110000100_010_0_101100001001;
      patterns[44067] = 29'b1_010110000100_011_1_011000010010;
      patterns[44068] = 29'b1_010110000100_100_0_101011000010;
      patterns[44069] = 29'b1_010110000100_101_0_010101100001;
      patterns[44070] = 29'b1_010110000100_110_1_010110000100;
      patterns[44071] = 29'b1_010110000100_111_1_010110000100;
      patterns[44072] = 29'b1_010110000101_000_1_010110000101;
      patterns[44073] = 29'b1_010110000101_001_1_000101010110;
      patterns[44074] = 29'b1_010110000101_010_0_101100001011;
      patterns[44075] = 29'b1_010110000101_011_1_011000010110;
      patterns[44076] = 29'b1_010110000101_100_1_101011000010;
      patterns[44077] = 29'b1_010110000101_101_0_110101100001;
      patterns[44078] = 29'b1_010110000101_110_1_010110000101;
      patterns[44079] = 29'b1_010110000101_111_1_010110000101;
      patterns[44080] = 29'b1_010110000110_000_1_010110000110;
      patterns[44081] = 29'b1_010110000110_001_1_000110010110;
      patterns[44082] = 29'b1_010110000110_010_0_101100001101;
      patterns[44083] = 29'b1_010110000110_011_1_011000011010;
      patterns[44084] = 29'b1_010110000110_100_0_101011000011;
      patterns[44085] = 29'b1_010110000110_101_1_010101100001;
      patterns[44086] = 29'b1_010110000110_110_1_010110000110;
      patterns[44087] = 29'b1_010110000110_111_1_010110000110;
      patterns[44088] = 29'b1_010110000111_000_1_010110000111;
      patterns[44089] = 29'b1_010110000111_001_1_000111010110;
      patterns[44090] = 29'b1_010110000111_010_0_101100001111;
      patterns[44091] = 29'b1_010110000111_011_1_011000011110;
      patterns[44092] = 29'b1_010110000111_100_1_101011000011;
      patterns[44093] = 29'b1_010110000111_101_1_110101100001;
      patterns[44094] = 29'b1_010110000111_110_1_010110000111;
      patterns[44095] = 29'b1_010110000111_111_1_010110000111;
      patterns[44096] = 29'b1_010110001000_000_1_010110001000;
      patterns[44097] = 29'b1_010110001000_001_1_001000010110;
      patterns[44098] = 29'b1_010110001000_010_0_101100010001;
      patterns[44099] = 29'b1_010110001000_011_1_011000100010;
      patterns[44100] = 29'b1_010110001000_100_0_101011000100;
      patterns[44101] = 29'b1_010110001000_101_0_010101100010;
      patterns[44102] = 29'b1_010110001000_110_1_010110001000;
      patterns[44103] = 29'b1_010110001000_111_1_010110001000;
      patterns[44104] = 29'b1_010110001001_000_1_010110001001;
      patterns[44105] = 29'b1_010110001001_001_1_001001010110;
      patterns[44106] = 29'b1_010110001001_010_0_101100010011;
      patterns[44107] = 29'b1_010110001001_011_1_011000100110;
      patterns[44108] = 29'b1_010110001001_100_1_101011000100;
      patterns[44109] = 29'b1_010110001001_101_0_110101100010;
      patterns[44110] = 29'b1_010110001001_110_1_010110001001;
      patterns[44111] = 29'b1_010110001001_111_1_010110001001;
      patterns[44112] = 29'b1_010110001010_000_1_010110001010;
      patterns[44113] = 29'b1_010110001010_001_1_001010010110;
      patterns[44114] = 29'b1_010110001010_010_0_101100010101;
      patterns[44115] = 29'b1_010110001010_011_1_011000101010;
      patterns[44116] = 29'b1_010110001010_100_0_101011000101;
      patterns[44117] = 29'b1_010110001010_101_1_010101100010;
      patterns[44118] = 29'b1_010110001010_110_1_010110001010;
      patterns[44119] = 29'b1_010110001010_111_1_010110001010;
      patterns[44120] = 29'b1_010110001011_000_1_010110001011;
      patterns[44121] = 29'b1_010110001011_001_1_001011010110;
      patterns[44122] = 29'b1_010110001011_010_0_101100010111;
      patterns[44123] = 29'b1_010110001011_011_1_011000101110;
      patterns[44124] = 29'b1_010110001011_100_1_101011000101;
      patterns[44125] = 29'b1_010110001011_101_1_110101100010;
      patterns[44126] = 29'b1_010110001011_110_1_010110001011;
      patterns[44127] = 29'b1_010110001011_111_1_010110001011;
      patterns[44128] = 29'b1_010110001100_000_1_010110001100;
      patterns[44129] = 29'b1_010110001100_001_1_001100010110;
      patterns[44130] = 29'b1_010110001100_010_0_101100011001;
      patterns[44131] = 29'b1_010110001100_011_1_011000110010;
      patterns[44132] = 29'b1_010110001100_100_0_101011000110;
      patterns[44133] = 29'b1_010110001100_101_0_010101100011;
      patterns[44134] = 29'b1_010110001100_110_1_010110001100;
      patterns[44135] = 29'b1_010110001100_111_1_010110001100;
      patterns[44136] = 29'b1_010110001101_000_1_010110001101;
      patterns[44137] = 29'b1_010110001101_001_1_001101010110;
      patterns[44138] = 29'b1_010110001101_010_0_101100011011;
      patterns[44139] = 29'b1_010110001101_011_1_011000110110;
      patterns[44140] = 29'b1_010110001101_100_1_101011000110;
      patterns[44141] = 29'b1_010110001101_101_0_110101100011;
      patterns[44142] = 29'b1_010110001101_110_1_010110001101;
      patterns[44143] = 29'b1_010110001101_111_1_010110001101;
      patterns[44144] = 29'b1_010110001110_000_1_010110001110;
      patterns[44145] = 29'b1_010110001110_001_1_001110010110;
      patterns[44146] = 29'b1_010110001110_010_0_101100011101;
      patterns[44147] = 29'b1_010110001110_011_1_011000111010;
      patterns[44148] = 29'b1_010110001110_100_0_101011000111;
      patterns[44149] = 29'b1_010110001110_101_1_010101100011;
      patterns[44150] = 29'b1_010110001110_110_1_010110001110;
      patterns[44151] = 29'b1_010110001110_111_1_010110001110;
      patterns[44152] = 29'b1_010110001111_000_1_010110001111;
      patterns[44153] = 29'b1_010110001111_001_1_001111010110;
      patterns[44154] = 29'b1_010110001111_010_0_101100011111;
      patterns[44155] = 29'b1_010110001111_011_1_011000111110;
      patterns[44156] = 29'b1_010110001111_100_1_101011000111;
      patterns[44157] = 29'b1_010110001111_101_1_110101100011;
      patterns[44158] = 29'b1_010110001111_110_1_010110001111;
      patterns[44159] = 29'b1_010110001111_111_1_010110001111;
      patterns[44160] = 29'b1_010110010000_000_1_010110010000;
      patterns[44161] = 29'b1_010110010000_001_1_010000010110;
      patterns[44162] = 29'b1_010110010000_010_0_101100100001;
      patterns[44163] = 29'b1_010110010000_011_1_011001000010;
      patterns[44164] = 29'b1_010110010000_100_0_101011001000;
      patterns[44165] = 29'b1_010110010000_101_0_010101100100;
      patterns[44166] = 29'b1_010110010000_110_1_010110010000;
      patterns[44167] = 29'b1_010110010000_111_1_010110010000;
      patterns[44168] = 29'b1_010110010001_000_1_010110010001;
      patterns[44169] = 29'b1_010110010001_001_1_010001010110;
      patterns[44170] = 29'b1_010110010001_010_0_101100100011;
      patterns[44171] = 29'b1_010110010001_011_1_011001000110;
      patterns[44172] = 29'b1_010110010001_100_1_101011001000;
      patterns[44173] = 29'b1_010110010001_101_0_110101100100;
      patterns[44174] = 29'b1_010110010001_110_1_010110010001;
      patterns[44175] = 29'b1_010110010001_111_1_010110010001;
      patterns[44176] = 29'b1_010110010010_000_1_010110010010;
      patterns[44177] = 29'b1_010110010010_001_1_010010010110;
      patterns[44178] = 29'b1_010110010010_010_0_101100100101;
      patterns[44179] = 29'b1_010110010010_011_1_011001001010;
      patterns[44180] = 29'b1_010110010010_100_0_101011001001;
      patterns[44181] = 29'b1_010110010010_101_1_010101100100;
      patterns[44182] = 29'b1_010110010010_110_1_010110010010;
      patterns[44183] = 29'b1_010110010010_111_1_010110010010;
      patterns[44184] = 29'b1_010110010011_000_1_010110010011;
      patterns[44185] = 29'b1_010110010011_001_1_010011010110;
      patterns[44186] = 29'b1_010110010011_010_0_101100100111;
      patterns[44187] = 29'b1_010110010011_011_1_011001001110;
      patterns[44188] = 29'b1_010110010011_100_1_101011001001;
      patterns[44189] = 29'b1_010110010011_101_1_110101100100;
      patterns[44190] = 29'b1_010110010011_110_1_010110010011;
      patterns[44191] = 29'b1_010110010011_111_1_010110010011;
      patterns[44192] = 29'b1_010110010100_000_1_010110010100;
      patterns[44193] = 29'b1_010110010100_001_1_010100010110;
      patterns[44194] = 29'b1_010110010100_010_0_101100101001;
      patterns[44195] = 29'b1_010110010100_011_1_011001010010;
      patterns[44196] = 29'b1_010110010100_100_0_101011001010;
      patterns[44197] = 29'b1_010110010100_101_0_010101100101;
      patterns[44198] = 29'b1_010110010100_110_1_010110010100;
      patterns[44199] = 29'b1_010110010100_111_1_010110010100;
      patterns[44200] = 29'b1_010110010101_000_1_010110010101;
      patterns[44201] = 29'b1_010110010101_001_1_010101010110;
      patterns[44202] = 29'b1_010110010101_010_0_101100101011;
      patterns[44203] = 29'b1_010110010101_011_1_011001010110;
      patterns[44204] = 29'b1_010110010101_100_1_101011001010;
      patterns[44205] = 29'b1_010110010101_101_0_110101100101;
      patterns[44206] = 29'b1_010110010101_110_1_010110010101;
      patterns[44207] = 29'b1_010110010101_111_1_010110010101;
      patterns[44208] = 29'b1_010110010110_000_1_010110010110;
      patterns[44209] = 29'b1_010110010110_001_1_010110010110;
      patterns[44210] = 29'b1_010110010110_010_0_101100101101;
      patterns[44211] = 29'b1_010110010110_011_1_011001011010;
      patterns[44212] = 29'b1_010110010110_100_0_101011001011;
      patterns[44213] = 29'b1_010110010110_101_1_010101100101;
      patterns[44214] = 29'b1_010110010110_110_1_010110010110;
      patterns[44215] = 29'b1_010110010110_111_1_010110010110;
      patterns[44216] = 29'b1_010110010111_000_1_010110010111;
      patterns[44217] = 29'b1_010110010111_001_1_010111010110;
      patterns[44218] = 29'b1_010110010111_010_0_101100101111;
      patterns[44219] = 29'b1_010110010111_011_1_011001011110;
      patterns[44220] = 29'b1_010110010111_100_1_101011001011;
      patterns[44221] = 29'b1_010110010111_101_1_110101100101;
      patterns[44222] = 29'b1_010110010111_110_1_010110010111;
      patterns[44223] = 29'b1_010110010111_111_1_010110010111;
      patterns[44224] = 29'b1_010110011000_000_1_010110011000;
      patterns[44225] = 29'b1_010110011000_001_1_011000010110;
      patterns[44226] = 29'b1_010110011000_010_0_101100110001;
      patterns[44227] = 29'b1_010110011000_011_1_011001100010;
      patterns[44228] = 29'b1_010110011000_100_0_101011001100;
      patterns[44229] = 29'b1_010110011000_101_0_010101100110;
      patterns[44230] = 29'b1_010110011000_110_1_010110011000;
      patterns[44231] = 29'b1_010110011000_111_1_010110011000;
      patterns[44232] = 29'b1_010110011001_000_1_010110011001;
      patterns[44233] = 29'b1_010110011001_001_1_011001010110;
      patterns[44234] = 29'b1_010110011001_010_0_101100110011;
      patterns[44235] = 29'b1_010110011001_011_1_011001100110;
      patterns[44236] = 29'b1_010110011001_100_1_101011001100;
      patterns[44237] = 29'b1_010110011001_101_0_110101100110;
      patterns[44238] = 29'b1_010110011001_110_1_010110011001;
      patterns[44239] = 29'b1_010110011001_111_1_010110011001;
      patterns[44240] = 29'b1_010110011010_000_1_010110011010;
      patterns[44241] = 29'b1_010110011010_001_1_011010010110;
      patterns[44242] = 29'b1_010110011010_010_0_101100110101;
      patterns[44243] = 29'b1_010110011010_011_1_011001101010;
      patterns[44244] = 29'b1_010110011010_100_0_101011001101;
      patterns[44245] = 29'b1_010110011010_101_1_010101100110;
      patterns[44246] = 29'b1_010110011010_110_1_010110011010;
      patterns[44247] = 29'b1_010110011010_111_1_010110011010;
      patterns[44248] = 29'b1_010110011011_000_1_010110011011;
      patterns[44249] = 29'b1_010110011011_001_1_011011010110;
      patterns[44250] = 29'b1_010110011011_010_0_101100110111;
      patterns[44251] = 29'b1_010110011011_011_1_011001101110;
      patterns[44252] = 29'b1_010110011011_100_1_101011001101;
      patterns[44253] = 29'b1_010110011011_101_1_110101100110;
      patterns[44254] = 29'b1_010110011011_110_1_010110011011;
      patterns[44255] = 29'b1_010110011011_111_1_010110011011;
      patterns[44256] = 29'b1_010110011100_000_1_010110011100;
      patterns[44257] = 29'b1_010110011100_001_1_011100010110;
      patterns[44258] = 29'b1_010110011100_010_0_101100111001;
      patterns[44259] = 29'b1_010110011100_011_1_011001110010;
      patterns[44260] = 29'b1_010110011100_100_0_101011001110;
      patterns[44261] = 29'b1_010110011100_101_0_010101100111;
      patterns[44262] = 29'b1_010110011100_110_1_010110011100;
      patterns[44263] = 29'b1_010110011100_111_1_010110011100;
      patterns[44264] = 29'b1_010110011101_000_1_010110011101;
      patterns[44265] = 29'b1_010110011101_001_1_011101010110;
      patterns[44266] = 29'b1_010110011101_010_0_101100111011;
      patterns[44267] = 29'b1_010110011101_011_1_011001110110;
      patterns[44268] = 29'b1_010110011101_100_1_101011001110;
      patterns[44269] = 29'b1_010110011101_101_0_110101100111;
      patterns[44270] = 29'b1_010110011101_110_1_010110011101;
      patterns[44271] = 29'b1_010110011101_111_1_010110011101;
      patterns[44272] = 29'b1_010110011110_000_1_010110011110;
      patterns[44273] = 29'b1_010110011110_001_1_011110010110;
      patterns[44274] = 29'b1_010110011110_010_0_101100111101;
      patterns[44275] = 29'b1_010110011110_011_1_011001111010;
      patterns[44276] = 29'b1_010110011110_100_0_101011001111;
      patterns[44277] = 29'b1_010110011110_101_1_010101100111;
      patterns[44278] = 29'b1_010110011110_110_1_010110011110;
      patterns[44279] = 29'b1_010110011110_111_1_010110011110;
      patterns[44280] = 29'b1_010110011111_000_1_010110011111;
      patterns[44281] = 29'b1_010110011111_001_1_011111010110;
      patterns[44282] = 29'b1_010110011111_010_0_101100111111;
      patterns[44283] = 29'b1_010110011111_011_1_011001111110;
      patterns[44284] = 29'b1_010110011111_100_1_101011001111;
      patterns[44285] = 29'b1_010110011111_101_1_110101100111;
      patterns[44286] = 29'b1_010110011111_110_1_010110011111;
      patterns[44287] = 29'b1_010110011111_111_1_010110011111;
      patterns[44288] = 29'b1_010110100000_000_1_010110100000;
      patterns[44289] = 29'b1_010110100000_001_1_100000010110;
      patterns[44290] = 29'b1_010110100000_010_0_101101000001;
      patterns[44291] = 29'b1_010110100000_011_1_011010000010;
      patterns[44292] = 29'b1_010110100000_100_0_101011010000;
      patterns[44293] = 29'b1_010110100000_101_0_010101101000;
      patterns[44294] = 29'b1_010110100000_110_1_010110100000;
      patterns[44295] = 29'b1_010110100000_111_1_010110100000;
      patterns[44296] = 29'b1_010110100001_000_1_010110100001;
      patterns[44297] = 29'b1_010110100001_001_1_100001010110;
      patterns[44298] = 29'b1_010110100001_010_0_101101000011;
      patterns[44299] = 29'b1_010110100001_011_1_011010000110;
      patterns[44300] = 29'b1_010110100001_100_1_101011010000;
      patterns[44301] = 29'b1_010110100001_101_0_110101101000;
      patterns[44302] = 29'b1_010110100001_110_1_010110100001;
      patterns[44303] = 29'b1_010110100001_111_1_010110100001;
      patterns[44304] = 29'b1_010110100010_000_1_010110100010;
      patterns[44305] = 29'b1_010110100010_001_1_100010010110;
      patterns[44306] = 29'b1_010110100010_010_0_101101000101;
      patterns[44307] = 29'b1_010110100010_011_1_011010001010;
      patterns[44308] = 29'b1_010110100010_100_0_101011010001;
      patterns[44309] = 29'b1_010110100010_101_1_010101101000;
      patterns[44310] = 29'b1_010110100010_110_1_010110100010;
      patterns[44311] = 29'b1_010110100010_111_1_010110100010;
      patterns[44312] = 29'b1_010110100011_000_1_010110100011;
      patterns[44313] = 29'b1_010110100011_001_1_100011010110;
      patterns[44314] = 29'b1_010110100011_010_0_101101000111;
      patterns[44315] = 29'b1_010110100011_011_1_011010001110;
      patterns[44316] = 29'b1_010110100011_100_1_101011010001;
      patterns[44317] = 29'b1_010110100011_101_1_110101101000;
      patterns[44318] = 29'b1_010110100011_110_1_010110100011;
      patterns[44319] = 29'b1_010110100011_111_1_010110100011;
      patterns[44320] = 29'b1_010110100100_000_1_010110100100;
      patterns[44321] = 29'b1_010110100100_001_1_100100010110;
      patterns[44322] = 29'b1_010110100100_010_0_101101001001;
      patterns[44323] = 29'b1_010110100100_011_1_011010010010;
      patterns[44324] = 29'b1_010110100100_100_0_101011010010;
      patterns[44325] = 29'b1_010110100100_101_0_010101101001;
      patterns[44326] = 29'b1_010110100100_110_1_010110100100;
      patterns[44327] = 29'b1_010110100100_111_1_010110100100;
      patterns[44328] = 29'b1_010110100101_000_1_010110100101;
      patterns[44329] = 29'b1_010110100101_001_1_100101010110;
      patterns[44330] = 29'b1_010110100101_010_0_101101001011;
      patterns[44331] = 29'b1_010110100101_011_1_011010010110;
      patterns[44332] = 29'b1_010110100101_100_1_101011010010;
      patterns[44333] = 29'b1_010110100101_101_0_110101101001;
      patterns[44334] = 29'b1_010110100101_110_1_010110100101;
      patterns[44335] = 29'b1_010110100101_111_1_010110100101;
      patterns[44336] = 29'b1_010110100110_000_1_010110100110;
      patterns[44337] = 29'b1_010110100110_001_1_100110010110;
      patterns[44338] = 29'b1_010110100110_010_0_101101001101;
      patterns[44339] = 29'b1_010110100110_011_1_011010011010;
      patterns[44340] = 29'b1_010110100110_100_0_101011010011;
      patterns[44341] = 29'b1_010110100110_101_1_010101101001;
      patterns[44342] = 29'b1_010110100110_110_1_010110100110;
      patterns[44343] = 29'b1_010110100110_111_1_010110100110;
      patterns[44344] = 29'b1_010110100111_000_1_010110100111;
      patterns[44345] = 29'b1_010110100111_001_1_100111010110;
      patterns[44346] = 29'b1_010110100111_010_0_101101001111;
      patterns[44347] = 29'b1_010110100111_011_1_011010011110;
      patterns[44348] = 29'b1_010110100111_100_1_101011010011;
      patterns[44349] = 29'b1_010110100111_101_1_110101101001;
      patterns[44350] = 29'b1_010110100111_110_1_010110100111;
      patterns[44351] = 29'b1_010110100111_111_1_010110100111;
      patterns[44352] = 29'b1_010110101000_000_1_010110101000;
      patterns[44353] = 29'b1_010110101000_001_1_101000010110;
      patterns[44354] = 29'b1_010110101000_010_0_101101010001;
      patterns[44355] = 29'b1_010110101000_011_1_011010100010;
      patterns[44356] = 29'b1_010110101000_100_0_101011010100;
      patterns[44357] = 29'b1_010110101000_101_0_010101101010;
      patterns[44358] = 29'b1_010110101000_110_1_010110101000;
      patterns[44359] = 29'b1_010110101000_111_1_010110101000;
      patterns[44360] = 29'b1_010110101001_000_1_010110101001;
      patterns[44361] = 29'b1_010110101001_001_1_101001010110;
      patterns[44362] = 29'b1_010110101001_010_0_101101010011;
      patterns[44363] = 29'b1_010110101001_011_1_011010100110;
      patterns[44364] = 29'b1_010110101001_100_1_101011010100;
      patterns[44365] = 29'b1_010110101001_101_0_110101101010;
      patterns[44366] = 29'b1_010110101001_110_1_010110101001;
      patterns[44367] = 29'b1_010110101001_111_1_010110101001;
      patterns[44368] = 29'b1_010110101010_000_1_010110101010;
      patterns[44369] = 29'b1_010110101010_001_1_101010010110;
      patterns[44370] = 29'b1_010110101010_010_0_101101010101;
      patterns[44371] = 29'b1_010110101010_011_1_011010101010;
      patterns[44372] = 29'b1_010110101010_100_0_101011010101;
      patterns[44373] = 29'b1_010110101010_101_1_010101101010;
      patterns[44374] = 29'b1_010110101010_110_1_010110101010;
      patterns[44375] = 29'b1_010110101010_111_1_010110101010;
      patterns[44376] = 29'b1_010110101011_000_1_010110101011;
      patterns[44377] = 29'b1_010110101011_001_1_101011010110;
      patterns[44378] = 29'b1_010110101011_010_0_101101010111;
      patterns[44379] = 29'b1_010110101011_011_1_011010101110;
      patterns[44380] = 29'b1_010110101011_100_1_101011010101;
      patterns[44381] = 29'b1_010110101011_101_1_110101101010;
      patterns[44382] = 29'b1_010110101011_110_1_010110101011;
      patterns[44383] = 29'b1_010110101011_111_1_010110101011;
      patterns[44384] = 29'b1_010110101100_000_1_010110101100;
      patterns[44385] = 29'b1_010110101100_001_1_101100010110;
      patterns[44386] = 29'b1_010110101100_010_0_101101011001;
      patterns[44387] = 29'b1_010110101100_011_1_011010110010;
      patterns[44388] = 29'b1_010110101100_100_0_101011010110;
      patterns[44389] = 29'b1_010110101100_101_0_010101101011;
      patterns[44390] = 29'b1_010110101100_110_1_010110101100;
      patterns[44391] = 29'b1_010110101100_111_1_010110101100;
      patterns[44392] = 29'b1_010110101101_000_1_010110101101;
      patterns[44393] = 29'b1_010110101101_001_1_101101010110;
      patterns[44394] = 29'b1_010110101101_010_0_101101011011;
      patterns[44395] = 29'b1_010110101101_011_1_011010110110;
      patterns[44396] = 29'b1_010110101101_100_1_101011010110;
      patterns[44397] = 29'b1_010110101101_101_0_110101101011;
      patterns[44398] = 29'b1_010110101101_110_1_010110101101;
      patterns[44399] = 29'b1_010110101101_111_1_010110101101;
      patterns[44400] = 29'b1_010110101110_000_1_010110101110;
      patterns[44401] = 29'b1_010110101110_001_1_101110010110;
      patterns[44402] = 29'b1_010110101110_010_0_101101011101;
      patterns[44403] = 29'b1_010110101110_011_1_011010111010;
      patterns[44404] = 29'b1_010110101110_100_0_101011010111;
      patterns[44405] = 29'b1_010110101110_101_1_010101101011;
      patterns[44406] = 29'b1_010110101110_110_1_010110101110;
      patterns[44407] = 29'b1_010110101110_111_1_010110101110;
      patterns[44408] = 29'b1_010110101111_000_1_010110101111;
      patterns[44409] = 29'b1_010110101111_001_1_101111010110;
      patterns[44410] = 29'b1_010110101111_010_0_101101011111;
      patterns[44411] = 29'b1_010110101111_011_1_011010111110;
      patterns[44412] = 29'b1_010110101111_100_1_101011010111;
      patterns[44413] = 29'b1_010110101111_101_1_110101101011;
      patterns[44414] = 29'b1_010110101111_110_1_010110101111;
      patterns[44415] = 29'b1_010110101111_111_1_010110101111;
      patterns[44416] = 29'b1_010110110000_000_1_010110110000;
      patterns[44417] = 29'b1_010110110000_001_1_110000010110;
      patterns[44418] = 29'b1_010110110000_010_0_101101100001;
      patterns[44419] = 29'b1_010110110000_011_1_011011000010;
      patterns[44420] = 29'b1_010110110000_100_0_101011011000;
      patterns[44421] = 29'b1_010110110000_101_0_010101101100;
      patterns[44422] = 29'b1_010110110000_110_1_010110110000;
      patterns[44423] = 29'b1_010110110000_111_1_010110110000;
      patterns[44424] = 29'b1_010110110001_000_1_010110110001;
      patterns[44425] = 29'b1_010110110001_001_1_110001010110;
      patterns[44426] = 29'b1_010110110001_010_0_101101100011;
      patterns[44427] = 29'b1_010110110001_011_1_011011000110;
      patterns[44428] = 29'b1_010110110001_100_1_101011011000;
      patterns[44429] = 29'b1_010110110001_101_0_110101101100;
      patterns[44430] = 29'b1_010110110001_110_1_010110110001;
      patterns[44431] = 29'b1_010110110001_111_1_010110110001;
      patterns[44432] = 29'b1_010110110010_000_1_010110110010;
      patterns[44433] = 29'b1_010110110010_001_1_110010010110;
      patterns[44434] = 29'b1_010110110010_010_0_101101100101;
      patterns[44435] = 29'b1_010110110010_011_1_011011001010;
      patterns[44436] = 29'b1_010110110010_100_0_101011011001;
      patterns[44437] = 29'b1_010110110010_101_1_010101101100;
      patterns[44438] = 29'b1_010110110010_110_1_010110110010;
      patterns[44439] = 29'b1_010110110010_111_1_010110110010;
      patterns[44440] = 29'b1_010110110011_000_1_010110110011;
      patterns[44441] = 29'b1_010110110011_001_1_110011010110;
      patterns[44442] = 29'b1_010110110011_010_0_101101100111;
      patterns[44443] = 29'b1_010110110011_011_1_011011001110;
      patterns[44444] = 29'b1_010110110011_100_1_101011011001;
      patterns[44445] = 29'b1_010110110011_101_1_110101101100;
      patterns[44446] = 29'b1_010110110011_110_1_010110110011;
      patterns[44447] = 29'b1_010110110011_111_1_010110110011;
      patterns[44448] = 29'b1_010110110100_000_1_010110110100;
      patterns[44449] = 29'b1_010110110100_001_1_110100010110;
      patterns[44450] = 29'b1_010110110100_010_0_101101101001;
      patterns[44451] = 29'b1_010110110100_011_1_011011010010;
      patterns[44452] = 29'b1_010110110100_100_0_101011011010;
      patterns[44453] = 29'b1_010110110100_101_0_010101101101;
      patterns[44454] = 29'b1_010110110100_110_1_010110110100;
      patterns[44455] = 29'b1_010110110100_111_1_010110110100;
      patterns[44456] = 29'b1_010110110101_000_1_010110110101;
      patterns[44457] = 29'b1_010110110101_001_1_110101010110;
      patterns[44458] = 29'b1_010110110101_010_0_101101101011;
      patterns[44459] = 29'b1_010110110101_011_1_011011010110;
      patterns[44460] = 29'b1_010110110101_100_1_101011011010;
      patterns[44461] = 29'b1_010110110101_101_0_110101101101;
      patterns[44462] = 29'b1_010110110101_110_1_010110110101;
      patterns[44463] = 29'b1_010110110101_111_1_010110110101;
      patterns[44464] = 29'b1_010110110110_000_1_010110110110;
      patterns[44465] = 29'b1_010110110110_001_1_110110010110;
      patterns[44466] = 29'b1_010110110110_010_0_101101101101;
      patterns[44467] = 29'b1_010110110110_011_1_011011011010;
      patterns[44468] = 29'b1_010110110110_100_0_101011011011;
      patterns[44469] = 29'b1_010110110110_101_1_010101101101;
      patterns[44470] = 29'b1_010110110110_110_1_010110110110;
      patterns[44471] = 29'b1_010110110110_111_1_010110110110;
      patterns[44472] = 29'b1_010110110111_000_1_010110110111;
      patterns[44473] = 29'b1_010110110111_001_1_110111010110;
      patterns[44474] = 29'b1_010110110111_010_0_101101101111;
      patterns[44475] = 29'b1_010110110111_011_1_011011011110;
      patterns[44476] = 29'b1_010110110111_100_1_101011011011;
      patterns[44477] = 29'b1_010110110111_101_1_110101101101;
      patterns[44478] = 29'b1_010110110111_110_1_010110110111;
      patterns[44479] = 29'b1_010110110111_111_1_010110110111;
      patterns[44480] = 29'b1_010110111000_000_1_010110111000;
      patterns[44481] = 29'b1_010110111000_001_1_111000010110;
      patterns[44482] = 29'b1_010110111000_010_0_101101110001;
      patterns[44483] = 29'b1_010110111000_011_1_011011100010;
      patterns[44484] = 29'b1_010110111000_100_0_101011011100;
      patterns[44485] = 29'b1_010110111000_101_0_010101101110;
      patterns[44486] = 29'b1_010110111000_110_1_010110111000;
      patterns[44487] = 29'b1_010110111000_111_1_010110111000;
      patterns[44488] = 29'b1_010110111001_000_1_010110111001;
      patterns[44489] = 29'b1_010110111001_001_1_111001010110;
      patterns[44490] = 29'b1_010110111001_010_0_101101110011;
      patterns[44491] = 29'b1_010110111001_011_1_011011100110;
      patterns[44492] = 29'b1_010110111001_100_1_101011011100;
      patterns[44493] = 29'b1_010110111001_101_0_110101101110;
      patterns[44494] = 29'b1_010110111001_110_1_010110111001;
      patterns[44495] = 29'b1_010110111001_111_1_010110111001;
      patterns[44496] = 29'b1_010110111010_000_1_010110111010;
      patterns[44497] = 29'b1_010110111010_001_1_111010010110;
      patterns[44498] = 29'b1_010110111010_010_0_101101110101;
      patterns[44499] = 29'b1_010110111010_011_1_011011101010;
      patterns[44500] = 29'b1_010110111010_100_0_101011011101;
      patterns[44501] = 29'b1_010110111010_101_1_010101101110;
      patterns[44502] = 29'b1_010110111010_110_1_010110111010;
      patterns[44503] = 29'b1_010110111010_111_1_010110111010;
      patterns[44504] = 29'b1_010110111011_000_1_010110111011;
      patterns[44505] = 29'b1_010110111011_001_1_111011010110;
      patterns[44506] = 29'b1_010110111011_010_0_101101110111;
      patterns[44507] = 29'b1_010110111011_011_1_011011101110;
      patterns[44508] = 29'b1_010110111011_100_1_101011011101;
      patterns[44509] = 29'b1_010110111011_101_1_110101101110;
      patterns[44510] = 29'b1_010110111011_110_1_010110111011;
      patterns[44511] = 29'b1_010110111011_111_1_010110111011;
      patterns[44512] = 29'b1_010110111100_000_1_010110111100;
      patterns[44513] = 29'b1_010110111100_001_1_111100010110;
      patterns[44514] = 29'b1_010110111100_010_0_101101111001;
      patterns[44515] = 29'b1_010110111100_011_1_011011110010;
      patterns[44516] = 29'b1_010110111100_100_0_101011011110;
      patterns[44517] = 29'b1_010110111100_101_0_010101101111;
      patterns[44518] = 29'b1_010110111100_110_1_010110111100;
      patterns[44519] = 29'b1_010110111100_111_1_010110111100;
      patterns[44520] = 29'b1_010110111101_000_1_010110111101;
      patterns[44521] = 29'b1_010110111101_001_1_111101010110;
      patterns[44522] = 29'b1_010110111101_010_0_101101111011;
      patterns[44523] = 29'b1_010110111101_011_1_011011110110;
      patterns[44524] = 29'b1_010110111101_100_1_101011011110;
      patterns[44525] = 29'b1_010110111101_101_0_110101101111;
      patterns[44526] = 29'b1_010110111101_110_1_010110111101;
      patterns[44527] = 29'b1_010110111101_111_1_010110111101;
      patterns[44528] = 29'b1_010110111110_000_1_010110111110;
      patterns[44529] = 29'b1_010110111110_001_1_111110010110;
      patterns[44530] = 29'b1_010110111110_010_0_101101111101;
      patterns[44531] = 29'b1_010110111110_011_1_011011111010;
      patterns[44532] = 29'b1_010110111110_100_0_101011011111;
      patterns[44533] = 29'b1_010110111110_101_1_010101101111;
      patterns[44534] = 29'b1_010110111110_110_1_010110111110;
      patterns[44535] = 29'b1_010110111110_111_1_010110111110;
      patterns[44536] = 29'b1_010110111111_000_1_010110111111;
      patterns[44537] = 29'b1_010110111111_001_1_111111010110;
      patterns[44538] = 29'b1_010110111111_010_0_101101111111;
      patterns[44539] = 29'b1_010110111111_011_1_011011111110;
      patterns[44540] = 29'b1_010110111111_100_1_101011011111;
      patterns[44541] = 29'b1_010110111111_101_1_110101101111;
      patterns[44542] = 29'b1_010110111111_110_1_010110111111;
      patterns[44543] = 29'b1_010110111111_111_1_010110111111;
      patterns[44544] = 29'b1_010111000000_000_1_010111000000;
      patterns[44545] = 29'b1_010111000000_001_1_000000010111;
      patterns[44546] = 29'b1_010111000000_010_0_101110000001;
      patterns[44547] = 29'b1_010111000000_011_1_011100000010;
      patterns[44548] = 29'b1_010111000000_100_0_101011100000;
      patterns[44549] = 29'b1_010111000000_101_0_010101110000;
      patterns[44550] = 29'b1_010111000000_110_1_010111000000;
      patterns[44551] = 29'b1_010111000000_111_1_010111000000;
      patterns[44552] = 29'b1_010111000001_000_1_010111000001;
      patterns[44553] = 29'b1_010111000001_001_1_000001010111;
      patterns[44554] = 29'b1_010111000001_010_0_101110000011;
      patterns[44555] = 29'b1_010111000001_011_1_011100000110;
      patterns[44556] = 29'b1_010111000001_100_1_101011100000;
      patterns[44557] = 29'b1_010111000001_101_0_110101110000;
      patterns[44558] = 29'b1_010111000001_110_1_010111000001;
      patterns[44559] = 29'b1_010111000001_111_1_010111000001;
      patterns[44560] = 29'b1_010111000010_000_1_010111000010;
      patterns[44561] = 29'b1_010111000010_001_1_000010010111;
      patterns[44562] = 29'b1_010111000010_010_0_101110000101;
      patterns[44563] = 29'b1_010111000010_011_1_011100001010;
      patterns[44564] = 29'b1_010111000010_100_0_101011100001;
      patterns[44565] = 29'b1_010111000010_101_1_010101110000;
      patterns[44566] = 29'b1_010111000010_110_1_010111000010;
      patterns[44567] = 29'b1_010111000010_111_1_010111000010;
      patterns[44568] = 29'b1_010111000011_000_1_010111000011;
      patterns[44569] = 29'b1_010111000011_001_1_000011010111;
      patterns[44570] = 29'b1_010111000011_010_0_101110000111;
      patterns[44571] = 29'b1_010111000011_011_1_011100001110;
      patterns[44572] = 29'b1_010111000011_100_1_101011100001;
      patterns[44573] = 29'b1_010111000011_101_1_110101110000;
      patterns[44574] = 29'b1_010111000011_110_1_010111000011;
      patterns[44575] = 29'b1_010111000011_111_1_010111000011;
      patterns[44576] = 29'b1_010111000100_000_1_010111000100;
      patterns[44577] = 29'b1_010111000100_001_1_000100010111;
      patterns[44578] = 29'b1_010111000100_010_0_101110001001;
      patterns[44579] = 29'b1_010111000100_011_1_011100010010;
      patterns[44580] = 29'b1_010111000100_100_0_101011100010;
      patterns[44581] = 29'b1_010111000100_101_0_010101110001;
      patterns[44582] = 29'b1_010111000100_110_1_010111000100;
      patterns[44583] = 29'b1_010111000100_111_1_010111000100;
      patterns[44584] = 29'b1_010111000101_000_1_010111000101;
      patterns[44585] = 29'b1_010111000101_001_1_000101010111;
      patterns[44586] = 29'b1_010111000101_010_0_101110001011;
      patterns[44587] = 29'b1_010111000101_011_1_011100010110;
      patterns[44588] = 29'b1_010111000101_100_1_101011100010;
      patterns[44589] = 29'b1_010111000101_101_0_110101110001;
      patterns[44590] = 29'b1_010111000101_110_1_010111000101;
      patterns[44591] = 29'b1_010111000101_111_1_010111000101;
      patterns[44592] = 29'b1_010111000110_000_1_010111000110;
      patterns[44593] = 29'b1_010111000110_001_1_000110010111;
      patterns[44594] = 29'b1_010111000110_010_0_101110001101;
      patterns[44595] = 29'b1_010111000110_011_1_011100011010;
      patterns[44596] = 29'b1_010111000110_100_0_101011100011;
      patterns[44597] = 29'b1_010111000110_101_1_010101110001;
      patterns[44598] = 29'b1_010111000110_110_1_010111000110;
      patterns[44599] = 29'b1_010111000110_111_1_010111000110;
      patterns[44600] = 29'b1_010111000111_000_1_010111000111;
      patterns[44601] = 29'b1_010111000111_001_1_000111010111;
      patterns[44602] = 29'b1_010111000111_010_0_101110001111;
      patterns[44603] = 29'b1_010111000111_011_1_011100011110;
      patterns[44604] = 29'b1_010111000111_100_1_101011100011;
      patterns[44605] = 29'b1_010111000111_101_1_110101110001;
      patterns[44606] = 29'b1_010111000111_110_1_010111000111;
      patterns[44607] = 29'b1_010111000111_111_1_010111000111;
      patterns[44608] = 29'b1_010111001000_000_1_010111001000;
      patterns[44609] = 29'b1_010111001000_001_1_001000010111;
      patterns[44610] = 29'b1_010111001000_010_0_101110010001;
      patterns[44611] = 29'b1_010111001000_011_1_011100100010;
      patterns[44612] = 29'b1_010111001000_100_0_101011100100;
      patterns[44613] = 29'b1_010111001000_101_0_010101110010;
      patterns[44614] = 29'b1_010111001000_110_1_010111001000;
      patterns[44615] = 29'b1_010111001000_111_1_010111001000;
      patterns[44616] = 29'b1_010111001001_000_1_010111001001;
      patterns[44617] = 29'b1_010111001001_001_1_001001010111;
      patterns[44618] = 29'b1_010111001001_010_0_101110010011;
      patterns[44619] = 29'b1_010111001001_011_1_011100100110;
      patterns[44620] = 29'b1_010111001001_100_1_101011100100;
      patterns[44621] = 29'b1_010111001001_101_0_110101110010;
      patterns[44622] = 29'b1_010111001001_110_1_010111001001;
      patterns[44623] = 29'b1_010111001001_111_1_010111001001;
      patterns[44624] = 29'b1_010111001010_000_1_010111001010;
      patterns[44625] = 29'b1_010111001010_001_1_001010010111;
      patterns[44626] = 29'b1_010111001010_010_0_101110010101;
      patterns[44627] = 29'b1_010111001010_011_1_011100101010;
      patterns[44628] = 29'b1_010111001010_100_0_101011100101;
      patterns[44629] = 29'b1_010111001010_101_1_010101110010;
      patterns[44630] = 29'b1_010111001010_110_1_010111001010;
      patterns[44631] = 29'b1_010111001010_111_1_010111001010;
      patterns[44632] = 29'b1_010111001011_000_1_010111001011;
      patterns[44633] = 29'b1_010111001011_001_1_001011010111;
      patterns[44634] = 29'b1_010111001011_010_0_101110010111;
      patterns[44635] = 29'b1_010111001011_011_1_011100101110;
      patterns[44636] = 29'b1_010111001011_100_1_101011100101;
      patterns[44637] = 29'b1_010111001011_101_1_110101110010;
      patterns[44638] = 29'b1_010111001011_110_1_010111001011;
      patterns[44639] = 29'b1_010111001011_111_1_010111001011;
      patterns[44640] = 29'b1_010111001100_000_1_010111001100;
      patterns[44641] = 29'b1_010111001100_001_1_001100010111;
      patterns[44642] = 29'b1_010111001100_010_0_101110011001;
      patterns[44643] = 29'b1_010111001100_011_1_011100110010;
      patterns[44644] = 29'b1_010111001100_100_0_101011100110;
      patterns[44645] = 29'b1_010111001100_101_0_010101110011;
      patterns[44646] = 29'b1_010111001100_110_1_010111001100;
      patterns[44647] = 29'b1_010111001100_111_1_010111001100;
      patterns[44648] = 29'b1_010111001101_000_1_010111001101;
      patterns[44649] = 29'b1_010111001101_001_1_001101010111;
      patterns[44650] = 29'b1_010111001101_010_0_101110011011;
      patterns[44651] = 29'b1_010111001101_011_1_011100110110;
      patterns[44652] = 29'b1_010111001101_100_1_101011100110;
      patterns[44653] = 29'b1_010111001101_101_0_110101110011;
      patterns[44654] = 29'b1_010111001101_110_1_010111001101;
      patterns[44655] = 29'b1_010111001101_111_1_010111001101;
      patterns[44656] = 29'b1_010111001110_000_1_010111001110;
      patterns[44657] = 29'b1_010111001110_001_1_001110010111;
      patterns[44658] = 29'b1_010111001110_010_0_101110011101;
      patterns[44659] = 29'b1_010111001110_011_1_011100111010;
      patterns[44660] = 29'b1_010111001110_100_0_101011100111;
      patterns[44661] = 29'b1_010111001110_101_1_010101110011;
      patterns[44662] = 29'b1_010111001110_110_1_010111001110;
      patterns[44663] = 29'b1_010111001110_111_1_010111001110;
      patterns[44664] = 29'b1_010111001111_000_1_010111001111;
      patterns[44665] = 29'b1_010111001111_001_1_001111010111;
      patterns[44666] = 29'b1_010111001111_010_0_101110011111;
      patterns[44667] = 29'b1_010111001111_011_1_011100111110;
      patterns[44668] = 29'b1_010111001111_100_1_101011100111;
      patterns[44669] = 29'b1_010111001111_101_1_110101110011;
      patterns[44670] = 29'b1_010111001111_110_1_010111001111;
      patterns[44671] = 29'b1_010111001111_111_1_010111001111;
      patterns[44672] = 29'b1_010111010000_000_1_010111010000;
      patterns[44673] = 29'b1_010111010000_001_1_010000010111;
      patterns[44674] = 29'b1_010111010000_010_0_101110100001;
      patterns[44675] = 29'b1_010111010000_011_1_011101000010;
      patterns[44676] = 29'b1_010111010000_100_0_101011101000;
      patterns[44677] = 29'b1_010111010000_101_0_010101110100;
      patterns[44678] = 29'b1_010111010000_110_1_010111010000;
      patterns[44679] = 29'b1_010111010000_111_1_010111010000;
      patterns[44680] = 29'b1_010111010001_000_1_010111010001;
      patterns[44681] = 29'b1_010111010001_001_1_010001010111;
      patterns[44682] = 29'b1_010111010001_010_0_101110100011;
      patterns[44683] = 29'b1_010111010001_011_1_011101000110;
      patterns[44684] = 29'b1_010111010001_100_1_101011101000;
      patterns[44685] = 29'b1_010111010001_101_0_110101110100;
      patterns[44686] = 29'b1_010111010001_110_1_010111010001;
      patterns[44687] = 29'b1_010111010001_111_1_010111010001;
      patterns[44688] = 29'b1_010111010010_000_1_010111010010;
      patterns[44689] = 29'b1_010111010010_001_1_010010010111;
      patterns[44690] = 29'b1_010111010010_010_0_101110100101;
      patterns[44691] = 29'b1_010111010010_011_1_011101001010;
      patterns[44692] = 29'b1_010111010010_100_0_101011101001;
      patterns[44693] = 29'b1_010111010010_101_1_010101110100;
      patterns[44694] = 29'b1_010111010010_110_1_010111010010;
      patterns[44695] = 29'b1_010111010010_111_1_010111010010;
      patterns[44696] = 29'b1_010111010011_000_1_010111010011;
      patterns[44697] = 29'b1_010111010011_001_1_010011010111;
      patterns[44698] = 29'b1_010111010011_010_0_101110100111;
      patterns[44699] = 29'b1_010111010011_011_1_011101001110;
      patterns[44700] = 29'b1_010111010011_100_1_101011101001;
      patterns[44701] = 29'b1_010111010011_101_1_110101110100;
      patterns[44702] = 29'b1_010111010011_110_1_010111010011;
      patterns[44703] = 29'b1_010111010011_111_1_010111010011;
      patterns[44704] = 29'b1_010111010100_000_1_010111010100;
      patterns[44705] = 29'b1_010111010100_001_1_010100010111;
      patterns[44706] = 29'b1_010111010100_010_0_101110101001;
      patterns[44707] = 29'b1_010111010100_011_1_011101010010;
      patterns[44708] = 29'b1_010111010100_100_0_101011101010;
      patterns[44709] = 29'b1_010111010100_101_0_010101110101;
      patterns[44710] = 29'b1_010111010100_110_1_010111010100;
      patterns[44711] = 29'b1_010111010100_111_1_010111010100;
      patterns[44712] = 29'b1_010111010101_000_1_010111010101;
      patterns[44713] = 29'b1_010111010101_001_1_010101010111;
      patterns[44714] = 29'b1_010111010101_010_0_101110101011;
      patterns[44715] = 29'b1_010111010101_011_1_011101010110;
      patterns[44716] = 29'b1_010111010101_100_1_101011101010;
      patterns[44717] = 29'b1_010111010101_101_0_110101110101;
      patterns[44718] = 29'b1_010111010101_110_1_010111010101;
      patterns[44719] = 29'b1_010111010101_111_1_010111010101;
      patterns[44720] = 29'b1_010111010110_000_1_010111010110;
      patterns[44721] = 29'b1_010111010110_001_1_010110010111;
      patterns[44722] = 29'b1_010111010110_010_0_101110101101;
      patterns[44723] = 29'b1_010111010110_011_1_011101011010;
      patterns[44724] = 29'b1_010111010110_100_0_101011101011;
      patterns[44725] = 29'b1_010111010110_101_1_010101110101;
      patterns[44726] = 29'b1_010111010110_110_1_010111010110;
      patterns[44727] = 29'b1_010111010110_111_1_010111010110;
      patterns[44728] = 29'b1_010111010111_000_1_010111010111;
      patterns[44729] = 29'b1_010111010111_001_1_010111010111;
      patterns[44730] = 29'b1_010111010111_010_0_101110101111;
      patterns[44731] = 29'b1_010111010111_011_1_011101011110;
      patterns[44732] = 29'b1_010111010111_100_1_101011101011;
      patterns[44733] = 29'b1_010111010111_101_1_110101110101;
      patterns[44734] = 29'b1_010111010111_110_1_010111010111;
      patterns[44735] = 29'b1_010111010111_111_1_010111010111;
      patterns[44736] = 29'b1_010111011000_000_1_010111011000;
      patterns[44737] = 29'b1_010111011000_001_1_011000010111;
      patterns[44738] = 29'b1_010111011000_010_0_101110110001;
      patterns[44739] = 29'b1_010111011000_011_1_011101100010;
      patterns[44740] = 29'b1_010111011000_100_0_101011101100;
      patterns[44741] = 29'b1_010111011000_101_0_010101110110;
      patterns[44742] = 29'b1_010111011000_110_1_010111011000;
      patterns[44743] = 29'b1_010111011000_111_1_010111011000;
      patterns[44744] = 29'b1_010111011001_000_1_010111011001;
      patterns[44745] = 29'b1_010111011001_001_1_011001010111;
      patterns[44746] = 29'b1_010111011001_010_0_101110110011;
      patterns[44747] = 29'b1_010111011001_011_1_011101100110;
      patterns[44748] = 29'b1_010111011001_100_1_101011101100;
      patterns[44749] = 29'b1_010111011001_101_0_110101110110;
      patterns[44750] = 29'b1_010111011001_110_1_010111011001;
      patterns[44751] = 29'b1_010111011001_111_1_010111011001;
      patterns[44752] = 29'b1_010111011010_000_1_010111011010;
      patterns[44753] = 29'b1_010111011010_001_1_011010010111;
      patterns[44754] = 29'b1_010111011010_010_0_101110110101;
      patterns[44755] = 29'b1_010111011010_011_1_011101101010;
      patterns[44756] = 29'b1_010111011010_100_0_101011101101;
      patterns[44757] = 29'b1_010111011010_101_1_010101110110;
      patterns[44758] = 29'b1_010111011010_110_1_010111011010;
      patterns[44759] = 29'b1_010111011010_111_1_010111011010;
      patterns[44760] = 29'b1_010111011011_000_1_010111011011;
      patterns[44761] = 29'b1_010111011011_001_1_011011010111;
      patterns[44762] = 29'b1_010111011011_010_0_101110110111;
      patterns[44763] = 29'b1_010111011011_011_1_011101101110;
      patterns[44764] = 29'b1_010111011011_100_1_101011101101;
      patterns[44765] = 29'b1_010111011011_101_1_110101110110;
      patterns[44766] = 29'b1_010111011011_110_1_010111011011;
      patterns[44767] = 29'b1_010111011011_111_1_010111011011;
      patterns[44768] = 29'b1_010111011100_000_1_010111011100;
      patterns[44769] = 29'b1_010111011100_001_1_011100010111;
      patterns[44770] = 29'b1_010111011100_010_0_101110111001;
      patterns[44771] = 29'b1_010111011100_011_1_011101110010;
      patterns[44772] = 29'b1_010111011100_100_0_101011101110;
      patterns[44773] = 29'b1_010111011100_101_0_010101110111;
      patterns[44774] = 29'b1_010111011100_110_1_010111011100;
      patterns[44775] = 29'b1_010111011100_111_1_010111011100;
      patterns[44776] = 29'b1_010111011101_000_1_010111011101;
      patterns[44777] = 29'b1_010111011101_001_1_011101010111;
      patterns[44778] = 29'b1_010111011101_010_0_101110111011;
      patterns[44779] = 29'b1_010111011101_011_1_011101110110;
      patterns[44780] = 29'b1_010111011101_100_1_101011101110;
      patterns[44781] = 29'b1_010111011101_101_0_110101110111;
      patterns[44782] = 29'b1_010111011101_110_1_010111011101;
      patterns[44783] = 29'b1_010111011101_111_1_010111011101;
      patterns[44784] = 29'b1_010111011110_000_1_010111011110;
      patterns[44785] = 29'b1_010111011110_001_1_011110010111;
      patterns[44786] = 29'b1_010111011110_010_0_101110111101;
      patterns[44787] = 29'b1_010111011110_011_1_011101111010;
      patterns[44788] = 29'b1_010111011110_100_0_101011101111;
      patterns[44789] = 29'b1_010111011110_101_1_010101110111;
      patterns[44790] = 29'b1_010111011110_110_1_010111011110;
      patterns[44791] = 29'b1_010111011110_111_1_010111011110;
      patterns[44792] = 29'b1_010111011111_000_1_010111011111;
      patterns[44793] = 29'b1_010111011111_001_1_011111010111;
      patterns[44794] = 29'b1_010111011111_010_0_101110111111;
      patterns[44795] = 29'b1_010111011111_011_1_011101111110;
      patterns[44796] = 29'b1_010111011111_100_1_101011101111;
      patterns[44797] = 29'b1_010111011111_101_1_110101110111;
      patterns[44798] = 29'b1_010111011111_110_1_010111011111;
      patterns[44799] = 29'b1_010111011111_111_1_010111011111;
      patterns[44800] = 29'b1_010111100000_000_1_010111100000;
      patterns[44801] = 29'b1_010111100000_001_1_100000010111;
      patterns[44802] = 29'b1_010111100000_010_0_101111000001;
      patterns[44803] = 29'b1_010111100000_011_1_011110000010;
      patterns[44804] = 29'b1_010111100000_100_0_101011110000;
      patterns[44805] = 29'b1_010111100000_101_0_010101111000;
      patterns[44806] = 29'b1_010111100000_110_1_010111100000;
      patterns[44807] = 29'b1_010111100000_111_1_010111100000;
      patterns[44808] = 29'b1_010111100001_000_1_010111100001;
      patterns[44809] = 29'b1_010111100001_001_1_100001010111;
      patterns[44810] = 29'b1_010111100001_010_0_101111000011;
      patterns[44811] = 29'b1_010111100001_011_1_011110000110;
      patterns[44812] = 29'b1_010111100001_100_1_101011110000;
      patterns[44813] = 29'b1_010111100001_101_0_110101111000;
      patterns[44814] = 29'b1_010111100001_110_1_010111100001;
      patterns[44815] = 29'b1_010111100001_111_1_010111100001;
      patterns[44816] = 29'b1_010111100010_000_1_010111100010;
      patterns[44817] = 29'b1_010111100010_001_1_100010010111;
      patterns[44818] = 29'b1_010111100010_010_0_101111000101;
      patterns[44819] = 29'b1_010111100010_011_1_011110001010;
      patterns[44820] = 29'b1_010111100010_100_0_101011110001;
      patterns[44821] = 29'b1_010111100010_101_1_010101111000;
      patterns[44822] = 29'b1_010111100010_110_1_010111100010;
      patterns[44823] = 29'b1_010111100010_111_1_010111100010;
      patterns[44824] = 29'b1_010111100011_000_1_010111100011;
      patterns[44825] = 29'b1_010111100011_001_1_100011010111;
      patterns[44826] = 29'b1_010111100011_010_0_101111000111;
      patterns[44827] = 29'b1_010111100011_011_1_011110001110;
      patterns[44828] = 29'b1_010111100011_100_1_101011110001;
      patterns[44829] = 29'b1_010111100011_101_1_110101111000;
      patterns[44830] = 29'b1_010111100011_110_1_010111100011;
      patterns[44831] = 29'b1_010111100011_111_1_010111100011;
      patterns[44832] = 29'b1_010111100100_000_1_010111100100;
      patterns[44833] = 29'b1_010111100100_001_1_100100010111;
      patterns[44834] = 29'b1_010111100100_010_0_101111001001;
      patterns[44835] = 29'b1_010111100100_011_1_011110010010;
      patterns[44836] = 29'b1_010111100100_100_0_101011110010;
      patterns[44837] = 29'b1_010111100100_101_0_010101111001;
      patterns[44838] = 29'b1_010111100100_110_1_010111100100;
      patterns[44839] = 29'b1_010111100100_111_1_010111100100;
      patterns[44840] = 29'b1_010111100101_000_1_010111100101;
      patterns[44841] = 29'b1_010111100101_001_1_100101010111;
      patterns[44842] = 29'b1_010111100101_010_0_101111001011;
      patterns[44843] = 29'b1_010111100101_011_1_011110010110;
      patterns[44844] = 29'b1_010111100101_100_1_101011110010;
      patterns[44845] = 29'b1_010111100101_101_0_110101111001;
      patterns[44846] = 29'b1_010111100101_110_1_010111100101;
      patterns[44847] = 29'b1_010111100101_111_1_010111100101;
      patterns[44848] = 29'b1_010111100110_000_1_010111100110;
      patterns[44849] = 29'b1_010111100110_001_1_100110010111;
      patterns[44850] = 29'b1_010111100110_010_0_101111001101;
      patterns[44851] = 29'b1_010111100110_011_1_011110011010;
      patterns[44852] = 29'b1_010111100110_100_0_101011110011;
      patterns[44853] = 29'b1_010111100110_101_1_010101111001;
      patterns[44854] = 29'b1_010111100110_110_1_010111100110;
      patterns[44855] = 29'b1_010111100110_111_1_010111100110;
      patterns[44856] = 29'b1_010111100111_000_1_010111100111;
      patterns[44857] = 29'b1_010111100111_001_1_100111010111;
      patterns[44858] = 29'b1_010111100111_010_0_101111001111;
      patterns[44859] = 29'b1_010111100111_011_1_011110011110;
      patterns[44860] = 29'b1_010111100111_100_1_101011110011;
      patterns[44861] = 29'b1_010111100111_101_1_110101111001;
      patterns[44862] = 29'b1_010111100111_110_1_010111100111;
      patterns[44863] = 29'b1_010111100111_111_1_010111100111;
      patterns[44864] = 29'b1_010111101000_000_1_010111101000;
      patterns[44865] = 29'b1_010111101000_001_1_101000010111;
      patterns[44866] = 29'b1_010111101000_010_0_101111010001;
      patterns[44867] = 29'b1_010111101000_011_1_011110100010;
      patterns[44868] = 29'b1_010111101000_100_0_101011110100;
      patterns[44869] = 29'b1_010111101000_101_0_010101111010;
      patterns[44870] = 29'b1_010111101000_110_1_010111101000;
      patterns[44871] = 29'b1_010111101000_111_1_010111101000;
      patterns[44872] = 29'b1_010111101001_000_1_010111101001;
      patterns[44873] = 29'b1_010111101001_001_1_101001010111;
      patterns[44874] = 29'b1_010111101001_010_0_101111010011;
      patterns[44875] = 29'b1_010111101001_011_1_011110100110;
      patterns[44876] = 29'b1_010111101001_100_1_101011110100;
      patterns[44877] = 29'b1_010111101001_101_0_110101111010;
      patterns[44878] = 29'b1_010111101001_110_1_010111101001;
      patterns[44879] = 29'b1_010111101001_111_1_010111101001;
      patterns[44880] = 29'b1_010111101010_000_1_010111101010;
      patterns[44881] = 29'b1_010111101010_001_1_101010010111;
      patterns[44882] = 29'b1_010111101010_010_0_101111010101;
      patterns[44883] = 29'b1_010111101010_011_1_011110101010;
      patterns[44884] = 29'b1_010111101010_100_0_101011110101;
      patterns[44885] = 29'b1_010111101010_101_1_010101111010;
      patterns[44886] = 29'b1_010111101010_110_1_010111101010;
      patterns[44887] = 29'b1_010111101010_111_1_010111101010;
      patterns[44888] = 29'b1_010111101011_000_1_010111101011;
      patterns[44889] = 29'b1_010111101011_001_1_101011010111;
      patterns[44890] = 29'b1_010111101011_010_0_101111010111;
      patterns[44891] = 29'b1_010111101011_011_1_011110101110;
      patterns[44892] = 29'b1_010111101011_100_1_101011110101;
      patterns[44893] = 29'b1_010111101011_101_1_110101111010;
      patterns[44894] = 29'b1_010111101011_110_1_010111101011;
      patterns[44895] = 29'b1_010111101011_111_1_010111101011;
      patterns[44896] = 29'b1_010111101100_000_1_010111101100;
      patterns[44897] = 29'b1_010111101100_001_1_101100010111;
      patterns[44898] = 29'b1_010111101100_010_0_101111011001;
      patterns[44899] = 29'b1_010111101100_011_1_011110110010;
      patterns[44900] = 29'b1_010111101100_100_0_101011110110;
      patterns[44901] = 29'b1_010111101100_101_0_010101111011;
      patterns[44902] = 29'b1_010111101100_110_1_010111101100;
      patterns[44903] = 29'b1_010111101100_111_1_010111101100;
      patterns[44904] = 29'b1_010111101101_000_1_010111101101;
      patterns[44905] = 29'b1_010111101101_001_1_101101010111;
      patterns[44906] = 29'b1_010111101101_010_0_101111011011;
      patterns[44907] = 29'b1_010111101101_011_1_011110110110;
      patterns[44908] = 29'b1_010111101101_100_1_101011110110;
      patterns[44909] = 29'b1_010111101101_101_0_110101111011;
      patterns[44910] = 29'b1_010111101101_110_1_010111101101;
      patterns[44911] = 29'b1_010111101101_111_1_010111101101;
      patterns[44912] = 29'b1_010111101110_000_1_010111101110;
      patterns[44913] = 29'b1_010111101110_001_1_101110010111;
      patterns[44914] = 29'b1_010111101110_010_0_101111011101;
      patterns[44915] = 29'b1_010111101110_011_1_011110111010;
      patterns[44916] = 29'b1_010111101110_100_0_101011110111;
      patterns[44917] = 29'b1_010111101110_101_1_010101111011;
      patterns[44918] = 29'b1_010111101110_110_1_010111101110;
      patterns[44919] = 29'b1_010111101110_111_1_010111101110;
      patterns[44920] = 29'b1_010111101111_000_1_010111101111;
      patterns[44921] = 29'b1_010111101111_001_1_101111010111;
      patterns[44922] = 29'b1_010111101111_010_0_101111011111;
      patterns[44923] = 29'b1_010111101111_011_1_011110111110;
      patterns[44924] = 29'b1_010111101111_100_1_101011110111;
      patterns[44925] = 29'b1_010111101111_101_1_110101111011;
      patterns[44926] = 29'b1_010111101111_110_1_010111101111;
      patterns[44927] = 29'b1_010111101111_111_1_010111101111;
      patterns[44928] = 29'b1_010111110000_000_1_010111110000;
      patterns[44929] = 29'b1_010111110000_001_1_110000010111;
      patterns[44930] = 29'b1_010111110000_010_0_101111100001;
      patterns[44931] = 29'b1_010111110000_011_1_011111000010;
      patterns[44932] = 29'b1_010111110000_100_0_101011111000;
      patterns[44933] = 29'b1_010111110000_101_0_010101111100;
      patterns[44934] = 29'b1_010111110000_110_1_010111110000;
      patterns[44935] = 29'b1_010111110000_111_1_010111110000;
      patterns[44936] = 29'b1_010111110001_000_1_010111110001;
      patterns[44937] = 29'b1_010111110001_001_1_110001010111;
      patterns[44938] = 29'b1_010111110001_010_0_101111100011;
      patterns[44939] = 29'b1_010111110001_011_1_011111000110;
      patterns[44940] = 29'b1_010111110001_100_1_101011111000;
      patterns[44941] = 29'b1_010111110001_101_0_110101111100;
      patterns[44942] = 29'b1_010111110001_110_1_010111110001;
      patterns[44943] = 29'b1_010111110001_111_1_010111110001;
      patterns[44944] = 29'b1_010111110010_000_1_010111110010;
      patterns[44945] = 29'b1_010111110010_001_1_110010010111;
      patterns[44946] = 29'b1_010111110010_010_0_101111100101;
      patterns[44947] = 29'b1_010111110010_011_1_011111001010;
      patterns[44948] = 29'b1_010111110010_100_0_101011111001;
      patterns[44949] = 29'b1_010111110010_101_1_010101111100;
      patterns[44950] = 29'b1_010111110010_110_1_010111110010;
      patterns[44951] = 29'b1_010111110010_111_1_010111110010;
      patterns[44952] = 29'b1_010111110011_000_1_010111110011;
      patterns[44953] = 29'b1_010111110011_001_1_110011010111;
      patterns[44954] = 29'b1_010111110011_010_0_101111100111;
      patterns[44955] = 29'b1_010111110011_011_1_011111001110;
      patterns[44956] = 29'b1_010111110011_100_1_101011111001;
      patterns[44957] = 29'b1_010111110011_101_1_110101111100;
      patterns[44958] = 29'b1_010111110011_110_1_010111110011;
      patterns[44959] = 29'b1_010111110011_111_1_010111110011;
      patterns[44960] = 29'b1_010111110100_000_1_010111110100;
      patterns[44961] = 29'b1_010111110100_001_1_110100010111;
      patterns[44962] = 29'b1_010111110100_010_0_101111101001;
      patterns[44963] = 29'b1_010111110100_011_1_011111010010;
      patterns[44964] = 29'b1_010111110100_100_0_101011111010;
      patterns[44965] = 29'b1_010111110100_101_0_010101111101;
      patterns[44966] = 29'b1_010111110100_110_1_010111110100;
      patterns[44967] = 29'b1_010111110100_111_1_010111110100;
      patterns[44968] = 29'b1_010111110101_000_1_010111110101;
      patterns[44969] = 29'b1_010111110101_001_1_110101010111;
      patterns[44970] = 29'b1_010111110101_010_0_101111101011;
      patterns[44971] = 29'b1_010111110101_011_1_011111010110;
      patterns[44972] = 29'b1_010111110101_100_1_101011111010;
      patterns[44973] = 29'b1_010111110101_101_0_110101111101;
      patterns[44974] = 29'b1_010111110101_110_1_010111110101;
      patterns[44975] = 29'b1_010111110101_111_1_010111110101;
      patterns[44976] = 29'b1_010111110110_000_1_010111110110;
      patterns[44977] = 29'b1_010111110110_001_1_110110010111;
      patterns[44978] = 29'b1_010111110110_010_0_101111101101;
      patterns[44979] = 29'b1_010111110110_011_1_011111011010;
      patterns[44980] = 29'b1_010111110110_100_0_101011111011;
      patterns[44981] = 29'b1_010111110110_101_1_010101111101;
      patterns[44982] = 29'b1_010111110110_110_1_010111110110;
      patterns[44983] = 29'b1_010111110110_111_1_010111110110;
      patterns[44984] = 29'b1_010111110111_000_1_010111110111;
      patterns[44985] = 29'b1_010111110111_001_1_110111010111;
      patterns[44986] = 29'b1_010111110111_010_0_101111101111;
      patterns[44987] = 29'b1_010111110111_011_1_011111011110;
      patterns[44988] = 29'b1_010111110111_100_1_101011111011;
      patterns[44989] = 29'b1_010111110111_101_1_110101111101;
      patterns[44990] = 29'b1_010111110111_110_1_010111110111;
      patterns[44991] = 29'b1_010111110111_111_1_010111110111;
      patterns[44992] = 29'b1_010111111000_000_1_010111111000;
      patterns[44993] = 29'b1_010111111000_001_1_111000010111;
      patterns[44994] = 29'b1_010111111000_010_0_101111110001;
      patterns[44995] = 29'b1_010111111000_011_1_011111100010;
      patterns[44996] = 29'b1_010111111000_100_0_101011111100;
      patterns[44997] = 29'b1_010111111000_101_0_010101111110;
      patterns[44998] = 29'b1_010111111000_110_1_010111111000;
      patterns[44999] = 29'b1_010111111000_111_1_010111111000;
      patterns[45000] = 29'b1_010111111001_000_1_010111111001;
      patterns[45001] = 29'b1_010111111001_001_1_111001010111;
      patterns[45002] = 29'b1_010111111001_010_0_101111110011;
      patterns[45003] = 29'b1_010111111001_011_1_011111100110;
      patterns[45004] = 29'b1_010111111001_100_1_101011111100;
      patterns[45005] = 29'b1_010111111001_101_0_110101111110;
      patterns[45006] = 29'b1_010111111001_110_1_010111111001;
      patterns[45007] = 29'b1_010111111001_111_1_010111111001;
      patterns[45008] = 29'b1_010111111010_000_1_010111111010;
      patterns[45009] = 29'b1_010111111010_001_1_111010010111;
      patterns[45010] = 29'b1_010111111010_010_0_101111110101;
      patterns[45011] = 29'b1_010111111010_011_1_011111101010;
      patterns[45012] = 29'b1_010111111010_100_0_101011111101;
      patterns[45013] = 29'b1_010111111010_101_1_010101111110;
      patterns[45014] = 29'b1_010111111010_110_1_010111111010;
      patterns[45015] = 29'b1_010111111010_111_1_010111111010;
      patterns[45016] = 29'b1_010111111011_000_1_010111111011;
      patterns[45017] = 29'b1_010111111011_001_1_111011010111;
      patterns[45018] = 29'b1_010111111011_010_0_101111110111;
      patterns[45019] = 29'b1_010111111011_011_1_011111101110;
      patterns[45020] = 29'b1_010111111011_100_1_101011111101;
      patterns[45021] = 29'b1_010111111011_101_1_110101111110;
      patterns[45022] = 29'b1_010111111011_110_1_010111111011;
      patterns[45023] = 29'b1_010111111011_111_1_010111111011;
      patterns[45024] = 29'b1_010111111100_000_1_010111111100;
      patterns[45025] = 29'b1_010111111100_001_1_111100010111;
      patterns[45026] = 29'b1_010111111100_010_0_101111111001;
      patterns[45027] = 29'b1_010111111100_011_1_011111110010;
      patterns[45028] = 29'b1_010111111100_100_0_101011111110;
      patterns[45029] = 29'b1_010111111100_101_0_010101111111;
      patterns[45030] = 29'b1_010111111100_110_1_010111111100;
      patterns[45031] = 29'b1_010111111100_111_1_010111111100;
      patterns[45032] = 29'b1_010111111101_000_1_010111111101;
      patterns[45033] = 29'b1_010111111101_001_1_111101010111;
      patterns[45034] = 29'b1_010111111101_010_0_101111111011;
      patterns[45035] = 29'b1_010111111101_011_1_011111110110;
      patterns[45036] = 29'b1_010111111101_100_1_101011111110;
      patterns[45037] = 29'b1_010111111101_101_0_110101111111;
      patterns[45038] = 29'b1_010111111101_110_1_010111111101;
      patterns[45039] = 29'b1_010111111101_111_1_010111111101;
      patterns[45040] = 29'b1_010111111110_000_1_010111111110;
      patterns[45041] = 29'b1_010111111110_001_1_111110010111;
      patterns[45042] = 29'b1_010111111110_010_0_101111111101;
      patterns[45043] = 29'b1_010111111110_011_1_011111111010;
      patterns[45044] = 29'b1_010111111110_100_0_101011111111;
      patterns[45045] = 29'b1_010111111110_101_1_010101111111;
      patterns[45046] = 29'b1_010111111110_110_1_010111111110;
      patterns[45047] = 29'b1_010111111110_111_1_010111111110;
      patterns[45048] = 29'b1_010111111111_000_1_010111111111;
      patterns[45049] = 29'b1_010111111111_001_1_111111010111;
      patterns[45050] = 29'b1_010111111111_010_0_101111111111;
      patterns[45051] = 29'b1_010111111111_011_1_011111111110;
      patterns[45052] = 29'b1_010111111111_100_1_101011111111;
      patterns[45053] = 29'b1_010111111111_101_1_110101111111;
      patterns[45054] = 29'b1_010111111111_110_1_010111111111;
      patterns[45055] = 29'b1_010111111111_111_1_010111111111;
      patterns[45056] = 29'b1_011000000000_000_1_011000000000;
      patterns[45057] = 29'b1_011000000000_001_1_000000011000;
      patterns[45058] = 29'b1_011000000000_010_0_110000000001;
      patterns[45059] = 29'b1_011000000000_011_1_100000000010;
      patterns[45060] = 29'b1_011000000000_100_0_101100000000;
      patterns[45061] = 29'b1_011000000000_101_0_010110000000;
      patterns[45062] = 29'b1_011000000000_110_1_011000000000;
      patterns[45063] = 29'b1_011000000000_111_1_011000000000;
      patterns[45064] = 29'b1_011000000001_000_1_011000000001;
      patterns[45065] = 29'b1_011000000001_001_1_000001011000;
      patterns[45066] = 29'b1_011000000001_010_0_110000000011;
      patterns[45067] = 29'b1_011000000001_011_1_100000000110;
      patterns[45068] = 29'b1_011000000001_100_1_101100000000;
      patterns[45069] = 29'b1_011000000001_101_0_110110000000;
      patterns[45070] = 29'b1_011000000001_110_1_011000000001;
      patterns[45071] = 29'b1_011000000001_111_1_011000000001;
      patterns[45072] = 29'b1_011000000010_000_1_011000000010;
      patterns[45073] = 29'b1_011000000010_001_1_000010011000;
      patterns[45074] = 29'b1_011000000010_010_0_110000000101;
      patterns[45075] = 29'b1_011000000010_011_1_100000001010;
      patterns[45076] = 29'b1_011000000010_100_0_101100000001;
      patterns[45077] = 29'b1_011000000010_101_1_010110000000;
      patterns[45078] = 29'b1_011000000010_110_1_011000000010;
      patterns[45079] = 29'b1_011000000010_111_1_011000000010;
      patterns[45080] = 29'b1_011000000011_000_1_011000000011;
      patterns[45081] = 29'b1_011000000011_001_1_000011011000;
      patterns[45082] = 29'b1_011000000011_010_0_110000000111;
      patterns[45083] = 29'b1_011000000011_011_1_100000001110;
      patterns[45084] = 29'b1_011000000011_100_1_101100000001;
      patterns[45085] = 29'b1_011000000011_101_1_110110000000;
      patterns[45086] = 29'b1_011000000011_110_1_011000000011;
      patterns[45087] = 29'b1_011000000011_111_1_011000000011;
      patterns[45088] = 29'b1_011000000100_000_1_011000000100;
      patterns[45089] = 29'b1_011000000100_001_1_000100011000;
      patterns[45090] = 29'b1_011000000100_010_0_110000001001;
      patterns[45091] = 29'b1_011000000100_011_1_100000010010;
      patterns[45092] = 29'b1_011000000100_100_0_101100000010;
      patterns[45093] = 29'b1_011000000100_101_0_010110000001;
      patterns[45094] = 29'b1_011000000100_110_1_011000000100;
      patterns[45095] = 29'b1_011000000100_111_1_011000000100;
      patterns[45096] = 29'b1_011000000101_000_1_011000000101;
      patterns[45097] = 29'b1_011000000101_001_1_000101011000;
      patterns[45098] = 29'b1_011000000101_010_0_110000001011;
      patterns[45099] = 29'b1_011000000101_011_1_100000010110;
      patterns[45100] = 29'b1_011000000101_100_1_101100000010;
      patterns[45101] = 29'b1_011000000101_101_0_110110000001;
      patterns[45102] = 29'b1_011000000101_110_1_011000000101;
      patterns[45103] = 29'b1_011000000101_111_1_011000000101;
      patterns[45104] = 29'b1_011000000110_000_1_011000000110;
      patterns[45105] = 29'b1_011000000110_001_1_000110011000;
      patterns[45106] = 29'b1_011000000110_010_0_110000001101;
      patterns[45107] = 29'b1_011000000110_011_1_100000011010;
      patterns[45108] = 29'b1_011000000110_100_0_101100000011;
      patterns[45109] = 29'b1_011000000110_101_1_010110000001;
      patterns[45110] = 29'b1_011000000110_110_1_011000000110;
      patterns[45111] = 29'b1_011000000110_111_1_011000000110;
      patterns[45112] = 29'b1_011000000111_000_1_011000000111;
      patterns[45113] = 29'b1_011000000111_001_1_000111011000;
      patterns[45114] = 29'b1_011000000111_010_0_110000001111;
      patterns[45115] = 29'b1_011000000111_011_1_100000011110;
      patterns[45116] = 29'b1_011000000111_100_1_101100000011;
      patterns[45117] = 29'b1_011000000111_101_1_110110000001;
      patterns[45118] = 29'b1_011000000111_110_1_011000000111;
      patterns[45119] = 29'b1_011000000111_111_1_011000000111;
      patterns[45120] = 29'b1_011000001000_000_1_011000001000;
      patterns[45121] = 29'b1_011000001000_001_1_001000011000;
      patterns[45122] = 29'b1_011000001000_010_0_110000010001;
      patterns[45123] = 29'b1_011000001000_011_1_100000100010;
      patterns[45124] = 29'b1_011000001000_100_0_101100000100;
      patterns[45125] = 29'b1_011000001000_101_0_010110000010;
      patterns[45126] = 29'b1_011000001000_110_1_011000001000;
      patterns[45127] = 29'b1_011000001000_111_1_011000001000;
      patterns[45128] = 29'b1_011000001001_000_1_011000001001;
      patterns[45129] = 29'b1_011000001001_001_1_001001011000;
      patterns[45130] = 29'b1_011000001001_010_0_110000010011;
      patterns[45131] = 29'b1_011000001001_011_1_100000100110;
      patterns[45132] = 29'b1_011000001001_100_1_101100000100;
      patterns[45133] = 29'b1_011000001001_101_0_110110000010;
      patterns[45134] = 29'b1_011000001001_110_1_011000001001;
      patterns[45135] = 29'b1_011000001001_111_1_011000001001;
      patterns[45136] = 29'b1_011000001010_000_1_011000001010;
      patterns[45137] = 29'b1_011000001010_001_1_001010011000;
      patterns[45138] = 29'b1_011000001010_010_0_110000010101;
      patterns[45139] = 29'b1_011000001010_011_1_100000101010;
      patterns[45140] = 29'b1_011000001010_100_0_101100000101;
      patterns[45141] = 29'b1_011000001010_101_1_010110000010;
      patterns[45142] = 29'b1_011000001010_110_1_011000001010;
      patterns[45143] = 29'b1_011000001010_111_1_011000001010;
      patterns[45144] = 29'b1_011000001011_000_1_011000001011;
      patterns[45145] = 29'b1_011000001011_001_1_001011011000;
      patterns[45146] = 29'b1_011000001011_010_0_110000010111;
      patterns[45147] = 29'b1_011000001011_011_1_100000101110;
      patterns[45148] = 29'b1_011000001011_100_1_101100000101;
      patterns[45149] = 29'b1_011000001011_101_1_110110000010;
      patterns[45150] = 29'b1_011000001011_110_1_011000001011;
      patterns[45151] = 29'b1_011000001011_111_1_011000001011;
      patterns[45152] = 29'b1_011000001100_000_1_011000001100;
      patterns[45153] = 29'b1_011000001100_001_1_001100011000;
      patterns[45154] = 29'b1_011000001100_010_0_110000011001;
      patterns[45155] = 29'b1_011000001100_011_1_100000110010;
      patterns[45156] = 29'b1_011000001100_100_0_101100000110;
      patterns[45157] = 29'b1_011000001100_101_0_010110000011;
      patterns[45158] = 29'b1_011000001100_110_1_011000001100;
      patterns[45159] = 29'b1_011000001100_111_1_011000001100;
      patterns[45160] = 29'b1_011000001101_000_1_011000001101;
      patterns[45161] = 29'b1_011000001101_001_1_001101011000;
      patterns[45162] = 29'b1_011000001101_010_0_110000011011;
      patterns[45163] = 29'b1_011000001101_011_1_100000110110;
      patterns[45164] = 29'b1_011000001101_100_1_101100000110;
      patterns[45165] = 29'b1_011000001101_101_0_110110000011;
      patterns[45166] = 29'b1_011000001101_110_1_011000001101;
      patterns[45167] = 29'b1_011000001101_111_1_011000001101;
      patterns[45168] = 29'b1_011000001110_000_1_011000001110;
      patterns[45169] = 29'b1_011000001110_001_1_001110011000;
      patterns[45170] = 29'b1_011000001110_010_0_110000011101;
      patterns[45171] = 29'b1_011000001110_011_1_100000111010;
      patterns[45172] = 29'b1_011000001110_100_0_101100000111;
      patterns[45173] = 29'b1_011000001110_101_1_010110000011;
      patterns[45174] = 29'b1_011000001110_110_1_011000001110;
      patterns[45175] = 29'b1_011000001110_111_1_011000001110;
      patterns[45176] = 29'b1_011000001111_000_1_011000001111;
      patterns[45177] = 29'b1_011000001111_001_1_001111011000;
      patterns[45178] = 29'b1_011000001111_010_0_110000011111;
      patterns[45179] = 29'b1_011000001111_011_1_100000111110;
      patterns[45180] = 29'b1_011000001111_100_1_101100000111;
      patterns[45181] = 29'b1_011000001111_101_1_110110000011;
      patterns[45182] = 29'b1_011000001111_110_1_011000001111;
      patterns[45183] = 29'b1_011000001111_111_1_011000001111;
      patterns[45184] = 29'b1_011000010000_000_1_011000010000;
      patterns[45185] = 29'b1_011000010000_001_1_010000011000;
      patterns[45186] = 29'b1_011000010000_010_0_110000100001;
      patterns[45187] = 29'b1_011000010000_011_1_100001000010;
      patterns[45188] = 29'b1_011000010000_100_0_101100001000;
      patterns[45189] = 29'b1_011000010000_101_0_010110000100;
      patterns[45190] = 29'b1_011000010000_110_1_011000010000;
      patterns[45191] = 29'b1_011000010000_111_1_011000010000;
      patterns[45192] = 29'b1_011000010001_000_1_011000010001;
      patterns[45193] = 29'b1_011000010001_001_1_010001011000;
      patterns[45194] = 29'b1_011000010001_010_0_110000100011;
      patterns[45195] = 29'b1_011000010001_011_1_100001000110;
      patterns[45196] = 29'b1_011000010001_100_1_101100001000;
      patterns[45197] = 29'b1_011000010001_101_0_110110000100;
      patterns[45198] = 29'b1_011000010001_110_1_011000010001;
      patterns[45199] = 29'b1_011000010001_111_1_011000010001;
      patterns[45200] = 29'b1_011000010010_000_1_011000010010;
      patterns[45201] = 29'b1_011000010010_001_1_010010011000;
      patterns[45202] = 29'b1_011000010010_010_0_110000100101;
      patterns[45203] = 29'b1_011000010010_011_1_100001001010;
      patterns[45204] = 29'b1_011000010010_100_0_101100001001;
      patterns[45205] = 29'b1_011000010010_101_1_010110000100;
      patterns[45206] = 29'b1_011000010010_110_1_011000010010;
      patterns[45207] = 29'b1_011000010010_111_1_011000010010;
      patterns[45208] = 29'b1_011000010011_000_1_011000010011;
      patterns[45209] = 29'b1_011000010011_001_1_010011011000;
      patterns[45210] = 29'b1_011000010011_010_0_110000100111;
      patterns[45211] = 29'b1_011000010011_011_1_100001001110;
      patterns[45212] = 29'b1_011000010011_100_1_101100001001;
      patterns[45213] = 29'b1_011000010011_101_1_110110000100;
      patterns[45214] = 29'b1_011000010011_110_1_011000010011;
      patterns[45215] = 29'b1_011000010011_111_1_011000010011;
      patterns[45216] = 29'b1_011000010100_000_1_011000010100;
      patterns[45217] = 29'b1_011000010100_001_1_010100011000;
      patterns[45218] = 29'b1_011000010100_010_0_110000101001;
      patterns[45219] = 29'b1_011000010100_011_1_100001010010;
      patterns[45220] = 29'b1_011000010100_100_0_101100001010;
      patterns[45221] = 29'b1_011000010100_101_0_010110000101;
      patterns[45222] = 29'b1_011000010100_110_1_011000010100;
      patterns[45223] = 29'b1_011000010100_111_1_011000010100;
      patterns[45224] = 29'b1_011000010101_000_1_011000010101;
      patterns[45225] = 29'b1_011000010101_001_1_010101011000;
      patterns[45226] = 29'b1_011000010101_010_0_110000101011;
      patterns[45227] = 29'b1_011000010101_011_1_100001010110;
      patterns[45228] = 29'b1_011000010101_100_1_101100001010;
      patterns[45229] = 29'b1_011000010101_101_0_110110000101;
      patterns[45230] = 29'b1_011000010101_110_1_011000010101;
      patterns[45231] = 29'b1_011000010101_111_1_011000010101;
      patterns[45232] = 29'b1_011000010110_000_1_011000010110;
      patterns[45233] = 29'b1_011000010110_001_1_010110011000;
      patterns[45234] = 29'b1_011000010110_010_0_110000101101;
      patterns[45235] = 29'b1_011000010110_011_1_100001011010;
      patterns[45236] = 29'b1_011000010110_100_0_101100001011;
      patterns[45237] = 29'b1_011000010110_101_1_010110000101;
      patterns[45238] = 29'b1_011000010110_110_1_011000010110;
      patterns[45239] = 29'b1_011000010110_111_1_011000010110;
      patterns[45240] = 29'b1_011000010111_000_1_011000010111;
      patterns[45241] = 29'b1_011000010111_001_1_010111011000;
      patterns[45242] = 29'b1_011000010111_010_0_110000101111;
      patterns[45243] = 29'b1_011000010111_011_1_100001011110;
      patterns[45244] = 29'b1_011000010111_100_1_101100001011;
      patterns[45245] = 29'b1_011000010111_101_1_110110000101;
      patterns[45246] = 29'b1_011000010111_110_1_011000010111;
      patterns[45247] = 29'b1_011000010111_111_1_011000010111;
      patterns[45248] = 29'b1_011000011000_000_1_011000011000;
      patterns[45249] = 29'b1_011000011000_001_1_011000011000;
      patterns[45250] = 29'b1_011000011000_010_0_110000110001;
      patterns[45251] = 29'b1_011000011000_011_1_100001100010;
      patterns[45252] = 29'b1_011000011000_100_0_101100001100;
      patterns[45253] = 29'b1_011000011000_101_0_010110000110;
      patterns[45254] = 29'b1_011000011000_110_1_011000011000;
      patterns[45255] = 29'b1_011000011000_111_1_011000011000;
      patterns[45256] = 29'b1_011000011001_000_1_011000011001;
      patterns[45257] = 29'b1_011000011001_001_1_011001011000;
      patterns[45258] = 29'b1_011000011001_010_0_110000110011;
      patterns[45259] = 29'b1_011000011001_011_1_100001100110;
      patterns[45260] = 29'b1_011000011001_100_1_101100001100;
      patterns[45261] = 29'b1_011000011001_101_0_110110000110;
      patterns[45262] = 29'b1_011000011001_110_1_011000011001;
      patterns[45263] = 29'b1_011000011001_111_1_011000011001;
      patterns[45264] = 29'b1_011000011010_000_1_011000011010;
      patterns[45265] = 29'b1_011000011010_001_1_011010011000;
      patterns[45266] = 29'b1_011000011010_010_0_110000110101;
      patterns[45267] = 29'b1_011000011010_011_1_100001101010;
      patterns[45268] = 29'b1_011000011010_100_0_101100001101;
      patterns[45269] = 29'b1_011000011010_101_1_010110000110;
      patterns[45270] = 29'b1_011000011010_110_1_011000011010;
      patterns[45271] = 29'b1_011000011010_111_1_011000011010;
      patterns[45272] = 29'b1_011000011011_000_1_011000011011;
      patterns[45273] = 29'b1_011000011011_001_1_011011011000;
      patterns[45274] = 29'b1_011000011011_010_0_110000110111;
      patterns[45275] = 29'b1_011000011011_011_1_100001101110;
      patterns[45276] = 29'b1_011000011011_100_1_101100001101;
      patterns[45277] = 29'b1_011000011011_101_1_110110000110;
      patterns[45278] = 29'b1_011000011011_110_1_011000011011;
      patterns[45279] = 29'b1_011000011011_111_1_011000011011;
      patterns[45280] = 29'b1_011000011100_000_1_011000011100;
      patterns[45281] = 29'b1_011000011100_001_1_011100011000;
      patterns[45282] = 29'b1_011000011100_010_0_110000111001;
      patterns[45283] = 29'b1_011000011100_011_1_100001110010;
      patterns[45284] = 29'b1_011000011100_100_0_101100001110;
      patterns[45285] = 29'b1_011000011100_101_0_010110000111;
      patterns[45286] = 29'b1_011000011100_110_1_011000011100;
      patterns[45287] = 29'b1_011000011100_111_1_011000011100;
      patterns[45288] = 29'b1_011000011101_000_1_011000011101;
      patterns[45289] = 29'b1_011000011101_001_1_011101011000;
      patterns[45290] = 29'b1_011000011101_010_0_110000111011;
      patterns[45291] = 29'b1_011000011101_011_1_100001110110;
      patterns[45292] = 29'b1_011000011101_100_1_101100001110;
      patterns[45293] = 29'b1_011000011101_101_0_110110000111;
      patterns[45294] = 29'b1_011000011101_110_1_011000011101;
      patterns[45295] = 29'b1_011000011101_111_1_011000011101;
      patterns[45296] = 29'b1_011000011110_000_1_011000011110;
      patterns[45297] = 29'b1_011000011110_001_1_011110011000;
      patterns[45298] = 29'b1_011000011110_010_0_110000111101;
      patterns[45299] = 29'b1_011000011110_011_1_100001111010;
      patterns[45300] = 29'b1_011000011110_100_0_101100001111;
      patterns[45301] = 29'b1_011000011110_101_1_010110000111;
      patterns[45302] = 29'b1_011000011110_110_1_011000011110;
      patterns[45303] = 29'b1_011000011110_111_1_011000011110;
      patterns[45304] = 29'b1_011000011111_000_1_011000011111;
      patterns[45305] = 29'b1_011000011111_001_1_011111011000;
      patterns[45306] = 29'b1_011000011111_010_0_110000111111;
      patterns[45307] = 29'b1_011000011111_011_1_100001111110;
      patterns[45308] = 29'b1_011000011111_100_1_101100001111;
      patterns[45309] = 29'b1_011000011111_101_1_110110000111;
      patterns[45310] = 29'b1_011000011111_110_1_011000011111;
      patterns[45311] = 29'b1_011000011111_111_1_011000011111;
      patterns[45312] = 29'b1_011000100000_000_1_011000100000;
      patterns[45313] = 29'b1_011000100000_001_1_100000011000;
      patterns[45314] = 29'b1_011000100000_010_0_110001000001;
      patterns[45315] = 29'b1_011000100000_011_1_100010000010;
      patterns[45316] = 29'b1_011000100000_100_0_101100010000;
      patterns[45317] = 29'b1_011000100000_101_0_010110001000;
      patterns[45318] = 29'b1_011000100000_110_1_011000100000;
      patterns[45319] = 29'b1_011000100000_111_1_011000100000;
      patterns[45320] = 29'b1_011000100001_000_1_011000100001;
      patterns[45321] = 29'b1_011000100001_001_1_100001011000;
      patterns[45322] = 29'b1_011000100001_010_0_110001000011;
      patterns[45323] = 29'b1_011000100001_011_1_100010000110;
      patterns[45324] = 29'b1_011000100001_100_1_101100010000;
      patterns[45325] = 29'b1_011000100001_101_0_110110001000;
      patterns[45326] = 29'b1_011000100001_110_1_011000100001;
      patterns[45327] = 29'b1_011000100001_111_1_011000100001;
      patterns[45328] = 29'b1_011000100010_000_1_011000100010;
      patterns[45329] = 29'b1_011000100010_001_1_100010011000;
      patterns[45330] = 29'b1_011000100010_010_0_110001000101;
      patterns[45331] = 29'b1_011000100010_011_1_100010001010;
      patterns[45332] = 29'b1_011000100010_100_0_101100010001;
      patterns[45333] = 29'b1_011000100010_101_1_010110001000;
      patterns[45334] = 29'b1_011000100010_110_1_011000100010;
      patterns[45335] = 29'b1_011000100010_111_1_011000100010;
      patterns[45336] = 29'b1_011000100011_000_1_011000100011;
      patterns[45337] = 29'b1_011000100011_001_1_100011011000;
      patterns[45338] = 29'b1_011000100011_010_0_110001000111;
      patterns[45339] = 29'b1_011000100011_011_1_100010001110;
      patterns[45340] = 29'b1_011000100011_100_1_101100010001;
      patterns[45341] = 29'b1_011000100011_101_1_110110001000;
      patterns[45342] = 29'b1_011000100011_110_1_011000100011;
      patterns[45343] = 29'b1_011000100011_111_1_011000100011;
      patterns[45344] = 29'b1_011000100100_000_1_011000100100;
      patterns[45345] = 29'b1_011000100100_001_1_100100011000;
      patterns[45346] = 29'b1_011000100100_010_0_110001001001;
      patterns[45347] = 29'b1_011000100100_011_1_100010010010;
      patterns[45348] = 29'b1_011000100100_100_0_101100010010;
      patterns[45349] = 29'b1_011000100100_101_0_010110001001;
      patterns[45350] = 29'b1_011000100100_110_1_011000100100;
      patterns[45351] = 29'b1_011000100100_111_1_011000100100;
      patterns[45352] = 29'b1_011000100101_000_1_011000100101;
      patterns[45353] = 29'b1_011000100101_001_1_100101011000;
      patterns[45354] = 29'b1_011000100101_010_0_110001001011;
      patterns[45355] = 29'b1_011000100101_011_1_100010010110;
      patterns[45356] = 29'b1_011000100101_100_1_101100010010;
      patterns[45357] = 29'b1_011000100101_101_0_110110001001;
      patterns[45358] = 29'b1_011000100101_110_1_011000100101;
      patterns[45359] = 29'b1_011000100101_111_1_011000100101;
      patterns[45360] = 29'b1_011000100110_000_1_011000100110;
      patterns[45361] = 29'b1_011000100110_001_1_100110011000;
      patterns[45362] = 29'b1_011000100110_010_0_110001001101;
      patterns[45363] = 29'b1_011000100110_011_1_100010011010;
      patterns[45364] = 29'b1_011000100110_100_0_101100010011;
      patterns[45365] = 29'b1_011000100110_101_1_010110001001;
      patterns[45366] = 29'b1_011000100110_110_1_011000100110;
      patterns[45367] = 29'b1_011000100110_111_1_011000100110;
      patterns[45368] = 29'b1_011000100111_000_1_011000100111;
      patterns[45369] = 29'b1_011000100111_001_1_100111011000;
      patterns[45370] = 29'b1_011000100111_010_0_110001001111;
      patterns[45371] = 29'b1_011000100111_011_1_100010011110;
      patterns[45372] = 29'b1_011000100111_100_1_101100010011;
      patterns[45373] = 29'b1_011000100111_101_1_110110001001;
      patterns[45374] = 29'b1_011000100111_110_1_011000100111;
      patterns[45375] = 29'b1_011000100111_111_1_011000100111;
      patterns[45376] = 29'b1_011000101000_000_1_011000101000;
      patterns[45377] = 29'b1_011000101000_001_1_101000011000;
      patterns[45378] = 29'b1_011000101000_010_0_110001010001;
      patterns[45379] = 29'b1_011000101000_011_1_100010100010;
      patterns[45380] = 29'b1_011000101000_100_0_101100010100;
      patterns[45381] = 29'b1_011000101000_101_0_010110001010;
      patterns[45382] = 29'b1_011000101000_110_1_011000101000;
      patterns[45383] = 29'b1_011000101000_111_1_011000101000;
      patterns[45384] = 29'b1_011000101001_000_1_011000101001;
      patterns[45385] = 29'b1_011000101001_001_1_101001011000;
      patterns[45386] = 29'b1_011000101001_010_0_110001010011;
      patterns[45387] = 29'b1_011000101001_011_1_100010100110;
      patterns[45388] = 29'b1_011000101001_100_1_101100010100;
      patterns[45389] = 29'b1_011000101001_101_0_110110001010;
      patterns[45390] = 29'b1_011000101001_110_1_011000101001;
      patterns[45391] = 29'b1_011000101001_111_1_011000101001;
      patterns[45392] = 29'b1_011000101010_000_1_011000101010;
      patterns[45393] = 29'b1_011000101010_001_1_101010011000;
      patterns[45394] = 29'b1_011000101010_010_0_110001010101;
      patterns[45395] = 29'b1_011000101010_011_1_100010101010;
      patterns[45396] = 29'b1_011000101010_100_0_101100010101;
      patterns[45397] = 29'b1_011000101010_101_1_010110001010;
      patterns[45398] = 29'b1_011000101010_110_1_011000101010;
      patterns[45399] = 29'b1_011000101010_111_1_011000101010;
      patterns[45400] = 29'b1_011000101011_000_1_011000101011;
      patterns[45401] = 29'b1_011000101011_001_1_101011011000;
      patterns[45402] = 29'b1_011000101011_010_0_110001010111;
      patterns[45403] = 29'b1_011000101011_011_1_100010101110;
      patterns[45404] = 29'b1_011000101011_100_1_101100010101;
      patterns[45405] = 29'b1_011000101011_101_1_110110001010;
      patterns[45406] = 29'b1_011000101011_110_1_011000101011;
      patterns[45407] = 29'b1_011000101011_111_1_011000101011;
      patterns[45408] = 29'b1_011000101100_000_1_011000101100;
      patterns[45409] = 29'b1_011000101100_001_1_101100011000;
      patterns[45410] = 29'b1_011000101100_010_0_110001011001;
      patterns[45411] = 29'b1_011000101100_011_1_100010110010;
      patterns[45412] = 29'b1_011000101100_100_0_101100010110;
      patterns[45413] = 29'b1_011000101100_101_0_010110001011;
      patterns[45414] = 29'b1_011000101100_110_1_011000101100;
      patterns[45415] = 29'b1_011000101100_111_1_011000101100;
      patterns[45416] = 29'b1_011000101101_000_1_011000101101;
      patterns[45417] = 29'b1_011000101101_001_1_101101011000;
      patterns[45418] = 29'b1_011000101101_010_0_110001011011;
      patterns[45419] = 29'b1_011000101101_011_1_100010110110;
      patterns[45420] = 29'b1_011000101101_100_1_101100010110;
      patterns[45421] = 29'b1_011000101101_101_0_110110001011;
      patterns[45422] = 29'b1_011000101101_110_1_011000101101;
      patterns[45423] = 29'b1_011000101101_111_1_011000101101;
      patterns[45424] = 29'b1_011000101110_000_1_011000101110;
      patterns[45425] = 29'b1_011000101110_001_1_101110011000;
      patterns[45426] = 29'b1_011000101110_010_0_110001011101;
      patterns[45427] = 29'b1_011000101110_011_1_100010111010;
      patterns[45428] = 29'b1_011000101110_100_0_101100010111;
      patterns[45429] = 29'b1_011000101110_101_1_010110001011;
      patterns[45430] = 29'b1_011000101110_110_1_011000101110;
      patterns[45431] = 29'b1_011000101110_111_1_011000101110;
      patterns[45432] = 29'b1_011000101111_000_1_011000101111;
      patterns[45433] = 29'b1_011000101111_001_1_101111011000;
      patterns[45434] = 29'b1_011000101111_010_0_110001011111;
      patterns[45435] = 29'b1_011000101111_011_1_100010111110;
      patterns[45436] = 29'b1_011000101111_100_1_101100010111;
      patterns[45437] = 29'b1_011000101111_101_1_110110001011;
      patterns[45438] = 29'b1_011000101111_110_1_011000101111;
      patterns[45439] = 29'b1_011000101111_111_1_011000101111;
      patterns[45440] = 29'b1_011000110000_000_1_011000110000;
      patterns[45441] = 29'b1_011000110000_001_1_110000011000;
      patterns[45442] = 29'b1_011000110000_010_0_110001100001;
      patterns[45443] = 29'b1_011000110000_011_1_100011000010;
      patterns[45444] = 29'b1_011000110000_100_0_101100011000;
      patterns[45445] = 29'b1_011000110000_101_0_010110001100;
      patterns[45446] = 29'b1_011000110000_110_1_011000110000;
      patterns[45447] = 29'b1_011000110000_111_1_011000110000;
      patterns[45448] = 29'b1_011000110001_000_1_011000110001;
      patterns[45449] = 29'b1_011000110001_001_1_110001011000;
      patterns[45450] = 29'b1_011000110001_010_0_110001100011;
      patterns[45451] = 29'b1_011000110001_011_1_100011000110;
      patterns[45452] = 29'b1_011000110001_100_1_101100011000;
      patterns[45453] = 29'b1_011000110001_101_0_110110001100;
      patterns[45454] = 29'b1_011000110001_110_1_011000110001;
      patterns[45455] = 29'b1_011000110001_111_1_011000110001;
      patterns[45456] = 29'b1_011000110010_000_1_011000110010;
      patterns[45457] = 29'b1_011000110010_001_1_110010011000;
      patterns[45458] = 29'b1_011000110010_010_0_110001100101;
      patterns[45459] = 29'b1_011000110010_011_1_100011001010;
      patterns[45460] = 29'b1_011000110010_100_0_101100011001;
      patterns[45461] = 29'b1_011000110010_101_1_010110001100;
      patterns[45462] = 29'b1_011000110010_110_1_011000110010;
      patterns[45463] = 29'b1_011000110010_111_1_011000110010;
      patterns[45464] = 29'b1_011000110011_000_1_011000110011;
      patterns[45465] = 29'b1_011000110011_001_1_110011011000;
      patterns[45466] = 29'b1_011000110011_010_0_110001100111;
      patterns[45467] = 29'b1_011000110011_011_1_100011001110;
      patterns[45468] = 29'b1_011000110011_100_1_101100011001;
      patterns[45469] = 29'b1_011000110011_101_1_110110001100;
      patterns[45470] = 29'b1_011000110011_110_1_011000110011;
      patterns[45471] = 29'b1_011000110011_111_1_011000110011;
      patterns[45472] = 29'b1_011000110100_000_1_011000110100;
      patterns[45473] = 29'b1_011000110100_001_1_110100011000;
      patterns[45474] = 29'b1_011000110100_010_0_110001101001;
      patterns[45475] = 29'b1_011000110100_011_1_100011010010;
      patterns[45476] = 29'b1_011000110100_100_0_101100011010;
      patterns[45477] = 29'b1_011000110100_101_0_010110001101;
      patterns[45478] = 29'b1_011000110100_110_1_011000110100;
      patterns[45479] = 29'b1_011000110100_111_1_011000110100;
      patterns[45480] = 29'b1_011000110101_000_1_011000110101;
      patterns[45481] = 29'b1_011000110101_001_1_110101011000;
      patterns[45482] = 29'b1_011000110101_010_0_110001101011;
      patterns[45483] = 29'b1_011000110101_011_1_100011010110;
      patterns[45484] = 29'b1_011000110101_100_1_101100011010;
      patterns[45485] = 29'b1_011000110101_101_0_110110001101;
      patterns[45486] = 29'b1_011000110101_110_1_011000110101;
      patterns[45487] = 29'b1_011000110101_111_1_011000110101;
      patterns[45488] = 29'b1_011000110110_000_1_011000110110;
      patterns[45489] = 29'b1_011000110110_001_1_110110011000;
      patterns[45490] = 29'b1_011000110110_010_0_110001101101;
      patterns[45491] = 29'b1_011000110110_011_1_100011011010;
      patterns[45492] = 29'b1_011000110110_100_0_101100011011;
      patterns[45493] = 29'b1_011000110110_101_1_010110001101;
      patterns[45494] = 29'b1_011000110110_110_1_011000110110;
      patterns[45495] = 29'b1_011000110110_111_1_011000110110;
      patterns[45496] = 29'b1_011000110111_000_1_011000110111;
      patterns[45497] = 29'b1_011000110111_001_1_110111011000;
      patterns[45498] = 29'b1_011000110111_010_0_110001101111;
      patterns[45499] = 29'b1_011000110111_011_1_100011011110;
      patterns[45500] = 29'b1_011000110111_100_1_101100011011;
      patterns[45501] = 29'b1_011000110111_101_1_110110001101;
      patterns[45502] = 29'b1_011000110111_110_1_011000110111;
      patterns[45503] = 29'b1_011000110111_111_1_011000110111;
      patterns[45504] = 29'b1_011000111000_000_1_011000111000;
      patterns[45505] = 29'b1_011000111000_001_1_111000011000;
      patterns[45506] = 29'b1_011000111000_010_0_110001110001;
      patterns[45507] = 29'b1_011000111000_011_1_100011100010;
      patterns[45508] = 29'b1_011000111000_100_0_101100011100;
      patterns[45509] = 29'b1_011000111000_101_0_010110001110;
      patterns[45510] = 29'b1_011000111000_110_1_011000111000;
      patterns[45511] = 29'b1_011000111000_111_1_011000111000;
      patterns[45512] = 29'b1_011000111001_000_1_011000111001;
      patterns[45513] = 29'b1_011000111001_001_1_111001011000;
      patterns[45514] = 29'b1_011000111001_010_0_110001110011;
      patterns[45515] = 29'b1_011000111001_011_1_100011100110;
      patterns[45516] = 29'b1_011000111001_100_1_101100011100;
      patterns[45517] = 29'b1_011000111001_101_0_110110001110;
      patterns[45518] = 29'b1_011000111001_110_1_011000111001;
      patterns[45519] = 29'b1_011000111001_111_1_011000111001;
      patterns[45520] = 29'b1_011000111010_000_1_011000111010;
      patterns[45521] = 29'b1_011000111010_001_1_111010011000;
      patterns[45522] = 29'b1_011000111010_010_0_110001110101;
      patterns[45523] = 29'b1_011000111010_011_1_100011101010;
      patterns[45524] = 29'b1_011000111010_100_0_101100011101;
      patterns[45525] = 29'b1_011000111010_101_1_010110001110;
      patterns[45526] = 29'b1_011000111010_110_1_011000111010;
      patterns[45527] = 29'b1_011000111010_111_1_011000111010;
      patterns[45528] = 29'b1_011000111011_000_1_011000111011;
      patterns[45529] = 29'b1_011000111011_001_1_111011011000;
      patterns[45530] = 29'b1_011000111011_010_0_110001110111;
      patterns[45531] = 29'b1_011000111011_011_1_100011101110;
      patterns[45532] = 29'b1_011000111011_100_1_101100011101;
      patterns[45533] = 29'b1_011000111011_101_1_110110001110;
      patterns[45534] = 29'b1_011000111011_110_1_011000111011;
      patterns[45535] = 29'b1_011000111011_111_1_011000111011;
      patterns[45536] = 29'b1_011000111100_000_1_011000111100;
      patterns[45537] = 29'b1_011000111100_001_1_111100011000;
      patterns[45538] = 29'b1_011000111100_010_0_110001111001;
      patterns[45539] = 29'b1_011000111100_011_1_100011110010;
      patterns[45540] = 29'b1_011000111100_100_0_101100011110;
      patterns[45541] = 29'b1_011000111100_101_0_010110001111;
      patterns[45542] = 29'b1_011000111100_110_1_011000111100;
      patterns[45543] = 29'b1_011000111100_111_1_011000111100;
      patterns[45544] = 29'b1_011000111101_000_1_011000111101;
      patterns[45545] = 29'b1_011000111101_001_1_111101011000;
      patterns[45546] = 29'b1_011000111101_010_0_110001111011;
      patterns[45547] = 29'b1_011000111101_011_1_100011110110;
      patterns[45548] = 29'b1_011000111101_100_1_101100011110;
      patterns[45549] = 29'b1_011000111101_101_0_110110001111;
      patterns[45550] = 29'b1_011000111101_110_1_011000111101;
      patterns[45551] = 29'b1_011000111101_111_1_011000111101;
      patterns[45552] = 29'b1_011000111110_000_1_011000111110;
      patterns[45553] = 29'b1_011000111110_001_1_111110011000;
      patterns[45554] = 29'b1_011000111110_010_0_110001111101;
      patterns[45555] = 29'b1_011000111110_011_1_100011111010;
      patterns[45556] = 29'b1_011000111110_100_0_101100011111;
      patterns[45557] = 29'b1_011000111110_101_1_010110001111;
      patterns[45558] = 29'b1_011000111110_110_1_011000111110;
      patterns[45559] = 29'b1_011000111110_111_1_011000111110;
      patterns[45560] = 29'b1_011000111111_000_1_011000111111;
      patterns[45561] = 29'b1_011000111111_001_1_111111011000;
      patterns[45562] = 29'b1_011000111111_010_0_110001111111;
      patterns[45563] = 29'b1_011000111111_011_1_100011111110;
      patterns[45564] = 29'b1_011000111111_100_1_101100011111;
      patterns[45565] = 29'b1_011000111111_101_1_110110001111;
      patterns[45566] = 29'b1_011000111111_110_1_011000111111;
      patterns[45567] = 29'b1_011000111111_111_1_011000111111;
      patterns[45568] = 29'b1_011001000000_000_1_011001000000;
      patterns[45569] = 29'b1_011001000000_001_1_000000011001;
      patterns[45570] = 29'b1_011001000000_010_0_110010000001;
      patterns[45571] = 29'b1_011001000000_011_1_100100000010;
      patterns[45572] = 29'b1_011001000000_100_0_101100100000;
      patterns[45573] = 29'b1_011001000000_101_0_010110010000;
      patterns[45574] = 29'b1_011001000000_110_1_011001000000;
      patterns[45575] = 29'b1_011001000000_111_1_011001000000;
      patterns[45576] = 29'b1_011001000001_000_1_011001000001;
      patterns[45577] = 29'b1_011001000001_001_1_000001011001;
      patterns[45578] = 29'b1_011001000001_010_0_110010000011;
      patterns[45579] = 29'b1_011001000001_011_1_100100000110;
      patterns[45580] = 29'b1_011001000001_100_1_101100100000;
      patterns[45581] = 29'b1_011001000001_101_0_110110010000;
      patterns[45582] = 29'b1_011001000001_110_1_011001000001;
      patterns[45583] = 29'b1_011001000001_111_1_011001000001;
      patterns[45584] = 29'b1_011001000010_000_1_011001000010;
      patterns[45585] = 29'b1_011001000010_001_1_000010011001;
      patterns[45586] = 29'b1_011001000010_010_0_110010000101;
      patterns[45587] = 29'b1_011001000010_011_1_100100001010;
      patterns[45588] = 29'b1_011001000010_100_0_101100100001;
      patterns[45589] = 29'b1_011001000010_101_1_010110010000;
      patterns[45590] = 29'b1_011001000010_110_1_011001000010;
      patterns[45591] = 29'b1_011001000010_111_1_011001000010;
      patterns[45592] = 29'b1_011001000011_000_1_011001000011;
      patterns[45593] = 29'b1_011001000011_001_1_000011011001;
      patterns[45594] = 29'b1_011001000011_010_0_110010000111;
      patterns[45595] = 29'b1_011001000011_011_1_100100001110;
      patterns[45596] = 29'b1_011001000011_100_1_101100100001;
      patterns[45597] = 29'b1_011001000011_101_1_110110010000;
      patterns[45598] = 29'b1_011001000011_110_1_011001000011;
      patterns[45599] = 29'b1_011001000011_111_1_011001000011;
      patterns[45600] = 29'b1_011001000100_000_1_011001000100;
      patterns[45601] = 29'b1_011001000100_001_1_000100011001;
      patterns[45602] = 29'b1_011001000100_010_0_110010001001;
      patterns[45603] = 29'b1_011001000100_011_1_100100010010;
      patterns[45604] = 29'b1_011001000100_100_0_101100100010;
      patterns[45605] = 29'b1_011001000100_101_0_010110010001;
      patterns[45606] = 29'b1_011001000100_110_1_011001000100;
      patterns[45607] = 29'b1_011001000100_111_1_011001000100;
      patterns[45608] = 29'b1_011001000101_000_1_011001000101;
      patterns[45609] = 29'b1_011001000101_001_1_000101011001;
      patterns[45610] = 29'b1_011001000101_010_0_110010001011;
      patterns[45611] = 29'b1_011001000101_011_1_100100010110;
      patterns[45612] = 29'b1_011001000101_100_1_101100100010;
      patterns[45613] = 29'b1_011001000101_101_0_110110010001;
      patterns[45614] = 29'b1_011001000101_110_1_011001000101;
      patterns[45615] = 29'b1_011001000101_111_1_011001000101;
      patterns[45616] = 29'b1_011001000110_000_1_011001000110;
      patterns[45617] = 29'b1_011001000110_001_1_000110011001;
      patterns[45618] = 29'b1_011001000110_010_0_110010001101;
      patterns[45619] = 29'b1_011001000110_011_1_100100011010;
      patterns[45620] = 29'b1_011001000110_100_0_101100100011;
      patterns[45621] = 29'b1_011001000110_101_1_010110010001;
      patterns[45622] = 29'b1_011001000110_110_1_011001000110;
      patterns[45623] = 29'b1_011001000110_111_1_011001000110;
      patterns[45624] = 29'b1_011001000111_000_1_011001000111;
      patterns[45625] = 29'b1_011001000111_001_1_000111011001;
      patterns[45626] = 29'b1_011001000111_010_0_110010001111;
      patterns[45627] = 29'b1_011001000111_011_1_100100011110;
      patterns[45628] = 29'b1_011001000111_100_1_101100100011;
      patterns[45629] = 29'b1_011001000111_101_1_110110010001;
      patterns[45630] = 29'b1_011001000111_110_1_011001000111;
      patterns[45631] = 29'b1_011001000111_111_1_011001000111;
      patterns[45632] = 29'b1_011001001000_000_1_011001001000;
      patterns[45633] = 29'b1_011001001000_001_1_001000011001;
      patterns[45634] = 29'b1_011001001000_010_0_110010010001;
      patterns[45635] = 29'b1_011001001000_011_1_100100100010;
      patterns[45636] = 29'b1_011001001000_100_0_101100100100;
      patterns[45637] = 29'b1_011001001000_101_0_010110010010;
      patterns[45638] = 29'b1_011001001000_110_1_011001001000;
      patterns[45639] = 29'b1_011001001000_111_1_011001001000;
      patterns[45640] = 29'b1_011001001001_000_1_011001001001;
      patterns[45641] = 29'b1_011001001001_001_1_001001011001;
      patterns[45642] = 29'b1_011001001001_010_0_110010010011;
      patterns[45643] = 29'b1_011001001001_011_1_100100100110;
      patterns[45644] = 29'b1_011001001001_100_1_101100100100;
      patterns[45645] = 29'b1_011001001001_101_0_110110010010;
      patterns[45646] = 29'b1_011001001001_110_1_011001001001;
      patterns[45647] = 29'b1_011001001001_111_1_011001001001;
      patterns[45648] = 29'b1_011001001010_000_1_011001001010;
      patterns[45649] = 29'b1_011001001010_001_1_001010011001;
      patterns[45650] = 29'b1_011001001010_010_0_110010010101;
      patterns[45651] = 29'b1_011001001010_011_1_100100101010;
      patterns[45652] = 29'b1_011001001010_100_0_101100100101;
      patterns[45653] = 29'b1_011001001010_101_1_010110010010;
      patterns[45654] = 29'b1_011001001010_110_1_011001001010;
      patterns[45655] = 29'b1_011001001010_111_1_011001001010;
      patterns[45656] = 29'b1_011001001011_000_1_011001001011;
      patterns[45657] = 29'b1_011001001011_001_1_001011011001;
      patterns[45658] = 29'b1_011001001011_010_0_110010010111;
      patterns[45659] = 29'b1_011001001011_011_1_100100101110;
      patterns[45660] = 29'b1_011001001011_100_1_101100100101;
      patterns[45661] = 29'b1_011001001011_101_1_110110010010;
      patterns[45662] = 29'b1_011001001011_110_1_011001001011;
      patterns[45663] = 29'b1_011001001011_111_1_011001001011;
      patterns[45664] = 29'b1_011001001100_000_1_011001001100;
      patterns[45665] = 29'b1_011001001100_001_1_001100011001;
      patterns[45666] = 29'b1_011001001100_010_0_110010011001;
      patterns[45667] = 29'b1_011001001100_011_1_100100110010;
      patterns[45668] = 29'b1_011001001100_100_0_101100100110;
      patterns[45669] = 29'b1_011001001100_101_0_010110010011;
      patterns[45670] = 29'b1_011001001100_110_1_011001001100;
      patterns[45671] = 29'b1_011001001100_111_1_011001001100;
      patterns[45672] = 29'b1_011001001101_000_1_011001001101;
      patterns[45673] = 29'b1_011001001101_001_1_001101011001;
      patterns[45674] = 29'b1_011001001101_010_0_110010011011;
      patterns[45675] = 29'b1_011001001101_011_1_100100110110;
      patterns[45676] = 29'b1_011001001101_100_1_101100100110;
      patterns[45677] = 29'b1_011001001101_101_0_110110010011;
      patterns[45678] = 29'b1_011001001101_110_1_011001001101;
      patterns[45679] = 29'b1_011001001101_111_1_011001001101;
      patterns[45680] = 29'b1_011001001110_000_1_011001001110;
      patterns[45681] = 29'b1_011001001110_001_1_001110011001;
      patterns[45682] = 29'b1_011001001110_010_0_110010011101;
      patterns[45683] = 29'b1_011001001110_011_1_100100111010;
      patterns[45684] = 29'b1_011001001110_100_0_101100100111;
      patterns[45685] = 29'b1_011001001110_101_1_010110010011;
      patterns[45686] = 29'b1_011001001110_110_1_011001001110;
      patterns[45687] = 29'b1_011001001110_111_1_011001001110;
      patterns[45688] = 29'b1_011001001111_000_1_011001001111;
      patterns[45689] = 29'b1_011001001111_001_1_001111011001;
      patterns[45690] = 29'b1_011001001111_010_0_110010011111;
      patterns[45691] = 29'b1_011001001111_011_1_100100111110;
      patterns[45692] = 29'b1_011001001111_100_1_101100100111;
      patterns[45693] = 29'b1_011001001111_101_1_110110010011;
      patterns[45694] = 29'b1_011001001111_110_1_011001001111;
      patterns[45695] = 29'b1_011001001111_111_1_011001001111;
      patterns[45696] = 29'b1_011001010000_000_1_011001010000;
      patterns[45697] = 29'b1_011001010000_001_1_010000011001;
      patterns[45698] = 29'b1_011001010000_010_0_110010100001;
      patterns[45699] = 29'b1_011001010000_011_1_100101000010;
      patterns[45700] = 29'b1_011001010000_100_0_101100101000;
      patterns[45701] = 29'b1_011001010000_101_0_010110010100;
      patterns[45702] = 29'b1_011001010000_110_1_011001010000;
      patterns[45703] = 29'b1_011001010000_111_1_011001010000;
      patterns[45704] = 29'b1_011001010001_000_1_011001010001;
      patterns[45705] = 29'b1_011001010001_001_1_010001011001;
      patterns[45706] = 29'b1_011001010001_010_0_110010100011;
      patterns[45707] = 29'b1_011001010001_011_1_100101000110;
      patterns[45708] = 29'b1_011001010001_100_1_101100101000;
      patterns[45709] = 29'b1_011001010001_101_0_110110010100;
      patterns[45710] = 29'b1_011001010001_110_1_011001010001;
      patterns[45711] = 29'b1_011001010001_111_1_011001010001;
      patterns[45712] = 29'b1_011001010010_000_1_011001010010;
      patterns[45713] = 29'b1_011001010010_001_1_010010011001;
      patterns[45714] = 29'b1_011001010010_010_0_110010100101;
      patterns[45715] = 29'b1_011001010010_011_1_100101001010;
      patterns[45716] = 29'b1_011001010010_100_0_101100101001;
      patterns[45717] = 29'b1_011001010010_101_1_010110010100;
      patterns[45718] = 29'b1_011001010010_110_1_011001010010;
      patterns[45719] = 29'b1_011001010010_111_1_011001010010;
      patterns[45720] = 29'b1_011001010011_000_1_011001010011;
      patterns[45721] = 29'b1_011001010011_001_1_010011011001;
      patterns[45722] = 29'b1_011001010011_010_0_110010100111;
      patterns[45723] = 29'b1_011001010011_011_1_100101001110;
      patterns[45724] = 29'b1_011001010011_100_1_101100101001;
      patterns[45725] = 29'b1_011001010011_101_1_110110010100;
      patterns[45726] = 29'b1_011001010011_110_1_011001010011;
      patterns[45727] = 29'b1_011001010011_111_1_011001010011;
      patterns[45728] = 29'b1_011001010100_000_1_011001010100;
      patterns[45729] = 29'b1_011001010100_001_1_010100011001;
      patterns[45730] = 29'b1_011001010100_010_0_110010101001;
      patterns[45731] = 29'b1_011001010100_011_1_100101010010;
      patterns[45732] = 29'b1_011001010100_100_0_101100101010;
      patterns[45733] = 29'b1_011001010100_101_0_010110010101;
      patterns[45734] = 29'b1_011001010100_110_1_011001010100;
      patterns[45735] = 29'b1_011001010100_111_1_011001010100;
      patterns[45736] = 29'b1_011001010101_000_1_011001010101;
      patterns[45737] = 29'b1_011001010101_001_1_010101011001;
      patterns[45738] = 29'b1_011001010101_010_0_110010101011;
      patterns[45739] = 29'b1_011001010101_011_1_100101010110;
      patterns[45740] = 29'b1_011001010101_100_1_101100101010;
      patterns[45741] = 29'b1_011001010101_101_0_110110010101;
      patterns[45742] = 29'b1_011001010101_110_1_011001010101;
      patterns[45743] = 29'b1_011001010101_111_1_011001010101;
      patterns[45744] = 29'b1_011001010110_000_1_011001010110;
      patterns[45745] = 29'b1_011001010110_001_1_010110011001;
      patterns[45746] = 29'b1_011001010110_010_0_110010101101;
      patterns[45747] = 29'b1_011001010110_011_1_100101011010;
      patterns[45748] = 29'b1_011001010110_100_0_101100101011;
      patterns[45749] = 29'b1_011001010110_101_1_010110010101;
      patterns[45750] = 29'b1_011001010110_110_1_011001010110;
      patterns[45751] = 29'b1_011001010110_111_1_011001010110;
      patterns[45752] = 29'b1_011001010111_000_1_011001010111;
      patterns[45753] = 29'b1_011001010111_001_1_010111011001;
      patterns[45754] = 29'b1_011001010111_010_0_110010101111;
      patterns[45755] = 29'b1_011001010111_011_1_100101011110;
      patterns[45756] = 29'b1_011001010111_100_1_101100101011;
      patterns[45757] = 29'b1_011001010111_101_1_110110010101;
      patterns[45758] = 29'b1_011001010111_110_1_011001010111;
      patterns[45759] = 29'b1_011001010111_111_1_011001010111;
      patterns[45760] = 29'b1_011001011000_000_1_011001011000;
      patterns[45761] = 29'b1_011001011000_001_1_011000011001;
      patterns[45762] = 29'b1_011001011000_010_0_110010110001;
      patterns[45763] = 29'b1_011001011000_011_1_100101100010;
      patterns[45764] = 29'b1_011001011000_100_0_101100101100;
      patterns[45765] = 29'b1_011001011000_101_0_010110010110;
      patterns[45766] = 29'b1_011001011000_110_1_011001011000;
      patterns[45767] = 29'b1_011001011000_111_1_011001011000;
      patterns[45768] = 29'b1_011001011001_000_1_011001011001;
      patterns[45769] = 29'b1_011001011001_001_1_011001011001;
      patterns[45770] = 29'b1_011001011001_010_0_110010110011;
      patterns[45771] = 29'b1_011001011001_011_1_100101100110;
      patterns[45772] = 29'b1_011001011001_100_1_101100101100;
      patterns[45773] = 29'b1_011001011001_101_0_110110010110;
      patterns[45774] = 29'b1_011001011001_110_1_011001011001;
      patterns[45775] = 29'b1_011001011001_111_1_011001011001;
      patterns[45776] = 29'b1_011001011010_000_1_011001011010;
      patterns[45777] = 29'b1_011001011010_001_1_011010011001;
      patterns[45778] = 29'b1_011001011010_010_0_110010110101;
      patterns[45779] = 29'b1_011001011010_011_1_100101101010;
      patterns[45780] = 29'b1_011001011010_100_0_101100101101;
      patterns[45781] = 29'b1_011001011010_101_1_010110010110;
      patterns[45782] = 29'b1_011001011010_110_1_011001011010;
      patterns[45783] = 29'b1_011001011010_111_1_011001011010;
      patterns[45784] = 29'b1_011001011011_000_1_011001011011;
      patterns[45785] = 29'b1_011001011011_001_1_011011011001;
      patterns[45786] = 29'b1_011001011011_010_0_110010110111;
      patterns[45787] = 29'b1_011001011011_011_1_100101101110;
      patterns[45788] = 29'b1_011001011011_100_1_101100101101;
      patterns[45789] = 29'b1_011001011011_101_1_110110010110;
      patterns[45790] = 29'b1_011001011011_110_1_011001011011;
      patterns[45791] = 29'b1_011001011011_111_1_011001011011;
      patterns[45792] = 29'b1_011001011100_000_1_011001011100;
      patterns[45793] = 29'b1_011001011100_001_1_011100011001;
      patterns[45794] = 29'b1_011001011100_010_0_110010111001;
      patterns[45795] = 29'b1_011001011100_011_1_100101110010;
      patterns[45796] = 29'b1_011001011100_100_0_101100101110;
      patterns[45797] = 29'b1_011001011100_101_0_010110010111;
      patterns[45798] = 29'b1_011001011100_110_1_011001011100;
      patterns[45799] = 29'b1_011001011100_111_1_011001011100;
      patterns[45800] = 29'b1_011001011101_000_1_011001011101;
      patterns[45801] = 29'b1_011001011101_001_1_011101011001;
      patterns[45802] = 29'b1_011001011101_010_0_110010111011;
      patterns[45803] = 29'b1_011001011101_011_1_100101110110;
      patterns[45804] = 29'b1_011001011101_100_1_101100101110;
      patterns[45805] = 29'b1_011001011101_101_0_110110010111;
      patterns[45806] = 29'b1_011001011101_110_1_011001011101;
      patterns[45807] = 29'b1_011001011101_111_1_011001011101;
      patterns[45808] = 29'b1_011001011110_000_1_011001011110;
      patterns[45809] = 29'b1_011001011110_001_1_011110011001;
      patterns[45810] = 29'b1_011001011110_010_0_110010111101;
      patterns[45811] = 29'b1_011001011110_011_1_100101111010;
      patterns[45812] = 29'b1_011001011110_100_0_101100101111;
      patterns[45813] = 29'b1_011001011110_101_1_010110010111;
      patterns[45814] = 29'b1_011001011110_110_1_011001011110;
      patterns[45815] = 29'b1_011001011110_111_1_011001011110;
      patterns[45816] = 29'b1_011001011111_000_1_011001011111;
      patterns[45817] = 29'b1_011001011111_001_1_011111011001;
      patterns[45818] = 29'b1_011001011111_010_0_110010111111;
      patterns[45819] = 29'b1_011001011111_011_1_100101111110;
      patterns[45820] = 29'b1_011001011111_100_1_101100101111;
      patterns[45821] = 29'b1_011001011111_101_1_110110010111;
      patterns[45822] = 29'b1_011001011111_110_1_011001011111;
      patterns[45823] = 29'b1_011001011111_111_1_011001011111;
      patterns[45824] = 29'b1_011001100000_000_1_011001100000;
      patterns[45825] = 29'b1_011001100000_001_1_100000011001;
      patterns[45826] = 29'b1_011001100000_010_0_110011000001;
      patterns[45827] = 29'b1_011001100000_011_1_100110000010;
      patterns[45828] = 29'b1_011001100000_100_0_101100110000;
      patterns[45829] = 29'b1_011001100000_101_0_010110011000;
      patterns[45830] = 29'b1_011001100000_110_1_011001100000;
      patterns[45831] = 29'b1_011001100000_111_1_011001100000;
      patterns[45832] = 29'b1_011001100001_000_1_011001100001;
      patterns[45833] = 29'b1_011001100001_001_1_100001011001;
      patterns[45834] = 29'b1_011001100001_010_0_110011000011;
      patterns[45835] = 29'b1_011001100001_011_1_100110000110;
      patterns[45836] = 29'b1_011001100001_100_1_101100110000;
      patterns[45837] = 29'b1_011001100001_101_0_110110011000;
      patterns[45838] = 29'b1_011001100001_110_1_011001100001;
      patterns[45839] = 29'b1_011001100001_111_1_011001100001;
      patterns[45840] = 29'b1_011001100010_000_1_011001100010;
      patterns[45841] = 29'b1_011001100010_001_1_100010011001;
      patterns[45842] = 29'b1_011001100010_010_0_110011000101;
      patterns[45843] = 29'b1_011001100010_011_1_100110001010;
      patterns[45844] = 29'b1_011001100010_100_0_101100110001;
      patterns[45845] = 29'b1_011001100010_101_1_010110011000;
      patterns[45846] = 29'b1_011001100010_110_1_011001100010;
      patterns[45847] = 29'b1_011001100010_111_1_011001100010;
      patterns[45848] = 29'b1_011001100011_000_1_011001100011;
      patterns[45849] = 29'b1_011001100011_001_1_100011011001;
      patterns[45850] = 29'b1_011001100011_010_0_110011000111;
      patterns[45851] = 29'b1_011001100011_011_1_100110001110;
      patterns[45852] = 29'b1_011001100011_100_1_101100110001;
      patterns[45853] = 29'b1_011001100011_101_1_110110011000;
      patterns[45854] = 29'b1_011001100011_110_1_011001100011;
      patterns[45855] = 29'b1_011001100011_111_1_011001100011;
      patterns[45856] = 29'b1_011001100100_000_1_011001100100;
      patterns[45857] = 29'b1_011001100100_001_1_100100011001;
      patterns[45858] = 29'b1_011001100100_010_0_110011001001;
      patterns[45859] = 29'b1_011001100100_011_1_100110010010;
      patterns[45860] = 29'b1_011001100100_100_0_101100110010;
      patterns[45861] = 29'b1_011001100100_101_0_010110011001;
      patterns[45862] = 29'b1_011001100100_110_1_011001100100;
      patterns[45863] = 29'b1_011001100100_111_1_011001100100;
      patterns[45864] = 29'b1_011001100101_000_1_011001100101;
      patterns[45865] = 29'b1_011001100101_001_1_100101011001;
      patterns[45866] = 29'b1_011001100101_010_0_110011001011;
      patterns[45867] = 29'b1_011001100101_011_1_100110010110;
      patterns[45868] = 29'b1_011001100101_100_1_101100110010;
      patterns[45869] = 29'b1_011001100101_101_0_110110011001;
      patterns[45870] = 29'b1_011001100101_110_1_011001100101;
      patterns[45871] = 29'b1_011001100101_111_1_011001100101;
      patterns[45872] = 29'b1_011001100110_000_1_011001100110;
      patterns[45873] = 29'b1_011001100110_001_1_100110011001;
      patterns[45874] = 29'b1_011001100110_010_0_110011001101;
      patterns[45875] = 29'b1_011001100110_011_1_100110011010;
      patterns[45876] = 29'b1_011001100110_100_0_101100110011;
      patterns[45877] = 29'b1_011001100110_101_1_010110011001;
      patterns[45878] = 29'b1_011001100110_110_1_011001100110;
      patterns[45879] = 29'b1_011001100110_111_1_011001100110;
      patterns[45880] = 29'b1_011001100111_000_1_011001100111;
      patterns[45881] = 29'b1_011001100111_001_1_100111011001;
      patterns[45882] = 29'b1_011001100111_010_0_110011001111;
      patterns[45883] = 29'b1_011001100111_011_1_100110011110;
      patterns[45884] = 29'b1_011001100111_100_1_101100110011;
      patterns[45885] = 29'b1_011001100111_101_1_110110011001;
      patterns[45886] = 29'b1_011001100111_110_1_011001100111;
      patterns[45887] = 29'b1_011001100111_111_1_011001100111;
      patterns[45888] = 29'b1_011001101000_000_1_011001101000;
      patterns[45889] = 29'b1_011001101000_001_1_101000011001;
      patterns[45890] = 29'b1_011001101000_010_0_110011010001;
      patterns[45891] = 29'b1_011001101000_011_1_100110100010;
      patterns[45892] = 29'b1_011001101000_100_0_101100110100;
      patterns[45893] = 29'b1_011001101000_101_0_010110011010;
      patterns[45894] = 29'b1_011001101000_110_1_011001101000;
      patterns[45895] = 29'b1_011001101000_111_1_011001101000;
      patterns[45896] = 29'b1_011001101001_000_1_011001101001;
      patterns[45897] = 29'b1_011001101001_001_1_101001011001;
      patterns[45898] = 29'b1_011001101001_010_0_110011010011;
      patterns[45899] = 29'b1_011001101001_011_1_100110100110;
      patterns[45900] = 29'b1_011001101001_100_1_101100110100;
      patterns[45901] = 29'b1_011001101001_101_0_110110011010;
      patterns[45902] = 29'b1_011001101001_110_1_011001101001;
      patterns[45903] = 29'b1_011001101001_111_1_011001101001;
      patterns[45904] = 29'b1_011001101010_000_1_011001101010;
      patterns[45905] = 29'b1_011001101010_001_1_101010011001;
      patterns[45906] = 29'b1_011001101010_010_0_110011010101;
      patterns[45907] = 29'b1_011001101010_011_1_100110101010;
      patterns[45908] = 29'b1_011001101010_100_0_101100110101;
      patterns[45909] = 29'b1_011001101010_101_1_010110011010;
      patterns[45910] = 29'b1_011001101010_110_1_011001101010;
      patterns[45911] = 29'b1_011001101010_111_1_011001101010;
      patterns[45912] = 29'b1_011001101011_000_1_011001101011;
      patterns[45913] = 29'b1_011001101011_001_1_101011011001;
      patterns[45914] = 29'b1_011001101011_010_0_110011010111;
      patterns[45915] = 29'b1_011001101011_011_1_100110101110;
      patterns[45916] = 29'b1_011001101011_100_1_101100110101;
      patterns[45917] = 29'b1_011001101011_101_1_110110011010;
      patterns[45918] = 29'b1_011001101011_110_1_011001101011;
      patterns[45919] = 29'b1_011001101011_111_1_011001101011;
      patterns[45920] = 29'b1_011001101100_000_1_011001101100;
      patterns[45921] = 29'b1_011001101100_001_1_101100011001;
      patterns[45922] = 29'b1_011001101100_010_0_110011011001;
      patterns[45923] = 29'b1_011001101100_011_1_100110110010;
      patterns[45924] = 29'b1_011001101100_100_0_101100110110;
      patterns[45925] = 29'b1_011001101100_101_0_010110011011;
      patterns[45926] = 29'b1_011001101100_110_1_011001101100;
      patterns[45927] = 29'b1_011001101100_111_1_011001101100;
      patterns[45928] = 29'b1_011001101101_000_1_011001101101;
      patterns[45929] = 29'b1_011001101101_001_1_101101011001;
      patterns[45930] = 29'b1_011001101101_010_0_110011011011;
      patterns[45931] = 29'b1_011001101101_011_1_100110110110;
      patterns[45932] = 29'b1_011001101101_100_1_101100110110;
      patterns[45933] = 29'b1_011001101101_101_0_110110011011;
      patterns[45934] = 29'b1_011001101101_110_1_011001101101;
      patterns[45935] = 29'b1_011001101101_111_1_011001101101;
      patterns[45936] = 29'b1_011001101110_000_1_011001101110;
      patterns[45937] = 29'b1_011001101110_001_1_101110011001;
      patterns[45938] = 29'b1_011001101110_010_0_110011011101;
      patterns[45939] = 29'b1_011001101110_011_1_100110111010;
      patterns[45940] = 29'b1_011001101110_100_0_101100110111;
      patterns[45941] = 29'b1_011001101110_101_1_010110011011;
      patterns[45942] = 29'b1_011001101110_110_1_011001101110;
      patterns[45943] = 29'b1_011001101110_111_1_011001101110;
      patterns[45944] = 29'b1_011001101111_000_1_011001101111;
      patterns[45945] = 29'b1_011001101111_001_1_101111011001;
      patterns[45946] = 29'b1_011001101111_010_0_110011011111;
      patterns[45947] = 29'b1_011001101111_011_1_100110111110;
      patterns[45948] = 29'b1_011001101111_100_1_101100110111;
      patterns[45949] = 29'b1_011001101111_101_1_110110011011;
      patterns[45950] = 29'b1_011001101111_110_1_011001101111;
      patterns[45951] = 29'b1_011001101111_111_1_011001101111;
      patterns[45952] = 29'b1_011001110000_000_1_011001110000;
      patterns[45953] = 29'b1_011001110000_001_1_110000011001;
      patterns[45954] = 29'b1_011001110000_010_0_110011100001;
      patterns[45955] = 29'b1_011001110000_011_1_100111000010;
      patterns[45956] = 29'b1_011001110000_100_0_101100111000;
      patterns[45957] = 29'b1_011001110000_101_0_010110011100;
      patterns[45958] = 29'b1_011001110000_110_1_011001110000;
      patterns[45959] = 29'b1_011001110000_111_1_011001110000;
      patterns[45960] = 29'b1_011001110001_000_1_011001110001;
      patterns[45961] = 29'b1_011001110001_001_1_110001011001;
      patterns[45962] = 29'b1_011001110001_010_0_110011100011;
      patterns[45963] = 29'b1_011001110001_011_1_100111000110;
      patterns[45964] = 29'b1_011001110001_100_1_101100111000;
      patterns[45965] = 29'b1_011001110001_101_0_110110011100;
      patterns[45966] = 29'b1_011001110001_110_1_011001110001;
      patterns[45967] = 29'b1_011001110001_111_1_011001110001;
      patterns[45968] = 29'b1_011001110010_000_1_011001110010;
      patterns[45969] = 29'b1_011001110010_001_1_110010011001;
      patterns[45970] = 29'b1_011001110010_010_0_110011100101;
      patterns[45971] = 29'b1_011001110010_011_1_100111001010;
      patterns[45972] = 29'b1_011001110010_100_0_101100111001;
      patterns[45973] = 29'b1_011001110010_101_1_010110011100;
      patterns[45974] = 29'b1_011001110010_110_1_011001110010;
      patterns[45975] = 29'b1_011001110010_111_1_011001110010;
      patterns[45976] = 29'b1_011001110011_000_1_011001110011;
      patterns[45977] = 29'b1_011001110011_001_1_110011011001;
      patterns[45978] = 29'b1_011001110011_010_0_110011100111;
      patterns[45979] = 29'b1_011001110011_011_1_100111001110;
      patterns[45980] = 29'b1_011001110011_100_1_101100111001;
      patterns[45981] = 29'b1_011001110011_101_1_110110011100;
      patterns[45982] = 29'b1_011001110011_110_1_011001110011;
      patterns[45983] = 29'b1_011001110011_111_1_011001110011;
      patterns[45984] = 29'b1_011001110100_000_1_011001110100;
      patterns[45985] = 29'b1_011001110100_001_1_110100011001;
      patterns[45986] = 29'b1_011001110100_010_0_110011101001;
      patterns[45987] = 29'b1_011001110100_011_1_100111010010;
      patterns[45988] = 29'b1_011001110100_100_0_101100111010;
      patterns[45989] = 29'b1_011001110100_101_0_010110011101;
      patterns[45990] = 29'b1_011001110100_110_1_011001110100;
      patterns[45991] = 29'b1_011001110100_111_1_011001110100;
      patterns[45992] = 29'b1_011001110101_000_1_011001110101;
      patterns[45993] = 29'b1_011001110101_001_1_110101011001;
      patterns[45994] = 29'b1_011001110101_010_0_110011101011;
      patterns[45995] = 29'b1_011001110101_011_1_100111010110;
      patterns[45996] = 29'b1_011001110101_100_1_101100111010;
      patterns[45997] = 29'b1_011001110101_101_0_110110011101;
      patterns[45998] = 29'b1_011001110101_110_1_011001110101;
      patterns[45999] = 29'b1_011001110101_111_1_011001110101;
      patterns[46000] = 29'b1_011001110110_000_1_011001110110;
      patterns[46001] = 29'b1_011001110110_001_1_110110011001;
      patterns[46002] = 29'b1_011001110110_010_0_110011101101;
      patterns[46003] = 29'b1_011001110110_011_1_100111011010;
      patterns[46004] = 29'b1_011001110110_100_0_101100111011;
      patterns[46005] = 29'b1_011001110110_101_1_010110011101;
      patterns[46006] = 29'b1_011001110110_110_1_011001110110;
      patterns[46007] = 29'b1_011001110110_111_1_011001110110;
      patterns[46008] = 29'b1_011001110111_000_1_011001110111;
      patterns[46009] = 29'b1_011001110111_001_1_110111011001;
      patterns[46010] = 29'b1_011001110111_010_0_110011101111;
      patterns[46011] = 29'b1_011001110111_011_1_100111011110;
      patterns[46012] = 29'b1_011001110111_100_1_101100111011;
      patterns[46013] = 29'b1_011001110111_101_1_110110011101;
      patterns[46014] = 29'b1_011001110111_110_1_011001110111;
      patterns[46015] = 29'b1_011001110111_111_1_011001110111;
      patterns[46016] = 29'b1_011001111000_000_1_011001111000;
      patterns[46017] = 29'b1_011001111000_001_1_111000011001;
      patterns[46018] = 29'b1_011001111000_010_0_110011110001;
      patterns[46019] = 29'b1_011001111000_011_1_100111100010;
      patterns[46020] = 29'b1_011001111000_100_0_101100111100;
      patterns[46021] = 29'b1_011001111000_101_0_010110011110;
      patterns[46022] = 29'b1_011001111000_110_1_011001111000;
      patterns[46023] = 29'b1_011001111000_111_1_011001111000;
      patterns[46024] = 29'b1_011001111001_000_1_011001111001;
      patterns[46025] = 29'b1_011001111001_001_1_111001011001;
      patterns[46026] = 29'b1_011001111001_010_0_110011110011;
      patterns[46027] = 29'b1_011001111001_011_1_100111100110;
      patterns[46028] = 29'b1_011001111001_100_1_101100111100;
      patterns[46029] = 29'b1_011001111001_101_0_110110011110;
      patterns[46030] = 29'b1_011001111001_110_1_011001111001;
      patterns[46031] = 29'b1_011001111001_111_1_011001111001;
      patterns[46032] = 29'b1_011001111010_000_1_011001111010;
      patterns[46033] = 29'b1_011001111010_001_1_111010011001;
      patterns[46034] = 29'b1_011001111010_010_0_110011110101;
      patterns[46035] = 29'b1_011001111010_011_1_100111101010;
      patterns[46036] = 29'b1_011001111010_100_0_101100111101;
      patterns[46037] = 29'b1_011001111010_101_1_010110011110;
      patterns[46038] = 29'b1_011001111010_110_1_011001111010;
      patterns[46039] = 29'b1_011001111010_111_1_011001111010;
      patterns[46040] = 29'b1_011001111011_000_1_011001111011;
      patterns[46041] = 29'b1_011001111011_001_1_111011011001;
      patterns[46042] = 29'b1_011001111011_010_0_110011110111;
      patterns[46043] = 29'b1_011001111011_011_1_100111101110;
      patterns[46044] = 29'b1_011001111011_100_1_101100111101;
      patterns[46045] = 29'b1_011001111011_101_1_110110011110;
      patterns[46046] = 29'b1_011001111011_110_1_011001111011;
      patterns[46047] = 29'b1_011001111011_111_1_011001111011;
      patterns[46048] = 29'b1_011001111100_000_1_011001111100;
      patterns[46049] = 29'b1_011001111100_001_1_111100011001;
      patterns[46050] = 29'b1_011001111100_010_0_110011111001;
      patterns[46051] = 29'b1_011001111100_011_1_100111110010;
      patterns[46052] = 29'b1_011001111100_100_0_101100111110;
      patterns[46053] = 29'b1_011001111100_101_0_010110011111;
      patterns[46054] = 29'b1_011001111100_110_1_011001111100;
      patterns[46055] = 29'b1_011001111100_111_1_011001111100;
      patterns[46056] = 29'b1_011001111101_000_1_011001111101;
      patterns[46057] = 29'b1_011001111101_001_1_111101011001;
      patterns[46058] = 29'b1_011001111101_010_0_110011111011;
      patterns[46059] = 29'b1_011001111101_011_1_100111110110;
      patterns[46060] = 29'b1_011001111101_100_1_101100111110;
      patterns[46061] = 29'b1_011001111101_101_0_110110011111;
      patterns[46062] = 29'b1_011001111101_110_1_011001111101;
      patterns[46063] = 29'b1_011001111101_111_1_011001111101;
      patterns[46064] = 29'b1_011001111110_000_1_011001111110;
      patterns[46065] = 29'b1_011001111110_001_1_111110011001;
      patterns[46066] = 29'b1_011001111110_010_0_110011111101;
      patterns[46067] = 29'b1_011001111110_011_1_100111111010;
      patterns[46068] = 29'b1_011001111110_100_0_101100111111;
      patterns[46069] = 29'b1_011001111110_101_1_010110011111;
      patterns[46070] = 29'b1_011001111110_110_1_011001111110;
      patterns[46071] = 29'b1_011001111110_111_1_011001111110;
      patterns[46072] = 29'b1_011001111111_000_1_011001111111;
      patterns[46073] = 29'b1_011001111111_001_1_111111011001;
      patterns[46074] = 29'b1_011001111111_010_0_110011111111;
      patterns[46075] = 29'b1_011001111111_011_1_100111111110;
      patterns[46076] = 29'b1_011001111111_100_1_101100111111;
      patterns[46077] = 29'b1_011001111111_101_1_110110011111;
      patterns[46078] = 29'b1_011001111111_110_1_011001111111;
      patterns[46079] = 29'b1_011001111111_111_1_011001111111;
      patterns[46080] = 29'b1_011010000000_000_1_011010000000;
      patterns[46081] = 29'b1_011010000000_001_1_000000011010;
      patterns[46082] = 29'b1_011010000000_010_0_110100000001;
      patterns[46083] = 29'b1_011010000000_011_1_101000000010;
      patterns[46084] = 29'b1_011010000000_100_0_101101000000;
      patterns[46085] = 29'b1_011010000000_101_0_010110100000;
      patterns[46086] = 29'b1_011010000000_110_1_011010000000;
      patterns[46087] = 29'b1_011010000000_111_1_011010000000;
      patterns[46088] = 29'b1_011010000001_000_1_011010000001;
      patterns[46089] = 29'b1_011010000001_001_1_000001011010;
      patterns[46090] = 29'b1_011010000001_010_0_110100000011;
      patterns[46091] = 29'b1_011010000001_011_1_101000000110;
      patterns[46092] = 29'b1_011010000001_100_1_101101000000;
      patterns[46093] = 29'b1_011010000001_101_0_110110100000;
      patterns[46094] = 29'b1_011010000001_110_1_011010000001;
      patterns[46095] = 29'b1_011010000001_111_1_011010000001;
      patterns[46096] = 29'b1_011010000010_000_1_011010000010;
      patterns[46097] = 29'b1_011010000010_001_1_000010011010;
      patterns[46098] = 29'b1_011010000010_010_0_110100000101;
      patterns[46099] = 29'b1_011010000010_011_1_101000001010;
      patterns[46100] = 29'b1_011010000010_100_0_101101000001;
      patterns[46101] = 29'b1_011010000010_101_1_010110100000;
      patterns[46102] = 29'b1_011010000010_110_1_011010000010;
      patterns[46103] = 29'b1_011010000010_111_1_011010000010;
      patterns[46104] = 29'b1_011010000011_000_1_011010000011;
      patterns[46105] = 29'b1_011010000011_001_1_000011011010;
      patterns[46106] = 29'b1_011010000011_010_0_110100000111;
      patterns[46107] = 29'b1_011010000011_011_1_101000001110;
      patterns[46108] = 29'b1_011010000011_100_1_101101000001;
      patterns[46109] = 29'b1_011010000011_101_1_110110100000;
      patterns[46110] = 29'b1_011010000011_110_1_011010000011;
      patterns[46111] = 29'b1_011010000011_111_1_011010000011;
      patterns[46112] = 29'b1_011010000100_000_1_011010000100;
      patterns[46113] = 29'b1_011010000100_001_1_000100011010;
      patterns[46114] = 29'b1_011010000100_010_0_110100001001;
      patterns[46115] = 29'b1_011010000100_011_1_101000010010;
      patterns[46116] = 29'b1_011010000100_100_0_101101000010;
      patterns[46117] = 29'b1_011010000100_101_0_010110100001;
      patterns[46118] = 29'b1_011010000100_110_1_011010000100;
      patterns[46119] = 29'b1_011010000100_111_1_011010000100;
      patterns[46120] = 29'b1_011010000101_000_1_011010000101;
      patterns[46121] = 29'b1_011010000101_001_1_000101011010;
      patterns[46122] = 29'b1_011010000101_010_0_110100001011;
      patterns[46123] = 29'b1_011010000101_011_1_101000010110;
      patterns[46124] = 29'b1_011010000101_100_1_101101000010;
      patterns[46125] = 29'b1_011010000101_101_0_110110100001;
      patterns[46126] = 29'b1_011010000101_110_1_011010000101;
      patterns[46127] = 29'b1_011010000101_111_1_011010000101;
      patterns[46128] = 29'b1_011010000110_000_1_011010000110;
      patterns[46129] = 29'b1_011010000110_001_1_000110011010;
      patterns[46130] = 29'b1_011010000110_010_0_110100001101;
      patterns[46131] = 29'b1_011010000110_011_1_101000011010;
      patterns[46132] = 29'b1_011010000110_100_0_101101000011;
      patterns[46133] = 29'b1_011010000110_101_1_010110100001;
      patterns[46134] = 29'b1_011010000110_110_1_011010000110;
      patterns[46135] = 29'b1_011010000110_111_1_011010000110;
      patterns[46136] = 29'b1_011010000111_000_1_011010000111;
      patterns[46137] = 29'b1_011010000111_001_1_000111011010;
      patterns[46138] = 29'b1_011010000111_010_0_110100001111;
      patterns[46139] = 29'b1_011010000111_011_1_101000011110;
      patterns[46140] = 29'b1_011010000111_100_1_101101000011;
      patterns[46141] = 29'b1_011010000111_101_1_110110100001;
      patterns[46142] = 29'b1_011010000111_110_1_011010000111;
      patterns[46143] = 29'b1_011010000111_111_1_011010000111;
      patterns[46144] = 29'b1_011010001000_000_1_011010001000;
      patterns[46145] = 29'b1_011010001000_001_1_001000011010;
      patterns[46146] = 29'b1_011010001000_010_0_110100010001;
      patterns[46147] = 29'b1_011010001000_011_1_101000100010;
      patterns[46148] = 29'b1_011010001000_100_0_101101000100;
      patterns[46149] = 29'b1_011010001000_101_0_010110100010;
      patterns[46150] = 29'b1_011010001000_110_1_011010001000;
      patterns[46151] = 29'b1_011010001000_111_1_011010001000;
      patterns[46152] = 29'b1_011010001001_000_1_011010001001;
      patterns[46153] = 29'b1_011010001001_001_1_001001011010;
      patterns[46154] = 29'b1_011010001001_010_0_110100010011;
      patterns[46155] = 29'b1_011010001001_011_1_101000100110;
      patterns[46156] = 29'b1_011010001001_100_1_101101000100;
      patterns[46157] = 29'b1_011010001001_101_0_110110100010;
      patterns[46158] = 29'b1_011010001001_110_1_011010001001;
      patterns[46159] = 29'b1_011010001001_111_1_011010001001;
      patterns[46160] = 29'b1_011010001010_000_1_011010001010;
      patterns[46161] = 29'b1_011010001010_001_1_001010011010;
      patterns[46162] = 29'b1_011010001010_010_0_110100010101;
      patterns[46163] = 29'b1_011010001010_011_1_101000101010;
      patterns[46164] = 29'b1_011010001010_100_0_101101000101;
      patterns[46165] = 29'b1_011010001010_101_1_010110100010;
      patterns[46166] = 29'b1_011010001010_110_1_011010001010;
      patterns[46167] = 29'b1_011010001010_111_1_011010001010;
      patterns[46168] = 29'b1_011010001011_000_1_011010001011;
      patterns[46169] = 29'b1_011010001011_001_1_001011011010;
      patterns[46170] = 29'b1_011010001011_010_0_110100010111;
      patterns[46171] = 29'b1_011010001011_011_1_101000101110;
      patterns[46172] = 29'b1_011010001011_100_1_101101000101;
      patterns[46173] = 29'b1_011010001011_101_1_110110100010;
      patterns[46174] = 29'b1_011010001011_110_1_011010001011;
      patterns[46175] = 29'b1_011010001011_111_1_011010001011;
      patterns[46176] = 29'b1_011010001100_000_1_011010001100;
      patterns[46177] = 29'b1_011010001100_001_1_001100011010;
      patterns[46178] = 29'b1_011010001100_010_0_110100011001;
      patterns[46179] = 29'b1_011010001100_011_1_101000110010;
      patterns[46180] = 29'b1_011010001100_100_0_101101000110;
      patterns[46181] = 29'b1_011010001100_101_0_010110100011;
      patterns[46182] = 29'b1_011010001100_110_1_011010001100;
      patterns[46183] = 29'b1_011010001100_111_1_011010001100;
      patterns[46184] = 29'b1_011010001101_000_1_011010001101;
      patterns[46185] = 29'b1_011010001101_001_1_001101011010;
      patterns[46186] = 29'b1_011010001101_010_0_110100011011;
      patterns[46187] = 29'b1_011010001101_011_1_101000110110;
      patterns[46188] = 29'b1_011010001101_100_1_101101000110;
      patterns[46189] = 29'b1_011010001101_101_0_110110100011;
      patterns[46190] = 29'b1_011010001101_110_1_011010001101;
      patterns[46191] = 29'b1_011010001101_111_1_011010001101;
      patterns[46192] = 29'b1_011010001110_000_1_011010001110;
      patterns[46193] = 29'b1_011010001110_001_1_001110011010;
      patterns[46194] = 29'b1_011010001110_010_0_110100011101;
      patterns[46195] = 29'b1_011010001110_011_1_101000111010;
      patterns[46196] = 29'b1_011010001110_100_0_101101000111;
      patterns[46197] = 29'b1_011010001110_101_1_010110100011;
      patterns[46198] = 29'b1_011010001110_110_1_011010001110;
      patterns[46199] = 29'b1_011010001110_111_1_011010001110;
      patterns[46200] = 29'b1_011010001111_000_1_011010001111;
      patterns[46201] = 29'b1_011010001111_001_1_001111011010;
      patterns[46202] = 29'b1_011010001111_010_0_110100011111;
      patterns[46203] = 29'b1_011010001111_011_1_101000111110;
      patterns[46204] = 29'b1_011010001111_100_1_101101000111;
      patterns[46205] = 29'b1_011010001111_101_1_110110100011;
      patterns[46206] = 29'b1_011010001111_110_1_011010001111;
      patterns[46207] = 29'b1_011010001111_111_1_011010001111;
      patterns[46208] = 29'b1_011010010000_000_1_011010010000;
      patterns[46209] = 29'b1_011010010000_001_1_010000011010;
      patterns[46210] = 29'b1_011010010000_010_0_110100100001;
      patterns[46211] = 29'b1_011010010000_011_1_101001000010;
      patterns[46212] = 29'b1_011010010000_100_0_101101001000;
      patterns[46213] = 29'b1_011010010000_101_0_010110100100;
      patterns[46214] = 29'b1_011010010000_110_1_011010010000;
      patterns[46215] = 29'b1_011010010000_111_1_011010010000;
      patterns[46216] = 29'b1_011010010001_000_1_011010010001;
      patterns[46217] = 29'b1_011010010001_001_1_010001011010;
      patterns[46218] = 29'b1_011010010001_010_0_110100100011;
      patterns[46219] = 29'b1_011010010001_011_1_101001000110;
      patterns[46220] = 29'b1_011010010001_100_1_101101001000;
      patterns[46221] = 29'b1_011010010001_101_0_110110100100;
      patterns[46222] = 29'b1_011010010001_110_1_011010010001;
      patterns[46223] = 29'b1_011010010001_111_1_011010010001;
      patterns[46224] = 29'b1_011010010010_000_1_011010010010;
      patterns[46225] = 29'b1_011010010010_001_1_010010011010;
      patterns[46226] = 29'b1_011010010010_010_0_110100100101;
      patterns[46227] = 29'b1_011010010010_011_1_101001001010;
      patterns[46228] = 29'b1_011010010010_100_0_101101001001;
      patterns[46229] = 29'b1_011010010010_101_1_010110100100;
      patterns[46230] = 29'b1_011010010010_110_1_011010010010;
      patterns[46231] = 29'b1_011010010010_111_1_011010010010;
      patterns[46232] = 29'b1_011010010011_000_1_011010010011;
      patterns[46233] = 29'b1_011010010011_001_1_010011011010;
      patterns[46234] = 29'b1_011010010011_010_0_110100100111;
      patterns[46235] = 29'b1_011010010011_011_1_101001001110;
      patterns[46236] = 29'b1_011010010011_100_1_101101001001;
      patterns[46237] = 29'b1_011010010011_101_1_110110100100;
      patterns[46238] = 29'b1_011010010011_110_1_011010010011;
      patterns[46239] = 29'b1_011010010011_111_1_011010010011;
      patterns[46240] = 29'b1_011010010100_000_1_011010010100;
      patterns[46241] = 29'b1_011010010100_001_1_010100011010;
      patterns[46242] = 29'b1_011010010100_010_0_110100101001;
      patterns[46243] = 29'b1_011010010100_011_1_101001010010;
      patterns[46244] = 29'b1_011010010100_100_0_101101001010;
      patterns[46245] = 29'b1_011010010100_101_0_010110100101;
      patterns[46246] = 29'b1_011010010100_110_1_011010010100;
      patterns[46247] = 29'b1_011010010100_111_1_011010010100;
      patterns[46248] = 29'b1_011010010101_000_1_011010010101;
      patterns[46249] = 29'b1_011010010101_001_1_010101011010;
      patterns[46250] = 29'b1_011010010101_010_0_110100101011;
      patterns[46251] = 29'b1_011010010101_011_1_101001010110;
      patterns[46252] = 29'b1_011010010101_100_1_101101001010;
      patterns[46253] = 29'b1_011010010101_101_0_110110100101;
      patterns[46254] = 29'b1_011010010101_110_1_011010010101;
      patterns[46255] = 29'b1_011010010101_111_1_011010010101;
      patterns[46256] = 29'b1_011010010110_000_1_011010010110;
      patterns[46257] = 29'b1_011010010110_001_1_010110011010;
      patterns[46258] = 29'b1_011010010110_010_0_110100101101;
      patterns[46259] = 29'b1_011010010110_011_1_101001011010;
      patterns[46260] = 29'b1_011010010110_100_0_101101001011;
      patterns[46261] = 29'b1_011010010110_101_1_010110100101;
      patterns[46262] = 29'b1_011010010110_110_1_011010010110;
      patterns[46263] = 29'b1_011010010110_111_1_011010010110;
      patterns[46264] = 29'b1_011010010111_000_1_011010010111;
      patterns[46265] = 29'b1_011010010111_001_1_010111011010;
      patterns[46266] = 29'b1_011010010111_010_0_110100101111;
      patterns[46267] = 29'b1_011010010111_011_1_101001011110;
      patterns[46268] = 29'b1_011010010111_100_1_101101001011;
      patterns[46269] = 29'b1_011010010111_101_1_110110100101;
      patterns[46270] = 29'b1_011010010111_110_1_011010010111;
      patterns[46271] = 29'b1_011010010111_111_1_011010010111;
      patterns[46272] = 29'b1_011010011000_000_1_011010011000;
      patterns[46273] = 29'b1_011010011000_001_1_011000011010;
      patterns[46274] = 29'b1_011010011000_010_0_110100110001;
      patterns[46275] = 29'b1_011010011000_011_1_101001100010;
      patterns[46276] = 29'b1_011010011000_100_0_101101001100;
      patterns[46277] = 29'b1_011010011000_101_0_010110100110;
      patterns[46278] = 29'b1_011010011000_110_1_011010011000;
      patterns[46279] = 29'b1_011010011000_111_1_011010011000;
      patterns[46280] = 29'b1_011010011001_000_1_011010011001;
      patterns[46281] = 29'b1_011010011001_001_1_011001011010;
      patterns[46282] = 29'b1_011010011001_010_0_110100110011;
      patterns[46283] = 29'b1_011010011001_011_1_101001100110;
      patterns[46284] = 29'b1_011010011001_100_1_101101001100;
      patterns[46285] = 29'b1_011010011001_101_0_110110100110;
      patterns[46286] = 29'b1_011010011001_110_1_011010011001;
      patterns[46287] = 29'b1_011010011001_111_1_011010011001;
      patterns[46288] = 29'b1_011010011010_000_1_011010011010;
      patterns[46289] = 29'b1_011010011010_001_1_011010011010;
      patterns[46290] = 29'b1_011010011010_010_0_110100110101;
      patterns[46291] = 29'b1_011010011010_011_1_101001101010;
      patterns[46292] = 29'b1_011010011010_100_0_101101001101;
      patterns[46293] = 29'b1_011010011010_101_1_010110100110;
      patterns[46294] = 29'b1_011010011010_110_1_011010011010;
      patterns[46295] = 29'b1_011010011010_111_1_011010011010;
      patterns[46296] = 29'b1_011010011011_000_1_011010011011;
      patterns[46297] = 29'b1_011010011011_001_1_011011011010;
      patterns[46298] = 29'b1_011010011011_010_0_110100110111;
      patterns[46299] = 29'b1_011010011011_011_1_101001101110;
      patterns[46300] = 29'b1_011010011011_100_1_101101001101;
      patterns[46301] = 29'b1_011010011011_101_1_110110100110;
      patterns[46302] = 29'b1_011010011011_110_1_011010011011;
      patterns[46303] = 29'b1_011010011011_111_1_011010011011;
      patterns[46304] = 29'b1_011010011100_000_1_011010011100;
      patterns[46305] = 29'b1_011010011100_001_1_011100011010;
      patterns[46306] = 29'b1_011010011100_010_0_110100111001;
      patterns[46307] = 29'b1_011010011100_011_1_101001110010;
      patterns[46308] = 29'b1_011010011100_100_0_101101001110;
      patterns[46309] = 29'b1_011010011100_101_0_010110100111;
      patterns[46310] = 29'b1_011010011100_110_1_011010011100;
      patterns[46311] = 29'b1_011010011100_111_1_011010011100;
      patterns[46312] = 29'b1_011010011101_000_1_011010011101;
      patterns[46313] = 29'b1_011010011101_001_1_011101011010;
      patterns[46314] = 29'b1_011010011101_010_0_110100111011;
      patterns[46315] = 29'b1_011010011101_011_1_101001110110;
      patterns[46316] = 29'b1_011010011101_100_1_101101001110;
      patterns[46317] = 29'b1_011010011101_101_0_110110100111;
      patterns[46318] = 29'b1_011010011101_110_1_011010011101;
      patterns[46319] = 29'b1_011010011101_111_1_011010011101;
      patterns[46320] = 29'b1_011010011110_000_1_011010011110;
      patterns[46321] = 29'b1_011010011110_001_1_011110011010;
      patterns[46322] = 29'b1_011010011110_010_0_110100111101;
      patterns[46323] = 29'b1_011010011110_011_1_101001111010;
      patterns[46324] = 29'b1_011010011110_100_0_101101001111;
      patterns[46325] = 29'b1_011010011110_101_1_010110100111;
      patterns[46326] = 29'b1_011010011110_110_1_011010011110;
      patterns[46327] = 29'b1_011010011110_111_1_011010011110;
      patterns[46328] = 29'b1_011010011111_000_1_011010011111;
      patterns[46329] = 29'b1_011010011111_001_1_011111011010;
      patterns[46330] = 29'b1_011010011111_010_0_110100111111;
      patterns[46331] = 29'b1_011010011111_011_1_101001111110;
      patterns[46332] = 29'b1_011010011111_100_1_101101001111;
      patterns[46333] = 29'b1_011010011111_101_1_110110100111;
      patterns[46334] = 29'b1_011010011111_110_1_011010011111;
      patterns[46335] = 29'b1_011010011111_111_1_011010011111;
      patterns[46336] = 29'b1_011010100000_000_1_011010100000;
      patterns[46337] = 29'b1_011010100000_001_1_100000011010;
      patterns[46338] = 29'b1_011010100000_010_0_110101000001;
      patterns[46339] = 29'b1_011010100000_011_1_101010000010;
      patterns[46340] = 29'b1_011010100000_100_0_101101010000;
      patterns[46341] = 29'b1_011010100000_101_0_010110101000;
      patterns[46342] = 29'b1_011010100000_110_1_011010100000;
      patterns[46343] = 29'b1_011010100000_111_1_011010100000;
      patterns[46344] = 29'b1_011010100001_000_1_011010100001;
      patterns[46345] = 29'b1_011010100001_001_1_100001011010;
      patterns[46346] = 29'b1_011010100001_010_0_110101000011;
      patterns[46347] = 29'b1_011010100001_011_1_101010000110;
      patterns[46348] = 29'b1_011010100001_100_1_101101010000;
      patterns[46349] = 29'b1_011010100001_101_0_110110101000;
      patterns[46350] = 29'b1_011010100001_110_1_011010100001;
      patterns[46351] = 29'b1_011010100001_111_1_011010100001;
      patterns[46352] = 29'b1_011010100010_000_1_011010100010;
      patterns[46353] = 29'b1_011010100010_001_1_100010011010;
      patterns[46354] = 29'b1_011010100010_010_0_110101000101;
      patterns[46355] = 29'b1_011010100010_011_1_101010001010;
      patterns[46356] = 29'b1_011010100010_100_0_101101010001;
      patterns[46357] = 29'b1_011010100010_101_1_010110101000;
      patterns[46358] = 29'b1_011010100010_110_1_011010100010;
      patterns[46359] = 29'b1_011010100010_111_1_011010100010;
      patterns[46360] = 29'b1_011010100011_000_1_011010100011;
      patterns[46361] = 29'b1_011010100011_001_1_100011011010;
      patterns[46362] = 29'b1_011010100011_010_0_110101000111;
      patterns[46363] = 29'b1_011010100011_011_1_101010001110;
      patterns[46364] = 29'b1_011010100011_100_1_101101010001;
      patterns[46365] = 29'b1_011010100011_101_1_110110101000;
      patterns[46366] = 29'b1_011010100011_110_1_011010100011;
      patterns[46367] = 29'b1_011010100011_111_1_011010100011;
      patterns[46368] = 29'b1_011010100100_000_1_011010100100;
      patterns[46369] = 29'b1_011010100100_001_1_100100011010;
      patterns[46370] = 29'b1_011010100100_010_0_110101001001;
      patterns[46371] = 29'b1_011010100100_011_1_101010010010;
      patterns[46372] = 29'b1_011010100100_100_0_101101010010;
      patterns[46373] = 29'b1_011010100100_101_0_010110101001;
      patterns[46374] = 29'b1_011010100100_110_1_011010100100;
      patterns[46375] = 29'b1_011010100100_111_1_011010100100;
      patterns[46376] = 29'b1_011010100101_000_1_011010100101;
      patterns[46377] = 29'b1_011010100101_001_1_100101011010;
      patterns[46378] = 29'b1_011010100101_010_0_110101001011;
      patterns[46379] = 29'b1_011010100101_011_1_101010010110;
      patterns[46380] = 29'b1_011010100101_100_1_101101010010;
      patterns[46381] = 29'b1_011010100101_101_0_110110101001;
      patterns[46382] = 29'b1_011010100101_110_1_011010100101;
      patterns[46383] = 29'b1_011010100101_111_1_011010100101;
      patterns[46384] = 29'b1_011010100110_000_1_011010100110;
      patterns[46385] = 29'b1_011010100110_001_1_100110011010;
      patterns[46386] = 29'b1_011010100110_010_0_110101001101;
      patterns[46387] = 29'b1_011010100110_011_1_101010011010;
      patterns[46388] = 29'b1_011010100110_100_0_101101010011;
      patterns[46389] = 29'b1_011010100110_101_1_010110101001;
      patterns[46390] = 29'b1_011010100110_110_1_011010100110;
      patterns[46391] = 29'b1_011010100110_111_1_011010100110;
      patterns[46392] = 29'b1_011010100111_000_1_011010100111;
      patterns[46393] = 29'b1_011010100111_001_1_100111011010;
      patterns[46394] = 29'b1_011010100111_010_0_110101001111;
      patterns[46395] = 29'b1_011010100111_011_1_101010011110;
      patterns[46396] = 29'b1_011010100111_100_1_101101010011;
      patterns[46397] = 29'b1_011010100111_101_1_110110101001;
      patterns[46398] = 29'b1_011010100111_110_1_011010100111;
      patterns[46399] = 29'b1_011010100111_111_1_011010100111;
      patterns[46400] = 29'b1_011010101000_000_1_011010101000;
      patterns[46401] = 29'b1_011010101000_001_1_101000011010;
      patterns[46402] = 29'b1_011010101000_010_0_110101010001;
      patterns[46403] = 29'b1_011010101000_011_1_101010100010;
      patterns[46404] = 29'b1_011010101000_100_0_101101010100;
      patterns[46405] = 29'b1_011010101000_101_0_010110101010;
      patterns[46406] = 29'b1_011010101000_110_1_011010101000;
      patterns[46407] = 29'b1_011010101000_111_1_011010101000;
      patterns[46408] = 29'b1_011010101001_000_1_011010101001;
      patterns[46409] = 29'b1_011010101001_001_1_101001011010;
      patterns[46410] = 29'b1_011010101001_010_0_110101010011;
      patterns[46411] = 29'b1_011010101001_011_1_101010100110;
      patterns[46412] = 29'b1_011010101001_100_1_101101010100;
      patterns[46413] = 29'b1_011010101001_101_0_110110101010;
      patterns[46414] = 29'b1_011010101001_110_1_011010101001;
      patterns[46415] = 29'b1_011010101001_111_1_011010101001;
      patterns[46416] = 29'b1_011010101010_000_1_011010101010;
      patterns[46417] = 29'b1_011010101010_001_1_101010011010;
      patterns[46418] = 29'b1_011010101010_010_0_110101010101;
      patterns[46419] = 29'b1_011010101010_011_1_101010101010;
      patterns[46420] = 29'b1_011010101010_100_0_101101010101;
      patterns[46421] = 29'b1_011010101010_101_1_010110101010;
      patterns[46422] = 29'b1_011010101010_110_1_011010101010;
      patterns[46423] = 29'b1_011010101010_111_1_011010101010;
      patterns[46424] = 29'b1_011010101011_000_1_011010101011;
      patterns[46425] = 29'b1_011010101011_001_1_101011011010;
      patterns[46426] = 29'b1_011010101011_010_0_110101010111;
      patterns[46427] = 29'b1_011010101011_011_1_101010101110;
      patterns[46428] = 29'b1_011010101011_100_1_101101010101;
      patterns[46429] = 29'b1_011010101011_101_1_110110101010;
      patterns[46430] = 29'b1_011010101011_110_1_011010101011;
      patterns[46431] = 29'b1_011010101011_111_1_011010101011;
      patterns[46432] = 29'b1_011010101100_000_1_011010101100;
      patterns[46433] = 29'b1_011010101100_001_1_101100011010;
      patterns[46434] = 29'b1_011010101100_010_0_110101011001;
      patterns[46435] = 29'b1_011010101100_011_1_101010110010;
      patterns[46436] = 29'b1_011010101100_100_0_101101010110;
      patterns[46437] = 29'b1_011010101100_101_0_010110101011;
      patterns[46438] = 29'b1_011010101100_110_1_011010101100;
      patterns[46439] = 29'b1_011010101100_111_1_011010101100;
      patterns[46440] = 29'b1_011010101101_000_1_011010101101;
      patterns[46441] = 29'b1_011010101101_001_1_101101011010;
      patterns[46442] = 29'b1_011010101101_010_0_110101011011;
      patterns[46443] = 29'b1_011010101101_011_1_101010110110;
      patterns[46444] = 29'b1_011010101101_100_1_101101010110;
      patterns[46445] = 29'b1_011010101101_101_0_110110101011;
      patterns[46446] = 29'b1_011010101101_110_1_011010101101;
      patterns[46447] = 29'b1_011010101101_111_1_011010101101;
      patterns[46448] = 29'b1_011010101110_000_1_011010101110;
      patterns[46449] = 29'b1_011010101110_001_1_101110011010;
      patterns[46450] = 29'b1_011010101110_010_0_110101011101;
      patterns[46451] = 29'b1_011010101110_011_1_101010111010;
      patterns[46452] = 29'b1_011010101110_100_0_101101010111;
      patterns[46453] = 29'b1_011010101110_101_1_010110101011;
      patterns[46454] = 29'b1_011010101110_110_1_011010101110;
      patterns[46455] = 29'b1_011010101110_111_1_011010101110;
      patterns[46456] = 29'b1_011010101111_000_1_011010101111;
      patterns[46457] = 29'b1_011010101111_001_1_101111011010;
      patterns[46458] = 29'b1_011010101111_010_0_110101011111;
      patterns[46459] = 29'b1_011010101111_011_1_101010111110;
      patterns[46460] = 29'b1_011010101111_100_1_101101010111;
      patterns[46461] = 29'b1_011010101111_101_1_110110101011;
      patterns[46462] = 29'b1_011010101111_110_1_011010101111;
      patterns[46463] = 29'b1_011010101111_111_1_011010101111;
      patterns[46464] = 29'b1_011010110000_000_1_011010110000;
      patterns[46465] = 29'b1_011010110000_001_1_110000011010;
      patterns[46466] = 29'b1_011010110000_010_0_110101100001;
      patterns[46467] = 29'b1_011010110000_011_1_101011000010;
      patterns[46468] = 29'b1_011010110000_100_0_101101011000;
      patterns[46469] = 29'b1_011010110000_101_0_010110101100;
      patterns[46470] = 29'b1_011010110000_110_1_011010110000;
      patterns[46471] = 29'b1_011010110000_111_1_011010110000;
      patterns[46472] = 29'b1_011010110001_000_1_011010110001;
      patterns[46473] = 29'b1_011010110001_001_1_110001011010;
      patterns[46474] = 29'b1_011010110001_010_0_110101100011;
      patterns[46475] = 29'b1_011010110001_011_1_101011000110;
      patterns[46476] = 29'b1_011010110001_100_1_101101011000;
      patterns[46477] = 29'b1_011010110001_101_0_110110101100;
      patterns[46478] = 29'b1_011010110001_110_1_011010110001;
      patterns[46479] = 29'b1_011010110001_111_1_011010110001;
      patterns[46480] = 29'b1_011010110010_000_1_011010110010;
      patterns[46481] = 29'b1_011010110010_001_1_110010011010;
      patterns[46482] = 29'b1_011010110010_010_0_110101100101;
      patterns[46483] = 29'b1_011010110010_011_1_101011001010;
      patterns[46484] = 29'b1_011010110010_100_0_101101011001;
      patterns[46485] = 29'b1_011010110010_101_1_010110101100;
      patterns[46486] = 29'b1_011010110010_110_1_011010110010;
      patterns[46487] = 29'b1_011010110010_111_1_011010110010;
      patterns[46488] = 29'b1_011010110011_000_1_011010110011;
      patterns[46489] = 29'b1_011010110011_001_1_110011011010;
      patterns[46490] = 29'b1_011010110011_010_0_110101100111;
      patterns[46491] = 29'b1_011010110011_011_1_101011001110;
      patterns[46492] = 29'b1_011010110011_100_1_101101011001;
      patterns[46493] = 29'b1_011010110011_101_1_110110101100;
      patterns[46494] = 29'b1_011010110011_110_1_011010110011;
      patterns[46495] = 29'b1_011010110011_111_1_011010110011;
      patterns[46496] = 29'b1_011010110100_000_1_011010110100;
      patterns[46497] = 29'b1_011010110100_001_1_110100011010;
      patterns[46498] = 29'b1_011010110100_010_0_110101101001;
      patterns[46499] = 29'b1_011010110100_011_1_101011010010;
      patterns[46500] = 29'b1_011010110100_100_0_101101011010;
      patterns[46501] = 29'b1_011010110100_101_0_010110101101;
      patterns[46502] = 29'b1_011010110100_110_1_011010110100;
      patterns[46503] = 29'b1_011010110100_111_1_011010110100;
      patterns[46504] = 29'b1_011010110101_000_1_011010110101;
      patterns[46505] = 29'b1_011010110101_001_1_110101011010;
      patterns[46506] = 29'b1_011010110101_010_0_110101101011;
      patterns[46507] = 29'b1_011010110101_011_1_101011010110;
      patterns[46508] = 29'b1_011010110101_100_1_101101011010;
      patterns[46509] = 29'b1_011010110101_101_0_110110101101;
      patterns[46510] = 29'b1_011010110101_110_1_011010110101;
      patterns[46511] = 29'b1_011010110101_111_1_011010110101;
      patterns[46512] = 29'b1_011010110110_000_1_011010110110;
      patterns[46513] = 29'b1_011010110110_001_1_110110011010;
      patterns[46514] = 29'b1_011010110110_010_0_110101101101;
      patterns[46515] = 29'b1_011010110110_011_1_101011011010;
      patterns[46516] = 29'b1_011010110110_100_0_101101011011;
      patterns[46517] = 29'b1_011010110110_101_1_010110101101;
      patterns[46518] = 29'b1_011010110110_110_1_011010110110;
      patterns[46519] = 29'b1_011010110110_111_1_011010110110;
      patterns[46520] = 29'b1_011010110111_000_1_011010110111;
      patterns[46521] = 29'b1_011010110111_001_1_110111011010;
      patterns[46522] = 29'b1_011010110111_010_0_110101101111;
      patterns[46523] = 29'b1_011010110111_011_1_101011011110;
      patterns[46524] = 29'b1_011010110111_100_1_101101011011;
      patterns[46525] = 29'b1_011010110111_101_1_110110101101;
      patterns[46526] = 29'b1_011010110111_110_1_011010110111;
      patterns[46527] = 29'b1_011010110111_111_1_011010110111;
      patterns[46528] = 29'b1_011010111000_000_1_011010111000;
      patterns[46529] = 29'b1_011010111000_001_1_111000011010;
      patterns[46530] = 29'b1_011010111000_010_0_110101110001;
      patterns[46531] = 29'b1_011010111000_011_1_101011100010;
      patterns[46532] = 29'b1_011010111000_100_0_101101011100;
      patterns[46533] = 29'b1_011010111000_101_0_010110101110;
      patterns[46534] = 29'b1_011010111000_110_1_011010111000;
      patterns[46535] = 29'b1_011010111000_111_1_011010111000;
      patterns[46536] = 29'b1_011010111001_000_1_011010111001;
      patterns[46537] = 29'b1_011010111001_001_1_111001011010;
      patterns[46538] = 29'b1_011010111001_010_0_110101110011;
      patterns[46539] = 29'b1_011010111001_011_1_101011100110;
      patterns[46540] = 29'b1_011010111001_100_1_101101011100;
      patterns[46541] = 29'b1_011010111001_101_0_110110101110;
      patterns[46542] = 29'b1_011010111001_110_1_011010111001;
      patterns[46543] = 29'b1_011010111001_111_1_011010111001;
      patterns[46544] = 29'b1_011010111010_000_1_011010111010;
      patterns[46545] = 29'b1_011010111010_001_1_111010011010;
      patterns[46546] = 29'b1_011010111010_010_0_110101110101;
      patterns[46547] = 29'b1_011010111010_011_1_101011101010;
      patterns[46548] = 29'b1_011010111010_100_0_101101011101;
      patterns[46549] = 29'b1_011010111010_101_1_010110101110;
      patterns[46550] = 29'b1_011010111010_110_1_011010111010;
      patterns[46551] = 29'b1_011010111010_111_1_011010111010;
      patterns[46552] = 29'b1_011010111011_000_1_011010111011;
      patterns[46553] = 29'b1_011010111011_001_1_111011011010;
      patterns[46554] = 29'b1_011010111011_010_0_110101110111;
      patterns[46555] = 29'b1_011010111011_011_1_101011101110;
      patterns[46556] = 29'b1_011010111011_100_1_101101011101;
      patterns[46557] = 29'b1_011010111011_101_1_110110101110;
      patterns[46558] = 29'b1_011010111011_110_1_011010111011;
      patterns[46559] = 29'b1_011010111011_111_1_011010111011;
      patterns[46560] = 29'b1_011010111100_000_1_011010111100;
      patterns[46561] = 29'b1_011010111100_001_1_111100011010;
      patterns[46562] = 29'b1_011010111100_010_0_110101111001;
      patterns[46563] = 29'b1_011010111100_011_1_101011110010;
      patterns[46564] = 29'b1_011010111100_100_0_101101011110;
      patterns[46565] = 29'b1_011010111100_101_0_010110101111;
      patterns[46566] = 29'b1_011010111100_110_1_011010111100;
      patterns[46567] = 29'b1_011010111100_111_1_011010111100;
      patterns[46568] = 29'b1_011010111101_000_1_011010111101;
      patterns[46569] = 29'b1_011010111101_001_1_111101011010;
      patterns[46570] = 29'b1_011010111101_010_0_110101111011;
      patterns[46571] = 29'b1_011010111101_011_1_101011110110;
      patterns[46572] = 29'b1_011010111101_100_1_101101011110;
      patterns[46573] = 29'b1_011010111101_101_0_110110101111;
      patterns[46574] = 29'b1_011010111101_110_1_011010111101;
      patterns[46575] = 29'b1_011010111101_111_1_011010111101;
      patterns[46576] = 29'b1_011010111110_000_1_011010111110;
      patterns[46577] = 29'b1_011010111110_001_1_111110011010;
      patterns[46578] = 29'b1_011010111110_010_0_110101111101;
      patterns[46579] = 29'b1_011010111110_011_1_101011111010;
      patterns[46580] = 29'b1_011010111110_100_0_101101011111;
      patterns[46581] = 29'b1_011010111110_101_1_010110101111;
      patterns[46582] = 29'b1_011010111110_110_1_011010111110;
      patterns[46583] = 29'b1_011010111110_111_1_011010111110;
      patterns[46584] = 29'b1_011010111111_000_1_011010111111;
      patterns[46585] = 29'b1_011010111111_001_1_111111011010;
      patterns[46586] = 29'b1_011010111111_010_0_110101111111;
      patterns[46587] = 29'b1_011010111111_011_1_101011111110;
      patterns[46588] = 29'b1_011010111111_100_1_101101011111;
      patterns[46589] = 29'b1_011010111111_101_1_110110101111;
      patterns[46590] = 29'b1_011010111111_110_1_011010111111;
      patterns[46591] = 29'b1_011010111111_111_1_011010111111;
      patterns[46592] = 29'b1_011011000000_000_1_011011000000;
      patterns[46593] = 29'b1_011011000000_001_1_000000011011;
      patterns[46594] = 29'b1_011011000000_010_0_110110000001;
      patterns[46595] = 29'b1_011011000000_011_1_101100000010;
      patterns[46596] = 29'b1_011011000000_100_0_101101100000;
      patterns[46597] = 29'b1_011011000000_101_0_010110110000;
      patterns[46598] = 29'b1_011011000000_110_1_011011000000;
      patterns[46599] = 29'b1_011011000000_111_1_011011000000;
      patterns[46600] = 29'b1_011011000001_000_1_011011000001;
      patterns[46601] = 29'b1_011011000001_001_1_000001011011;
      patterns[46602] = 29'b1_011011000001_010_0_110110000011;
      patterns[46603] = 29'b1_011011000001_011_1_101100000110;
      patterns[46604] = 29'b1_011011000001_100_1_101101100000;
      patterns[46605] = 29'b1_011011000001_101_0_110110110000;
      patterns[46606] = 29'b1_011011000001_110_1_011011000001;
      patterns[46607] = 29'b1_011011000001_111_1_011011000001;
      patterns[46608] = 29'b1_011011000010_000_1_011011000010;
      patterns[46609] = 29'b1_011011000010_001_1_000010011011;
      patterns[46610] = 29'b1_011011000010_010_0_110110000101;
      patterns[46611] = 29'b1_011011000010_011_1_101100001010;
      patterns[46612] = 29'b1_011011000010_100_0_101101100001;
      patterns[46613] = 29'b1_011011000010_101_1_010110110000;
      patterns[46614] = 29'b1_011011000010_110_1_011011000010;
      patterns[46615] = 29'b1_011011000010_111_1_011011000010;
      patterns[46616] = 29'b1_011011000011_000_1_011011000011;
      patterns[46617] = 29'b1_011011000011_001_1_000011011011;
      patterns[46618] = 29'b1_011011000011_010_0_110110000111;
      patterns[46619] = 29'b1_011011000011_011_1_101100001110;
      patterns[46620] = 29'b1_011011000011_100_1_101101100001;
      patterns[46621] = 29'b1_011011000011_101_1_110110110000;
      patterns[46622] = 29'b1_011011000011_110_1_011011000011;
      patterns[46623] = 29'b1_011011000011_111_1_011011000011;
      patterns[46624] = 29'b1_011011000100_000_1_011011000100;
      patterns[46625] = 29'b1_011011000100_001_1_000100011011;
      patterns[46626] = 29'b1_011011000100_010_0_110110001001;
      patterns[46627] = 29'b1_011011000100_011_1_101100010010;
      patterns[46628] = 29'b1_011011000100_100_0_101101100010;
      patterns[46629] = 29'b1_011011000100_101_0_010110110001;
      patterns[46630] = 29'b1_011011000100_110_1_011011000100;
      patterns[46631] = 29'b1_011011000100_111_1_011011000100;
      patterns[46632] = 29'b1_011011000101_000_1_011011000101;
      patterns[46633] = 29'b1_011011000101_001_1_000101011011;
      patterns[46634] = 29'b1_011011000101_010_0_110110001011;
      patterns[46635] = 29'b1_011011000101_011_1_101100010110;
      patterns[46636] = 29'b1_011011000101_100_1_101101100010;
      patterns[46637] = 29'b1_011011000101_101_0_110110110001;
      patterns[46638] = 29'b1_011011000101_110_1_011011000101;
      patterns[46639] = 29'b1_011011000101_111_1_011011000101;
      patterns[46640] = 29'b1_011011000110_000_1_011011000110;
      patterns[46641] = 29'b1_011011000110_001_1_000110011011;
      patterns[46642] = 29'b1_011011000110_010_0_110110001101;
      patterns[46643] = 29'b1_011011000110_011_1_101100011010;
      patterns[46644] = 29'b1_011011000110_100_0_101101100011;
      patterns[46645] = 29'b1_011011000110_101_1_010110110001;
      patterns[46646] = 29'b1_011011000110_110_1_011011000110;
      patterns[46647] = 29'b1_011011000110_111_1_011011000110;
      patterns[46648] = 29'b1_011011000111_000_1_011011000111;
      patterns[46649] = 29'b1_011011000111_001_1_000111011011;
      patterns[46650] = 29'b1_011011000111_010_0_110110001111;
      patterns[46651] = 29'b1_011011000111_011_1_101100011110;
      patterns[46652] = 29'b1_011011000111_100_1_101101100011;
      patterns[46653] = 29'b1_011011000111_101_1_110110110001;
      patterns[46654] = 29'b1_011011000111_110_1_011011000111;
      patterns[46655] = 29'b1_011011000111_111_1_011011000111;
      patterns[46656] = 29'b1_011011001000_000_1_011011001000;
      patterns[46657] = 29'b1_011011001000_001_1_001000011011;
      patterns[46658] = 29'b1_011011001000_010_0_110110010001;
      patterns[46659] = 29'b1_011011001000_011_1_101100100010;
      patterns[46660] = 29'b1_011011001000_100_0_101101100100;
      patterns[46661] = 29'b1_011011001000_101_0_010110110010;
      patterns[46662] = 29'b1_011011001000_110_1_011011001000;
      patterns[46663] = 29'b1_011011001000_111_1_011011001000;
      patterns[46664] = 29'b1_011011001001_000_1_011011001001;
      patterns[46665] = 29'b1_011011001001_001_1_001001011011;
      patterns[46666] = 29'b1_011011001001_010_0_110110010011;
      patterns[46667] = 29'b1_011011001001_011_1_101100100110;
      patterns[46668] = 29'b1_011011001001_100_1_101101100100;
      patterns[46669] = 29'b1_011011001001_101_0_110110110010;
      patterns[46670] = 29'b1_011011001001_110_1_011011001001;
      patterns[46671] = 29'b1_011011001001_111_1_011011001001;
      patterns[46672] = 29'b1_011011001010_000_1_011011001010;
      patterns[46673] = 29'b1_011011001010_001_1_001010011011;
      patterns[46674] = 29'b1_011011001010_010_0_110110010101;
      patterns[46675] = 29'b1_011011001010_011_1_101100101010;
      patterns[46676] = 29'b1_011011001010_100_0_101101100101;
      patterns[46677] = 29'b1_011011001010_101_1_010110110010;
      patterns[46678] = 29'b1_011011001010_110_1_011011001010;
      patterns[46679] = 29'b1_011011001010_111_1_011011001010;
      patterns[46680] = 29'b1_011011001011_000_1_011011001011;
      patterns[46681] = 29'b1_011011001011_001_1_001011011011;
      patterns[46682] = 29'b1_011011001011_010_0_110110010111;
      patterns[46683] = 29'b1_011011001011_011_1_101100101110;
      patterns[46684] = 29'b1_011011001011_100_1_101101100101;
      patterns[46685] = 29'b1_011011001011_101_1_110110110010;
      patterns[46686] = 29'b1_011011001011_110_1_011011001011;
      patterns[46687] = 29'b1_011011001011_111_1_011011001011;
      patterns[46688] = 29'b1_011011001100_000_1_011011001100;
      patterns[46689] = 29'b1_011011001100_001_1_001100011011;
      patterns[46690] = 29'b1_011011001100_010_0_110110011001;
      patterns[46691] = 29'b1_011011001100_011_1_101100110010;
      patterns[46692] = 29'b1_011011001100_100_0_101101100110;
      patterns[46693] = 29'b1_011011001100_101_0_010110110011;
      patterns[46694] = 29'b1_011011001100_110_1_011011001100;
      patterns[46695] = 29'b1_011011001100_111_1_011011001100;
      patterns[46696] = 29'b1_011011001101_000_1_011011001101;
      patterns[46697] = 29'b1_011011001101_001_1_001101011011;
      patterns[46698] = 29'b1_011011001101_010_0_110110011011;
      patterns[46699] = 29'b1_011011001101_011_1_101100110110;
      patterns[46700] = 29'b1_011011001101_100_1_101101100110;
      patterns[46701] = 29'b1_011011001101_101_0_110110110011;
      patterns[46702] = 29'b1_011011001101_110_1_011011001101;
      patterns[46703] = 29'b1_011011001101_111_1_011011001101;
      patterns[46704] = 29'b1_011011001110_000_1_011011001110;
      patterns[46705] = 29'b1_011011001110_001_1_001110011011;
      patterns[46706] = 29'b1_011011001110_010_0_110110011101;
      patterns[46707] = 29'b1_011011001110_011_1_101100111010;
      patterns[46708] = 29'b1_011011001110_100_0_101101100111;
      patterns[46709] = 29'b1_011011001110_101_1_010110110011;
      patterns[46710] = 29'b1_011011001110_110_1_011011001110;
      patterns[46711] = 29'b1_011011001110_111_1_011011001110;
      patterns[46712] = 29'b1_011011001111_000_1_011011001111;
      patterns[46713] = 29'b1_011011001111_001_1_001111011011;
      patterns[46714] = 29'b1_011011001111_010_0_110110011111;
      patterns[46715] = 29'b1_011011001111_011_1_101100111110;
      patterns[46716] = 29'b1_011011001111_100_1_101101100111;
      patterns[46717] = 29'b1_011011001111_101_1_110110110011;
      patterns[46718] = 29'b1_011011001111_110_1_011011001111;
      patterns[46719] = 29'b1_011011001111_111_1_011011001111;
      patterns[46720] = 29'b1_011011010000_000_1_011011010000;
      patterns[46721] = 29'b1_011011010000_001_1_010000011011;
      patterns[46722] = 29'b1_011011010000_010_0_110110100001;
      patterns[46723] = 29'b1_011011010000_011_1_101101000010;
      patterns[46724] = 29'b1_011011010000_100_0_101101101000;
      patterns[46725] = 29'b1_011011010000_101_0_010110110100;
      patterns[46726] = 29'b1_011011010000_110_1_011011010000;
      patterns[46727] = 29'b1_011011010000_111_1_011011010000;
      patterns[46728] = 29'b1_011011010001_000_1_011011010001;
      patterns[46729] = 29'b1_011011010001_001_1_010001011011;
      patterns[46730] = 29'b1_011011010001_010_0_110110100011;
      patterns[46731] = 29'b1_011011010001_011_1_101101000110;
      patterns[46732] = 29'b1_011011010001_100_1_101101101000;
      patterns[46733] = 29'b1_011011010001_101_0_110110110100;
      patterns[46734] = 29'b1_011011010001_110_1_011011010001;
      patterns[46735] = 29'b1_011011010001_111_1_011011010001;
      patterns[46736] = 29'b1_011011010010_000_1_011011010010;
      patterns[46737] = 29'b1_011011010010_001_1_010010011011;
      patterns[46738] = 29'b1_011011010010_010_0_110110100101;
      patterns[46739] = 29'b1_011011010010_011_1_101101001010;
      patterns[46740] = 29'b1_011011010010_100_0_101101101001;
      patterns[46741] = 29'b1_011011010010_101_1_010110110100;
      patterns[46742] = 29'b1_011011010010_110_1_011011010010;
      patterns[46743] = 29'b1_011011010010_111_1_011011010010;
      patterns[46744] = 29'b1_011011010011_000_1_011011010011;
      patterns[46745] = 29'b1_011011010011_001_1_010011011011;
      patterns[46746] = 29'b1_011011010011_010_0_110110100111;
      patterns[46747] = 29'b1_011011010011_011_1_101101001110;
      patterns[46748] = 29'b1_011011010011_100_1_101101101001;
      patterns[46749] = 29'b1_011011010011_101_1_110110110100;
      patterns[46750] = 29'b1_011011010011_110_1_011011010011;
      patterns[46751] = 29'b1_011011010011_111_1_011011010011;
      patterns[46752] = 29'b1_011011010100_000_1_011011010100;
      patterns[46753] = 29'b1_011011010100_001_1_010100011011;
      patterns[46754] = 29'b1_011011010100_010_0_110110101001;
      patterns[46755] = 29'b1_011011010100_011_1_101101010010;
      patterns[46756] = 29'b1_011011010100_100_0_101101101010;
      patterns[46757] = 29'b1_011011010100_101_0_010110110101;
      patterns[46758] = 29'b1_011011010100_110_1_011011010100;
      patterns[46759] = 29'b1_011011010100_111_1_011011010100;
      patterns[46760] = 29'b1_011011010101_000_1_011011010101;
      patterns[46761] = 29'b1_011011010101_001_1_010101011011;
      patterns[46762] = 29'b1_011011010101_010_0_110110101011;
      patterns[46763] = 29'b1_011011010101_011_1_101101010110;
      patterns[46764] = 29'b1_011011010101_100_1_101101101010;
      patterns[46765] = 29'b1_011011010101_101_0_110110110101;
      patterns[46766] = 29'b1_011011010101_110_1_011011010101;
      patterns[46767] = 29'b1_011011010101_111_1_011011010101;
      patterns[46768] = 29'b1_011011010110_000_1_011011010110;
      patterns[46769] = 29'b1_011011010110_001_1_010110011011;
      patterns[46770] = 29'b1_011011010110_010_0_110110101101;
      patterns[46771] = 29'b1_011011010110_011_1_101101011010;
      patterns[46772] = 29'b1_011011010110_100_0_101101101011;
      patterns[46773] = 29'b1_011011010110_101_1_010110110101;
      patterns[46774] = 29'b1_011011010110_110_1_011011010110;
      patterns[46775] = 29'b1_011011010110_111_1_011011010110;
      patterns[46776] = 29'b1_011011010111_000_1_011011010111;
      patterns[46777] = 29'b1_011011010111_001_1_010111011011;
      patterns[46778] = 29'b1_011011010111_010_0_110110101111;
      patterns[46779] = 29'b1_011011010111_011_1_101101011110;
      patterns[46780] = 29'b1_011011010111_100_1_101101101011;
      patterns[46781] = 29'b1_011011010111_101_1_110110110101;
      patterns[46782] = 29'b1_011011010111_110_1_011011010111;
      patterns[46783] = 29'b1_011011010111_111_1_011011010111;
      patterns[46784] = 29'b1_011011011000_000_1_011011011000;
      patterns[46785] = 29'b1_011011011000_001_1_011000011011;
      patterns[46786] = 29'b1_011011011000_010_0_110110110001;
      patterns[46787] = 29'b1_011011011000_011_1_101101100010;
      patterns[46788] = 29'b1_011011011000_100_0_101101101100;
      patterns[46789] = 29'b1_011011011000_101_0_010110110110;
      patterns[46790] = 29'b1_011011011000_110_1_011011011000;
      patterns[46791] = 29'b1_011011011000_111_1_011011011000;
      patterns[46792] = 29'b1_011011011001_000_1_011011011001;
      patterns[46793] = 29'b1_011011011001_001_1_011001011011;
      patterns[46794] = 29'b1_011011011001_010_0_110110110011;
      patterns[46795] = 29'b1_011011011001_011_1_101101100110;
      patterns[46796] = 29'b1_011011011001_100_1_101101101100;
      patterns[46797] = 29'b1_011011011001_101_0_110110110110;
      patterns[46798] = 29'b1_011011011001_110_1_011011011001;
      patterns[46799] = 29'b1_011011011001_111_1_011011011001;
      patterns[46800] = 29'b1_011011011010_000_1_011011011010;
      patterns[46801] = 29'b1_011011011010_001_1_011010011011;
      patterns[46802] = 29'b1_011011011010_010_0_110110110101;
      patterns[46803] = 29'b1_011011011010_011_1_101101101010;
      patterns[46804] = 29'b1_011011011010_100_0_101101101101;
      patterns[46805] = 29'b1_011011011010_101_1_010110110110;
      patterns[46806] = 29'b1_011011011010_110_1_011011011010;
      patterns[46807] = 29'b1_011011011010_111_1_011011011010;
      patterns[46808] = 29'b1_011011011011_000_1_011011011011;
      patterns[46809] = 29'b1_011011011011_001_1_011011011011;
      patterns[46810] = 29'b1_011011011011_010_0_110110110111;
      patterns[46811] = 29'b1_011011011011_011_1_101101101110;
      patterns[46812] = 29'b1_011011011011_100_1_101101101101;
      patterns[46813] = 29'b1_011011011011_101_1_110110110110;
      patterns[46814] = 29'b1_011011011011_110_1_011011011011;
      patterns[46815] = 29'b1_011011011011_111_1_011011011011;
      patterns[46816] = 29'b1_011011011100_000_1_011011011100;
      patterns[46817] = 29'b1_011011011100_001_1_011100011011;
      patterns[46818] = 29'b1_011011011100_010_0_110110111001;
      patterns[46819] = 29'b1_011011011100_011_1_101101110010;
      patterns[46820] = 29'b1_011011011100_100_0_101101101110;
      patterns[46821] = 29'b1_011011011100_101_0_010110110111;
      patterns[46822] = 29'b1_011011011100_110_1_011011011100;
      patterns[46823] = 29'b1_011011011100_111_1_011011011100;
      patterns[46824] = 29'b1_011011011101_000_1_011011011101;
      patterns[46825] = 29'b1_011011011101_001_1_011101011011;
      patterns[46826] = 29'b1_011011011101_010_0_110110111011;
      patterns[46827] = 29'b1_011011011101_011_1_101101110110;
      patterns[46828] = 29'b1_011011011101_100_1_101101101110;
      patterns[46829] = 29'b1_011011011101_101_0_110110110111;
      patterns[46830] = 29'b1_011011011101_110_1_011011011101;
      patterns[46831] = 29'b1_011011011101_111_1_011011011101;
      patterns[46832] = 29'b1_011011011110_000_1_011011011110;
      patterns[46833] = 29'b1_011011011110_001_1_011110011011;
      patterns[46834] = 29'b1_011011011110_010_0_110110111101;
      patterns[46835] = 29'b1_011011011110_011_1_101101111010;
      patterns[46836] = 29'b1_011011011110_100_0_101101101111;
      patterns[46837] = 29'b1_011011011110_101_1_010110110111;
      patterns[46838] = 29'b1_011011011110_110_1_011011011110;
      patterns[46839] = 29'b1_011011011110_111_1_011011011110;
      patterns[46840] = 29'b1_011011011111_000_1_011011011111;
      patterns[46841] = 29'b1_011011011111_001_1_011111011011;
      patterns[46842] = 29'b1_011011011111_010_0_110110111111;
      patterns[46843] = 29'b1_011011011111_011_1_101101111110;
      patterns[46844] = 29'b1_011011011111_100_1_101101101111;
      patterns[46845] = 29'b1_011011011111_101_1_110110110111;
      patterns[46846] = 29'b1_011011011111_110_1_011011011111;
      patterns[46847] = 29'b1_011011011111_111_1_011011011111;
      patterns[46848] = 29'b1_011011100000_000_1_011011100000;
      patterns[46849] = 29'b1_011011100000_001_1_100000011011;
      patterns[46850] = 29'b1_011011100000_010_0_110111000001;
      patterns[46851] = 29'b1_011011100000_011_1_101110000010;
      patterns[46852] = 29'b1_011011100000_100_0_101101110000;
      patterns[46853] = 29'b1_011011100000_101_0_010110111000;
      patterns[46854] = 29'b1_011011100000_110_1_011011100000;
      patterns[46855] = 29'b1_011011100000_111_1_011011100000;
      patterns[46856] = 29'b1_011011100001_000_1_011011100001;
      patterns[46857] = 29'b1_011011100001_001_1_100001011011;
      patterns[46858] = 29'b1_011011100001_010_0_110111000011;
      patterns[46859] = 29'b1_011011100001_011_1_101110000110;
      patterns[46860] = 29'b1_011011100001_100_1_101101110000;
      patterns[46861] = 29'b1_011011100001_101_0_110110111000;
      patterns[46862] = 29'b1_011011100001_110_1_011011100001;
      patterns[46863] = 29'b1_011011100001_111_1_011011100001;
      patterns[46864] = 29'b1_011011100010_000_1_011011100010;
      patterns[46865] = 29'b1_011011100010_001_1_100010011011;
      patterns[46866] = 29'b1_011011100010_010_0_110111000101;
      patterns[46867] = 29'b1_011011100010_011_1_101110001010;
      patterns[46868] = 29'b1_011011100010_100_0_101101110001;
      patterns[46869] = 29'b1_011011100010_101_1_010110111000;
      patterns[46870] = 29'b1_011011100010_110_1_011011100010;
      patterns[46871] = 29'b1_011011100010_111_1_011011100010;
      patterns[46872] = 29'b1_011011100011_000_1_011011100011;
      patterns[46873] = 29'b1_011011100011_001_1_100011011011;
      patterns[46874] = 29'b1_011011100011_010_0_110111000111;
      patterns[46875] = 29'b1_011011100011_011_1_101110001110;
      patterns[46876] = 29'b1_011011100011_100_1_101101110001;
      patterns[46877] = 29'b1_011011100011_101_1_110110111000;
      patterns[46878] = 29'b1_011011100011_110_1_011011100011;
      patterns[46879] = 29'b1_011011100011_111_1_011011100011;
      patterns[46880] = 29'b1_011011100100_000_1_011011100100;
      patterns[46881] = 29'b1_011011100100_001_1_100100011011;
      patterns[46882] = 29'b1_011011100100_010_0_110111001001;
      patterns[46883] = 29'b1_011011100100_011_1_101110010010;
      patterns[46884] = 29'b1_011011100100_100_0_101101110010;
      patterns[46885] = 29'b1_011011100100_101_0_010110111001;
      patterns[46886] = 29'b1_011011100100_110_1_011011100100;
      patterns[46887] = 29'b1_011011100100_111_1_011011100100;
      patterns[46888] = 29'b1_011011100101_000_1_011011100101;
      patterns[46889] = 29'b1_011011100101_001_1_100101011011;
      patterns[46890] = 29'b1_011011100101_010_0_110111001011;
      patterns[46891] = 29'b1_011011100101_011_1_101110010110;
      patterns[46892] = 29'b1_011011100101_100_1_101101110010;
      patterns[46893] = 29'b1_011011100101_101_0_110110111001;
      patterns[46894] = 29'b1_011011100101_110_1_011011100101;
      patterns[46895] = 29'b1_011011100101_111_1_011011100101;
      patterns[46896] = 29'b1_011011100110_000_1_011011100110;
      patterns[46897] = 29'b1_011011100110_001_1_100110011011;
      patterns[46898] = 29'b1_011011100110_010_0_110111001101;
      patterns[46899] = 29'b1_011011100110_011_1_101110011010;
      patterns[46900] = 29'b1_011011100110_100_0_101101110011;
      patterns[46901] = 29'b1_011011100110_101_1_010110111001;
      patterns[46902] = 29'b1_011011100110_110_1_011011100110;
      patterns[46903] = 29'b1_011011100110_111_1_011011100110;
      patterns[46904] = 29'b1_011011100111_000_1_011011100111;
      patterns[46905] = 29'b1_011011100111_001_1_100111011011;
      patterns[46906] = 29'b1_011011100111_010_0_110111001111;
      patterns[46907] = 29'b1_011011100111_011_1_101110011110;
      patterns[46908] = 29'b1_011011100111_100_1_101101110011;
      patterns[46909] = 29'b1_011011100111_101_1_110110111001;
      patterns[46910] = 29'b1_011011100111_110_1_011011100111;
      patterns[46911] = 29'b1_011011100111_111_1_011011100111;
      patterns[46912] = 29'b1_011011101000_000_1_011011101000;
      patterns[46913] = 29'b1_011011101000_001_1_101000011011;
      patterns[46914] = 29'b1_011011101000_010_0_110111010001;
      patterns[46915] = 29'b1_011011101000_011_1_101110100010;
      patterns[46916] = 29'b1_011011101000_100_0_101101110100;
      patterns[46917] = 29'b1_011011101000_101_0_010110111010;
      patterns[46918] = 29'b1_011011101000_110_1_011011101000;
      patterns[46919] = 29'b1_011011101000_111_1_011011101000;
      patterns[46920] = 29'b1_011011101001_000_1_011011101001;
      patterns[46921] = 29'b1_011011101001_001_1_101001011011;
      patterns[46922] = 29'b1_011011101001_010_0_110111010011;
      patterns[46923] = 29'b1_011011101001_011_1_101110100110;
      patterns[46924] = 29'b1_011011101001_100_1_101101110100;
      patterns[46925] = 29'b1_011011101001_101_0_110110111010;
      patterns[46926] = 29'b1_011011101001_110_1_011011101001;
      patterns[46927] = 29'b1_011011101001_111_1_011011101001;
      patterns[46928] = 29'b1_011011101010_000_1_011011101010;
      patterns[46929] = 29'b1_011011101010_001_1_101010011011;
      patterns[46930] = 29'b1_011011101010_010_0_110111010101;
      patterns[46931] = 29'b1_011011101010_011_1_101110101010;
      patterns[46932] = 29'b1_011011101010_100_0_101101110101;
      patterns[46933] = 29'b1_011011101010_101_1_010110111010;
      patterns[46934] = 29'b1_011011101010_110_1_011011101010;
      patterns[46935] = 29'b1_011011101010_111_1_011011101010;
      patterns[46936] = 29'b1_011011101011_000_1_011011101011;
      patterns[46937] = 29'b1_011011101011_001_1_101011011011;
      patterns[46938] = 29'b1_011011101011_010_0_110111010111;
      patterns[46939] = 29'b1_011011101011_011_1_101110101110;
      patterns[46940] = 29'b1_011011101011_100_1_101101110101;
      patterns[46941] = 29'b1_011011101011_101_1_110110111010;
      patterns[46942] = 29'b1_011011101011_110_1_011011101011;
      patterns[46943] = 29'b1_011011101011_111_1_011011101011;
      patterns[46944] = 29'b1_011011101100_000_1_011011101100;
      patterns[46945] = 29'b1_011011101100_001_1_101100011011;
      patterns[46946] = 29'b1_011011101100_010_0_110111011001;
      patterns[46947] = 29'b1_011011101100_011_1_101110110010;
      patterns[46948] = 29'b1_011011101100_100_0_101101110110;
      patterns[46949] = 29'b1_011011101100_101_0_010110111011;
      patterns[46950] = 29'b1_011011101100_110_1_011011101100;
      patterns[46951] = 29'b1_011011101100_111_1_011011101100;
      patterns[46952] = 29'b1_011011101101_000_1_011011101101;
      patterns[46953] = 29'b1_011011101101_001_1_101101011011;
      patterns[46954] = 29'b1_011011101101_010_0_110111011011;
      patterns[46955] = 29'b1_011011101101_011_1_101110110110;
      patterns[46956] = 29'b1_011011101101_100_1_101101110110;
      patterns[46957] = 29'b1_011011101101_101_0_110110111011;
      patterns[46958] = 29'b1_011011101101_110_1_011011101101;
      patterns[46959] = 29'b1_011011101101_111_1_011011101101;
      patterns[46960] = 29'b1_011011101110_000_1_011011101110;
      patterns[46961] = 29'b1_011011101110_001_1_101110011011;
      patterns[46962] = 29'b1_011011101110_010_0_110111011101;
      patterns[46963] = 29'b1_011011101110_011_1_101110111010;
      patterns[46964] = 29'b1_011011101110_100_0_101101110111;
      patterns[46965] = 29'b1_011011101110_101_1_010110111011;
      patterns[46966] = 29'b1_011011101110_110_1_011011101110;
      patterns[46967] = 29'b1_011011101110_111_1_011011101110;
      patterns[46968] = 29'b1_011011101111_000_1_011011101111;
      patterns[46969] = 29'b1_011011101111_001_1_101111011011;
      patterns[46970] = 29'b1_011011101111_010_0_110111011111;
      patterns[46971] = 29'b1_011011101111_011_1_101110111110;
      patterns[46972] = 29'b1_011011101111_100_1_101101110111;
      patterns[46973] = 29'b1_011011101111_101_1_110110111011;
      patterns[46974] = 29'b1_011011101111_110_1_011011101111;
      patterns[46975] = 29'b1_011011101111_111_1_011011101111;
      patterns[46976] = 29'b1_011011110000_000_1_011011110000;
      patterns[46977] = 29'b1_011011110000_001_1_110000011011;
      patterns[46978] = 29'b1_011011110000_010_0_110111100001;
      patterns[46979] = 29'b1_011011110000_011_1_101111000010;
      patterns[46980] = 29'b1_011011110000_100_0_101101111000;
      patterns[46981] = 29'b1_011011110000_101_0_010110111100;
      patterns[46982] = 29'b1_011011110000_110_1_011011110000;
      patterns[46983] = 29'b1_011011110000_111_1_011011110000;
      patterns[46984] = 29'b1_011011110001_000_1_011011110001;
      patterns[46985] = 29'b1_011011110001_001_1_110001011011;
      patterns[46986] = 29'b1_011011110001_010_0_110111100011;
      patterns[46987] = 29'b1_011011110001_011_1_101111000110;
      patterns[46988] = 29'b1_011011110001_100_1_101101111000;
      patterns[46989] = 29'b1_011011110001_101_0_110110111100;
      patterns[46990] = 29'b1_011011110001_110_1_011011110001;
      patterns[46991] = 29'b1_011011110001_111_1_011011110001;
      patterns[46992] = 29'b1_011011110010_000_1_011011110010;
      patterns[46993] = 29'b1_011011110010_001_1_110010011011;
      patterns[46994] = 29'b1_011011110010_010_0_110111100101;
      patterns[46995] = 29'b1_011011110010_011_1_101111001010;
      patterns[46996] = 29'b1_011011110010_100_0_101101111001;
      patterns[46997] = 29'b1_011011110010_101_1_010110111100;
      patterns[46998] = 29'b1_011011110010_110_1_011011110010;
      patterns[46999] = 29'b1_011011110010_111_1_011011110010;
      patterns[47000] = 29'b1_011011110011_000_1_011011110011;
      patterns[47001] = 29'b1_011011110011_001_1_110011011011;
      patterns[47002] = 29'b1_011011110011_010_0_110111100111;
      patterns[47003] = 29'b1_011011110011_011_1_101111001110;
      patterns[47004] = 29'b1_011011110011_100_1_101101111001;
      patterns[47005] = 29'b1_011011110011_101_1_110110111100;
      patterns[47006] = 29'b1_011011110011_110_1_011011110011;
      patterns[47007] = 29'b1_011011110011_111_1_011011110011;
      patterns[47008] = 29'b1_011011110100_000_1_011011110100;
      patterns[47009] = 29'b1_011011110100_001_1_110100011011;
      patterns[47010] = 29'b1_011011110100_010_0_110111101001;
      patterns[47011] = 29'b1_011011110100_011_1_101111010010;
      patterns[47012] = 29'b1_011011110100_100_0_101101111010;
      patterns[47013] = 29'b1_011011110100_101_0_010110111101;
      patterns[47014] = 29'b1_011011110100_110_1_011011110100;
      patterns[47015] = 29'b1_011011110100_111_1_011011110100;
      patterns[47016] = 29'b1_011011110101_000_1_011011110101;
      patterns[47017] = 29'b1_011011110101_001_1_110101011011;
      patterns[47018] = 29'b1_011011110101_010_0_110111101011;
      patterns[47019] = 29'b1_011011110101_011_1_101111010110;
      patterns[47020] = 29'b1_011011110101_100_1_101101111010;
      patterns[47021] = 29'b1_011011110101_101_0_110110111101;
      patterns[47022] = 29'b1_011011110101_110_1_011011110101;
      patterns[47023] = 29'b1_011011110101_111_1_011011110101;
      patterns[47024] = 29'b1_011011110110_000_1_011011110110;
      patterns[47025] = 29'b1_011011110110_001_1_110110011011;
      patterns[47026] = 29'b1_011011110110_010_0_110111101101;
      patterns[47027] = 29'b1_011011110110_011_1_101111011010;
      patterns[47028] = 29'b1_011011110110_100_0_101101111011;
      patterns[47029] = 29'b1_011011110110_101_1_010110111101;
      patterns[47030] = 29'b1_011011110110_110_1_011011110110;
      patterns[47031] = 29'b1_011011110110_111_1_011011110110;
      patterns[47032] = 29'b1_011011110111_000_1_011011110111;
      patterns[47033] = 29'b1_011011110111_001_1_110111011011;
      patterns[47034] = 29'b1_011011110111_010_0_110111101111;
      patterns[47035] = 29'b1_011011110111_011_1_101111011110;
      patterns[47036] = 29'b1_011011110111_100_1_101101111011;
      patterns[47037] = 29'b1_011011110111_101_1_110110111101;
      patterns[47038] = 29'b1_011011110111_110_1_011011110111;
      patterns[47039] = 29'b1_011011110111_111_1_011011110111;
      patterns[47040] = 29'b1_011011111000_000_1_011011111000;
      patterns[47041] = 29'b1_011011111000_001_1_111000011011;
      patterns[47042] = 29'b1_011011111000_010_0_110111110001;
      patterns[47043] = 29'b1_011011111000_011_1_101111100010;
      patterns[47044] = 29'b1_011011111000_100_0_101101111100;
      patterns[47045] = 29'b1_011011111000_101_0_010110111110;
      patterns[47046] = 29'b1_011011111000_110_1_011011111000;
      patterns[47047] = 29'b1_011011111000_111_1_011011111000;
      patterns[47048] = 29'b1_011011111001_000_1_011011111001;
      patterns[47049] = 29'b1_011011111001_001_1_111001011011;
      patterns[47050] = 29'b1_011011111001_010_0_110111110011;
      patterns[47051] = 29'b1_011011111001_011_1_101111100110;
      patterns[47052] = 29'b1_011011111001_100_1_101101111100;
      patterns[47053] = 29'b1_011011111001_101_0_110110111110;
      patterns[47054] = 29'b1_011011111001_110_1_011011111001;
      patterns[47055] = 29'b1_011011111001_111_1_011011111001;
      patterns[47056] = 29'b1_011011111010_000_1_011011111010;
      patterns[47057] = 29'b1_011011111010_001_1_111010011011;
      patterns[47058] = 29'b1_011011111010_010_0_110111110101;
      patterns[47059] = 29'b1_011011111010_011_1_101111101010;
      patterns[47060] = 29'b1_011011111010_100_0_101101111101;
      patterns[47061] = 29'b1_011011111010_101_1_010110111110;
      patterns[47062] = 29'b1_011011111010_110_1_011011111010;
      patterns[47063] = 29'b1_011011111010_111_1_011011111010;
      patterns[47064] = 29'b1_011011111011_000_1_011011111011;
      patterns[47065] = 29'b1_011011111011_001_1_111011011011;
      patterns[47066] = 29'b1_011011111011_010_0_110111110111;
      patterns[47067] = 29'b1_011011111011_011_1_101111101110;
      patterns[47068] = 29'b1_011011111011_100_1_101101111101;
      patterns[47069] = 29'b1_011011111011_101_1_110110111110;
      patterns[47070] = 29'b1_011011111011_110_1_011011111011;
      patterns[47071] = 29'b1_011011111011_111_1_011011111011;
      patterns[47072] = 29'b1_011011111100_000_1_011011111100;
      patterns[47073] = 29'b1_011011111100_001_1_111100011011;
      patterns[47074] = 29'b1_011011111100_010_0_110111111001;
      patterns[47075] = 29'b1_011011111100_011_1_101111110010;
      patterns[47076] = 29'b1_011011111100_100_0_101101111110;
      patterns[47077] = 29'b1_011011111100_101_0_010110111111;
      patterns[47078] = 29'b1_011011111100_110_1_011011111100;
      patterns[47079] = 29'b1_011011111100_111_1_011011111100;
      patterns[47080] = 29'b1_011011111101_000_1_011011111101;
      patterns[47081] = 29'b1_011011111101_001_1_111101011011;
      patterns[47082] = 29'b1_011011111101_010_0_110111111011;
      patterns[47083] = 29'b1_011011111101_011_1_101111110110;
      patterns[47084] = 29'b1_011011111101_100_1_101101111110;
      patterns[47085] = 29'b1_011011111101_101_0_110110111111;
      patterns[47086] = 29'b1_011011111101_110_1_011011111101;
      patterns[47087] = 29'b1_011011111101_111_1_011011111101;
      patterns[47088] = 29'b1_011011111110_000_1_011011111110;
      patterns[47089] = 29'b1_011011111110_001_1_111110011011;
      patterns[47090] = 29'b1_011011111110_010_0_110111111101;
      patterns[47091] = 29'b1_011011111110_011_1_101111111010;
      patterns[47092] = 29'b1_011011111110_100_0_101101111111;
      patterns[47093] = 29'b1_011011111110_101_1_010110111111;
      patterns[47094] = 29'b1_011011111110_110_1_011011111110;
      patterns[47095] = 29'b1_011011111110_111_1_011011111110;
      patterns[47096] = 29'b1_011011111111_000_1_011011111111;
      patterns[47097] = 29'b1_011011111111_001_1_111111011011;
      patterns[47098] = 29'b1_011011111111_010_0_110111111111;
      patterns[47099] = 29'b1_011011111111_011_1_101111111110;
      patterns[47100] = 29'b1_011011111111_100_1_101101111111;
      patterns[47101] = 29'b1_011011111111_101_1_110110111111;
      patterns[47102] = 29'b1_011011111111_110_1_011011111111;
      patterns[47103] = 29'b1_011011111111_111_1_011011111111;
      patterns[47104] = 29'b1_011100000000_000_1_011100000000;
      patterns[47105] = 29'b1_011100000000_001_1_000000011100;
      patterns[47106] = 29'b1_011100000000_010_0_111000000001;
      patterns[47107] = 29'b1_011100000000_011_1_110000000010;
      patterns[47108] = 29'b1_011100000000_100_0_101110000000;
      patterns[47109] = 29'b1_011100000000_101_0_010111000000;
      patterns[47110] = 29'b1_011100000000_110_1_011100000000;
      patterns[47111] = 29'b1_011100000000_111_1_011100000000;
      patterns[47112] = 29'b1_011100000001_000_1_011100000001;
      patterns[47113] = 29'b1_011100000001_001_1_000001011100;
      patterns[47114] = 29'b1_011100000001_010_0_111000000011;
      patterns[47115] = 29'b1_011100000001_011_1_110000000110;
      patterns[47116] = 29'b1_011100000001_100_1_101110000000;
      patterns[47117] = 29'b1_011100000001_101_0_110111000000;
      patterns[47118] = 29'b1_011100000001_110_1_011100000001;
      patterns[47119] = 29'b1_011100000001_111_1_011100000001;
      patterns[47120] = 29'b1_011100000010_000_1_011100000010;
      patterns[47121] = 29'b1_011100000010_001_1_000010011100;
      patterns[47122] = 29'b1_011100000010_010_0_111000000101;
      patterns[47123] = 29'b1_011100000010_011_1_110000001010;
      patterns[47124] = 29'b1_011100000010_100_0_101110000001;
      patterns[47125] = 29'b1_011100000010_101_1_010111000000;
      patterns[47126] = 29'b1_011100000010_110_1_011100000010;
      patterns[47127] = 29'b1_011100000010_111_1_011100000010;
      patterns[47128] = 29'b1_011100000011_000_1_011100000011;
      patterns[47129] = 29'b1_011100000011_001_1_000011011100;
      patterns[47130] = 29'b1_011100000011_010_0_111000000111;
      patterns[47131] = 29'b1_011100000011_011_1_110000001110;
      patterns[47132] = 29'b1_011100000011_100_1_101110000001;
      patterns[47133] = 29'b1_011100000011_101_1_110111000000;
      patterns[47134] = 29'b1_011100000011_110_1_011100000011;
      patterns[47135] = 29'b1_011100000011_111_1_011100000011;
      patterns[47136] = 29'b1_011100000100_000_1_011100000100;
      patterns[47137] = 29'b1_011100000100_001_1_000100011100;
      patterns[47138] = 29'b1_011100000100_010_0_111000001001;
      patterns[47139] = 29'b1_011100000100_011_1_110000010010;
      patterns[47140] = 29'b1_011100000100_100_0_101110000010;
      patterns[47141] = 29'b1_011100000100_101_0_010111000001;
      patterns[47142] = 29'b1_011100000100_110_1_011100000100;
      patterns[47143] = 29'b1_011100000100_111_1_011100000100;
      patterns[47144] = 29'b1_011100000101_000_1_011100000101;
      patterns[47145] = 29'b1_011100000101_001_1_000101011100;
      patterns[47146] = 29'b1_011100000101_010_0_111000001011;
      patterns[47147] = 29'b1_011100000101_011_1_110000010110;
      patterns[47148] = 29'b1_011100000101_100_1_101110000010;
      patterns[47149] = 29'b1_011100000101_101_0_110111000001;
      patterns[47150] = 29'b1_011100000101_110_1_011100000101;
      patterns[47151] = 29'b1_011100000101_111_1_011100000101;
      patterns[47152] = 29'b1_011100000110_000_1_011100000110;
      patterns[47153] = 29'b1_011100000110_001_1_000110011100;
      patterns[47154] = 29'b1_011100000110_010_0_111000001101;
      patterns[47155] = 29'b1_011100000110_011_1_110000011010;
      patterns[47156] = 29'b1_011100000110_100_0_101110000011;
      patterns[47157] = 29'b1_011100000110_101_1_010111000001;
      patterns[47158] = 29'b1_011100000110_110_1_011100000110;
      patterns[47159] = 29'b1_011100000110_111_1_011100000110;
      patterns[47160] = 29'b1_011100000111_000_1_011100000111;
      patterns[47161] = 29'b1_011100000111_001_1_000111011100;
      patterns[47162] = 29'b1_011100000111_010_0_111000001111;
      patterns[47163] = 29'b1_011100000111_011_1_110000011110;
      patterns[47164] = 29'b1_011100000111_100_1_101110000011;
      patterns[47165] = 29'b1_011100000111_101_1_110111000001;
      patterns[47166] = 29'b1_011100000111_110_1_011100000111;
      patterns[47167] = 29'b1_011100000111_111_1_011100000111;
      patterns[47168] = 29'b1_011100001000_000_1_011100001000;
      patterns[47169] = 29'b1_011100001000_001_1_001000011100;
      patterns[47170] = 29'b1_011100001000_010_0_111000010001;
      patterns[47171] = 29'b1_011100001000_011_1_110000100010;
      patterns[47172] = 29'b1_011100001000_100_0_101110000100;
      patterns[47173] = 29'b1_011100001000_101_0_010111000010;
      patterns[47174] = 29'b1_011100001000_110_1_011100001000;
      patterns[47175] = 29'b1_011100001000_111_1_011100001000;
      patterns[47176] = 29'b1_011100001001_000_1_011100001001;
      patterns[47177] = 29'b1_011100001001_001_1_001001011100;
      patterns[47178] = 29'b1_011100001001_010_0_111000010011;
      patterns[47179] = 29'b1_011100001001_011_1_110000100110;
      patterns[47180] = 29'b1_011100001001_100_1_101110000100;
      patterns[47181] = 29'b1_011100001001_101_0_110111000010;
      patterns[47182] = 29'b1_011100001001_110_1_011100001001;
      patterns[47183] = 29'b1_011100001001_111_1_011100001001;
      patterns[47184] = 29'b1_011100001010_000_1_011100001010;
      patterns[47185] = 29'b1_011100001010_001_1_001010011100;
      patterns[47186] = 29'b1_011100001010_010_0_111000010101;
      patterns[47187] = 29'b1_011100001010_011_1_110000101010;
      patterns[47188] = 29'b1_011100001010_100_0_101110000101;
      patterns[47189] = 29'b1_011100001010_101_1_010111000010;
      patterns[47190] = 29'b1_011100001010_110_1_011100001010;
      patterns[47191] = 29'b1_011100001010_111_1_011100001010;
      patterns[47192] = 29'b1_011100001011_000_1_011100001011;
      patterns[47193] = 29'b1_011100001011_001_1_001011011100;
      patterns[47194] = 29'b1_011100001011_010_0_111000010111;
      patterns[47195] = 29'b1_011100001011_011_1_110000101110;
      patterns[47196] = 29'b1_011100001011_100_1_101110000101;
      patterns[47197] = 29'b1_011100001011_101_1_110111000010;
      patterns[47198] = 29'b1_011100001011_110_1_011100001011;
      patterns[47199] = 29'b1_011100001011_111_1_011100001011;
      patterns[47200] = 29'b1_011100001100_000_1_011100001100;
      patterns[47201] = 29'b1_011100001100_001_1_001100011100;
      patterns[47202] = 29'b1_011100001100_010_0_111000011001;
      patterns[47203] = 29'b1_011100001100_011_1_110000110010;
      patterns[47204] = 29'b1_011100001100_100_0_101110000110;
      patterns[47205] = 29'b1_011100001100_101_0_010111000011;
      patterns[47206] = 29'b1_011100001100_110_1_011100001100;
      patterns[47207] = 29'b1_011100001100_111_1_011100001100;
      patterns[47208] = 29'b1_011100001101_000_1_011100001101;
      patterns[47209] = 29'b1_011100001101_001_1_001101011100;
      patterns[47210] = 29'b1_011100001101_010_0_111000011011;
      patterns[47211] = 29'b1_011100001101_011_1_110000110110;
      patterns[47212] = 29'b1_011100001101_100_1_101110000110;
      patterns[47213] = 29'b1_011100001101_101_0_110111000011;
      patterns[47214] = 29'b1_011100001101_110_1_011100001101;
      patterns[47215] = 29'b1_011100001101_111_1_011100001101;
      patterns[47216] = 29'b1_011100001110_000_1_011100001110;
      patterns[47217] = 29'b1_011100001110_001_1_001110011100;
      patterns[47218] = 29'b1_011100001110_010_0_111000011101;
      patterns[47219] = 29'b1_011100001110_011_1_110000111010;
      patterns[47220] = 29'b1_011100001110_100_0_101110000111;
      patterns[47221] = 29'b1_011100001110_101_1_010111000011;
      patterns[47222] = 29'b1_011100001110_110_1_011100001110;
      patterns[47223] = 29'b1_011100001110_111_1_011100001110;
      patterns[47224] = 29'b1_011100001111_000_1_011100001111;
      patterns[47225] = 29'b1_011100001111_001_1_001111011100;
      patterns[47226] = 29'b1_011100001111_010_0_111000011111;
      patterns[47227] = 29'b1_011100001111_011_1_110000111110;
      patterns[47228] = 29'b1_011100001111_100_1_101110000111;
      patterns[47229] = 29'b1_011100001111_101_1_110111000011;
      patterns[47230] = 29'b1_011100001111_110_1_011100001111;
      patterns[47231] = 29'b1_011100001111_111_1_011100001111;
      patterns[47232] = 29'b1_011100010000_000_1_011100010000;
      patterns[47233] = 29'b1_011100010000_001_1_010000011100;
      patterns[47234] = 29'b1_011100010000_010_0_111000100001;
      patterns[47235] = 29'b1_011100010000_011_1_110001000010;
      patterns[47236] = 29'b1_011100010000_100_0_101110001000;
      patterns[47237] = 29'b1_011100010000_101_0_010111000100;
      patterns[47238] = 29'b1_011100010000_110_1_011100010000;
      patterns[47239] = 29'b1_011100010000_111_1_011100010000;
      patterns[47240] = 29'b1_011100010001_000_1_011100010001;
      patterns[47241] = 29'b1_011100010001_001_1_010001011100;
      patterns[47242] = 29'b1_011100010001_010_0_111000100011;
      patterns[47243] = 29'b1_011100010001_011_1_110001000110;
      patterns[47244] = 29'b1_011100010001_100_1_101110001000;
      patterns[47245] = 29'b1_011100010001_101_0_110111000100;
      patterns[47246] = 29'b1_011100010001_110_1_011100010001;
      patterns[47247] = 29'b1_011100010001_111_1_011100010001;
      patterns[47248] = 29'b1_011100010010_000_1_011100010010;
      patterns[47249] = 29'b1_011100010010_001_1_010010011100;
      patterns[47250] = 29'b1_011100010010_010_0_111000100101;
      patterns[47251] = 29'b1_011100010010_011_1_110001001010;
      patterns[47252] = 29'b1_011100010010_100_0_101110001001;
      patterns[47253] = 29'b1_011100010010_101_1_010111000100;
      patterns[47254] = 29'b1_011100010010_110_1_011100010010;
      patterns[47255] = 29'b1_011100010010_111_1_011100010010;
      patterns[47256] = 29'b1_011100010011_000_1_011100010011;
      patterns[47257] = 29'b1_011100010011_001_1_010011011100;
      patterns[47258] = 29'b1_011100010011_010_0_111000100111;
      patterns[47259] = 29'b1_011100010011_011_1_110001001110;
      patterns[47260] = 29'b1_011100010011_100_1_101110001001;
      patterns[47261] = 29'b1_011100010011_101_1_110111000100;
      patterns[47262] = 29'b1_011100010011_110_1_011100010011;
      patterns[47263] = 29'b1_011100010011_111_1_011100010011;
      patterns[47264] = 29'b1_011100010100_000_1_011100010100;
      patterns[47265] = 29'b1_011100010100_001_1_010100011100;
      patterns[47266] = 29'b1_011100010100_010_0_111000101001;
      patterns[47267] = 29'b1_011100010100_011_1_110001010010;
      patterns[47268] = 29'b1_011100010100_100_0_101110001010;
      patterns[47269] = 29'b1_011100010100_101_0_010111000101;
      patterns[47270] = 29'b1_011100010100_110_1_011100010100;
      patterns[47271] = 29'b1_011100010100_111_1_011100010100;
      patterns[47272] = 29'b1_011100010101_000_1_011100010101;
      patterns[47273] = 29'b1_011100010101_001_1_010101011100;
      patterns[47274] = 29'b1_011100010101_010_0_111000101011;
      patterns[47275] = 29'b1_011100010101_011_1_110001010110;
      patterns[47276] = 29'b1_011100010101_100_1_101110001010;
      patterns[47277] = 29'b1_011100010101_101_0_110111000101;
      patterns[47278] = 29'b1_011100010101_110_1_011100010101;
      patterns[47279] = 29'b1_011100010101_111_1_011100010101;
      patterns[47280] = 29'b1_011100010110_000_1_011100010110;
      patterns[47281] = 29'b1_011100010110_001_1_010110011100;
      patterns[47282] = 29'b1_011100010110_010_0_111000101101;
      patterns[47283] = 29'b1_011100010110_011_1_110001011010;
      patterns[47284] = 29'b1_011100010110_100_0_101110001011;
      patterns[47285] = 29'b1_011100010110_101_1_010111000101;
      patterns[47286] = 29'b1_011100010110_110_1_011100010110;
      patterns[47287] = 29'b1_011100010110_111_1_011100010110;
      patterns[47288] = 29'b1_011100010111_000_1_011100010111;
      patterns[47289] = 29'b1_011100010111_001_1_010111011100;
      patterns[47290] = 29'b1_011100010111_010_0_111000101111;
      patterns[47291] = 29'b1_011100010111_011_1_110001011110;
      patterns[47292] = 29'b1_011100010111_100_1_101110001011;
      patterns[47293] = 29'b1_011100010111_101_1_110111000101;
      patterns[47294] = 29'b1_011100010111_110_1_011100010111;
      patterns[47295] = 29'b1_011100010111_111_1_011100010111;
      patterns[47296] = 29'b1_011100011000_000_1_011100011000;
      patterns[47297] = 29'b1_011100011000_001_1_011000011100;
      patterns[47298] = 29'b1_011100011000_010_0_111000110001;
      patterns[47299] = 29'b1_011100011000_011_1_110001100010;
      patterns[47300] = 29'b1_011100011000_100_0_101110001100;
      patterns[47301] = 29'b1_011100011000_101_0_010111000110;
      patterns[47302] = 29'b1_011100011000_110_1_011100011000;
      patterns[47303] = 29'b1_011100011000_111_1_011100011000;
      patterns[47304] = 29'b1_011100011001_000_1_011100011001;
      patterns[47305] = 29'b1_011100011001_001_1_011001011100;
      patterns[47306] = 29'b1_011100011001_010_0_111000110011;
      patterns[47307] = 29'b1_011100011001_011_1_110001100110;
      patterns[47308] = 29'b1_011100011001_100_1_101110001100;
      patterns[47309] = 29'b1_011100011001_101_0_110111000110;
      patterns[47310] = 29'b1_011100011001_110_1_011100011001;
      patterns[47311] = 29'b1_011100011001_111_1_011100011001;
      patterns[47312] = 29'b1_011100011010_000_1_011100011010;
      patterns[47313] = 29'b1_011100011010_001_1_011010011100;
      patterns[47314] = 29'b1_011100011010_010_0_111000110101;
      patterns[47315] = 29'b1_011100011010_011_1_110001101010;
      patterns[47316] = 29'b1_011100011010_100_0_101110001101;
      patterns[47317] = 29'b1_011100011010_101_1_010111000110;
      patterns[47318] = 29'b1_011100011010_110_1_011100011010;
      patterns[47319] = 29'b1_011100011010_111_1_011100011010;
      patterns[47320] = 29'b1_011100011011_000_1_011100011011;
      patterns[47321] = 29'b1_011100011011_001_1_011011011100;
      patterns[47322] = 29'b1_011100011011_010_0_111000110111;
      patterns[47323] = 29'b1_011100011011_011_1_110001101110;
      patterns[47324] = 29'b1_011100011011_100_1_101110001101;
      patterns[47325] = 29'b1_011100011011_101_1_110111000110;
      patterns[47326] = 29'b1_011100011011_110_1_011100011011;
      patterns[47327] = 29'b1_011100011011_111_1_011100011011;
      patterns[47328] = 29'b1_011100011100_000_1_011100011100;
      patterns[47329] = 29'b1_011100011100_001_1_011100011100;
      patterns[47330] = 29'b1_011100011100_010_0_111000111001;
      patterns[47331] = 29'b1_011100011100_011_1_110001110010;
      patterns[47332] = 29'b1_011100011100_100_0_101110001110;
      patterns[47333] = 29'b1_011100011100_101_0_010111000111;
      patterns[47334] = 29'b1_011100011100_110_1_011100011100;
      patterns[47335] = 29'b1_011100011100_111_1_011100011100;
      patterns[47336] = 29'b1_011100011101_000_1_011100011101;
      patterns[47337] = 29'b1_011100011101_001_1_011101011100;
      patterns[47338] = 29'b1_011100011101_010_0_111000111011;
      patterns[47339] = 29'b1_011100011101_011_1_110001110110;
      patterns[47340] = 29'b1_011100011101_100_1_101110001110;
      patterns[47341] = 29'b1_011100011101_101_0_110111000111;
      patterns[47342] = 29'b1_011100011101_110_1_011100011101;
      patterns[47343] = 29'b1_011100011101_111_1_011100011101;
      patterns[47344] = 29'b1_011100011110_000_1_011100011110;
      patterns[47345] = 29'b1_011100011110_001_1_011110011100;
      patterns[47346] = 29'b1_011100011110_010_0_111000111101;
      patterns[47347] = 29'b1_011100011110_011_1_110001111010;
      patterns[47348] = 29'b1_011100011110_100_0_101110001111;
      patterns[47349] = 29'b1_011100011110_101_1_010111000111;
      patterns[47350] = 29'b1_011100011110_110_1_011100011110;
      patterns[47351] = 29'b1_011100011110_111_1_011100011110;
      patterns[47352] = 29'b1_011100011111_000_1_011100011111;
      patterns[47353] = 29'b1_011100011111_001_1_011111011100;
      patterns[47354] = 29'b1_011100011111_010_0_111000111111;
      patterns[47355] = 29'b1_011100011111_011_1_110001111110;
      patterns[47356] = 29'b1_011100011111_100_1_101110001111;
      patterns[47357] = 29'b1_011100011111_101_1_110111000111;
      patterns[47358] = 29'b1_011100011111_110_1_011100011111;
      patterns[47359] = 29'b1_011100011111_111_1_011100011111;
      patterns[47360] = 29'b1_011100100000_000_1_011100100000;
      patterns[47361] = 29'b1_011100100000_001_1_100000011100;
      patterns[47362] = 29'b1_011100100000_010_0_111001000001;
      patterns[47363] = 29'b1_011100100000_011_1_110010000010;
      patterns[47364] = 29'b1_011100100000_100_0_101110010000;
      patterns[47365] = 29'b1_011100100000_101_0_010111001000;
      patterns[47366] = 29'b1_011100100000_110_1_011100100000;
      patterns[47367] = 29'b1_011100100000_111_1_011100100000;
      patterns[47368] = 29'b1_011100100001_000_1_011100100001;
      patterns[47369] = 29'b1_011100100001_001_1_100001011100;
      patterns[47370] = 29'b1_011100100001_010_0_111001000011;
      patterns[47371] = 29'b1_011100100001_011_1_110010000110;
      patterns[47372] = 29'b1_011100100001_100_1_101110010000;
      patterns[47373] = 29'b1_011100100001_101_0_110111001000;
      patterns[47374] = 29'b1_011100100001_110_1_011100100001;
      patterns[47375] = 29'b1_011100100001_111_1_011100100001;
      patterns[47376] = 29'b1_011100100010_000_1_011100100010;
      patterns[47377] = 29'b1_011100100010_001_1_100010011100;
      patterns[47378] = 29'b1_011100100010_010_0_111001000101;
      patterns[47379] = 29'b1_011100100010_011_1_110010001010;
      patterns[47380] = 29'b1_011100100010_100_0_101110010001;
      patterns[47381] = 29'b1_011100100010_101_1_010111001000;
      patterns[47382] = 29'b1_011100100010_110_1_011100100010;
      patterns[47383] = 29'b1_011100100010_111_1_011100100010;
      patterns[47384] = 29'b1_011100100011_000_1_011100100011;
      patterns[47385] = 29'b1_011100100011_001_1_100011011100;
      patterns[47386] = 29'b1_011100100011_010_0_111001000111;
      patterns[47387] = 29'b1_011100100011_011_1_110010001110;
      patterns[47388] = 29'b1_011100100011_100_1_101110010001;
      patterns[47389] = 29'b1_011100100011_101_1_110111001000;
      patterns[47390] = 29'b1_011100100011_110_1_011100100011;
      patterns[47391] = 29'b1_011100100011_111_1_011100100011;
      patterns[47392] = 29'b1_011100100100_000_1_011100100100;
      patterns[47393] = 29'b1_011100100100_001_1_100100011100;
      patterns[47394] = 29'b1_011100100100_010_0_111001001001;
      patterns[47395] = 29'b1_011100100100_011_1_110010010010;
      patterns[47396] = 29'b1_011100100100_100_0_101110010010;
      patterns[47397] = 29'b1_011100100100_101_0_010111001001;
      patterns[47398] = 29'b1_011100100100_110_1_011100100100;
      patterns[47399] = 29'b1_011100100100_111_1_011100100100;
      patterns[47400] = 29'b1_011100100101_000_1_011100100101;
      patterns[47401] = 29'b1_011100100101_001_1_100101011100;
      patterns[47402] = 29'b1_011100100101_010_0_111001001011;
      patterns[47403] = 29'b1_011100100101_011_1_110010010110;
      patterns[47404] = 29'b1_011100100101_100_1_101110010010;
      patterns[47405] = 29'b1_011100100101_101_0_110111001001;
      patterns[47406] = 29'b1_011100100101_110_1_011100100101;
      patterns[47407] = 29'b1_011100100101_111_1_011100100101;
      patterns[47408] = 29'b1_011100100110_000_1_011100100110;
      patterns[47409] = 29'b1_011100100110_001_1_100110011100;
      patterns[47410] = 29'b1_011100100110_010_0_111001001101;
      patterns[47411] = 29'b1_011100100110_011_1_110010011010;
      patterns[47412] = 29'b1_011100100110_100_0_101110010011;
      patterns[47413] = 29'b1_011100100110_101_1_010111001001;
      patterns[47414] = 29'b1_011100100110_110_1_011100100110;
      patterns[47415] = 29'b1_011100100110_111_1_011100100110;
      patterns[47416] = 29'b1_011100100111_000_1_011100100111;
      patterns[47417] = 29'b1_011100100111_001_1_100111011100;
      patterns[47418] = 29'b1_011100100111_010_0_111001001111;
      patterns[47419] = 29'b1_011100100111_011_1_110010011110;
      patterns[47420] = 29'b1_011100100111_100_1_101110010011;
      patterns[47421] = 29'b1_011100100111_101_1_110111001001;
      patterns[47422] = 29'b1_011100100111_110_1_011100100111;
      patterns[47423] = 29'b1_011100100111_111_1_011100100111;
      patterns[47424] = 29'b1_011100101000_000_1_011100101000;
      patterns[47425] = 29'b1_011100101000_001_1_101000011100;
      patterns[47426] = 29'b1_011100101000_010_0_111001010001;
      patterns[47427] = 29'b1_011100101000_011_1_110010100010;
      patterns[47428] = 29'b1_011100101000_100_0_101110010100;
      patterns[47429] = 29'b1_011100101000_101_0_010111001010;
      patterns[47430] = 29'b1_011100101000_110_1_011100101000;
      patterns[47431] = 29'b1_011100101000_111_1_011100101000;
      patterns[47432] = 29'b1_011100101001_000_1_011100101001;
      patterns[47433] = 29'b1_011100101001_001_1_101001011100;
      patterns[47434] = 29'b1_011100101001_010_0_111001010011;
      patterns[47435] = 29'b1_011100101001_011_1_110010100110;
      patterns[47436] = 29'b1_011100101001_100_1_101110010100;
      patterns[47437] = 29'b1_011100101001_101_0_110111001010;
      patterns[47438] = 29'b1_011100101001_110_1_011100101001;
      patterns[47439] = 29'b1_011100101001_111_1_011100101001;
      patterns[47440] = 29'b1_011100101010_000_1_011100101010;
      patterns[47441] = 29'b1_011100101010_001_1_101010011100;
      patterns[47442] = 29'b1_011100101010_010_0_111001010101;
      patterns[47443] = 29'b1_011100101010_011_1_110010101010;
      patterns[47444] = 29'b1_011100101010_100_0_101110010101;
      patterns[47445] = 29'b1_011100101010_101_1_010111001010;
      patterns[47446] = 29'b1_011100101010_110_1_011100101010;
      patterns[47447] = 29'b1_011100101010_111_1_011100101010;
      patterns[47448] = 29'b1_011100101011_000_1_011100101011;
      patterns[47449] = 29'b1_011100101011_001_1_101011011100;
      patterns[47450] = 29'b1_011100101011_010_0_111001010111;
      patterns[47451] = 29'b1_011100101011_011_1_110010101110;
      patterns[47452] = 29'b1_011100101011_100_1_101110010101;
      patterns[47453] = 29'b1_011100101011_101_1_110111001010;
      patterns[47454] = 29'b1_011100101011_110_1_011100101011;
      patterns[47455] = 29'b1_011100101011_111_1_011100101011;
      patterns[47456] = 29'b1_011100101100_000_1_011100101100;
      patterns[47457] = 29'b1_011100101100_001_1_101100011100;
      patterns[47458] = 29'b1_011100101100_010_0_111001011001;
      patterns[47459] = 29'b1_011100101100_011_1_110010110010;
      patterns[47460] = 29'b1_011100101100_100_0_101110010110;
      patterns[47461] = 29'b1_011100101100_101_0_010111001011;
      patterns[47462] = 29'b1_011100101100_110_1_011100101100;
      patterns[47463] = 29'b1_011100101100_111_1_011100101100;
      patterns[47464] = 29'b1_011100101101_000_1_011100101101;
      patterns[47465] = 29'b1_011100101101_001_1_101101011100;
      patterns[47466] = 29'b1_011100101101_010_0_111001011011;
      patterns[47467] = 29'b1_011100101101_011_1_110010110110;
      patterns[47468] = 29'b1_011100101101_100_1_101110010110;
      patterns[47469] = 29'b1_011100101101_101_0_110111001011;
      patterns[47470] = 29'b1_011100101101_110_1_011100101101;
      patterns[47471] = 29'b1_011100101101_111_1_011100101101;
      patterns[47472] = 29'b1_011100101110_000_1_011100101110;
      patterns[47473] = 29'b1_011100101110_001_1_101110011100;
      patterns[47474] = 29'b1_011100101110_010_0_111001011101;
      patterns[47475] = 29'b1_011100101110_011_1_110010111010;
      patterns[47476] = 29'b1_011100101110_100_0_101110010111;
      patterns[47477] = 29'b1_011100101110_101_1_010111001011;
      patterns[47478] = 29'b1_011100101110_110_1_011100101110;
      patterns[47479] = 29'b1_011100101110_111_1_011100101110;
      patterns[47480] = 29'b1_011100101111_000_1_011100101111;
      patterns[47481] = 29'b1_011100101111_001_1_101111011100;
      patterns[47482] = 29'b1_011100101111_010_0_111001011111;
      patterns[47483] = 29'b1_011100101111_011_1_110010111110;
      patterns[47484] = 29'b1_011100101111_100_1_101110010111;
      patterns[47485] = 29'b1_011100101111_101_1_110111001011;
      patterns[47486] = 29'b1_011100101111_110_1_011100101111;
      patterns[47487] = 29'b1_011100101111_111_1_011100101111;
      patterns[47488] = 29'b1_011100110000_000_1_011100110000;
      patterns[47489] = 29'b1_011100110000_001_1_110000011100;
      patterns[47490] = 29'b1_011100110000_010_0_111001100001;
      patterns[47491] = 29'b1_011100110000_011_1_110011000010;
      patterns[47492] = 29'b1_011100110000_100_0_101110011000;
      patterns[47493] = 29'b1_011100110000_101_0_010111001100;
      patterns[47494] = 29'b1_011100110000_110_1_011100110000;
      patterns[47495] = 29'b1_011100110000_111_1_011100110000;
      patterns[47496] = 29'b1_011100110001_000_1_011100110001;
      patterns[47497] = 29'b1_011100110001_001_1_110001011100;
      patterns[47498] = 29'b1_011100110001_010_0_111001100011;
      patterns[47499] = 29'b1_011100110001_011_1_110011000110;
      patterns[47500] = 29'b1_011100110001_100_1_101110011000;
      patterns[47501] = 29'b1_011100110001_101_0_110111001100;
      patterns[47502] = 29'b1_011100110001_110_1_011100110001;
      patterns[47503] = 29'b1_011100110001_111_1_011100110001;
      patterns[47504] = 29'b1_011100110010_000_1_011100110010;
      patterns[47505] = 29'b1_011100110010_001_1_110010011100;
      patterns[47506] = 29'b1_011100110010_010_0_111001100101;
      patterns[47507] = 29'b1_011100110010_011_1_110011001010;
      patterns[47508] = 29'b1_011100110010_100_0_101110011001;
      patterns[47509] = 29'b1_011100110010_101_1_010111001100;
      patterns[47510] = 29'b1_011100110010_110_1_011100110010;
      patterns[47511] = 29'b1_011100110010_111_1_011100110010;
      patterns[47512] = 29'b1_011100110011_000_1_011100110011;
      patterns[47513] = 29'b1_011100110011_001_1_110011011100;
      patterns[47514] = 29'b1_011100110011_010_0_111001100111;
      patterns[47515] = 29'b1_011100110011_011_1_110011001110;
      patterns[47516] = 29'b1_011100110011_100_1_101110011001;
      patterns[47517] = 29'b1_011100110011_101_1_110111001100;
      patterns[47518] = 29'b1_011100110011_110_1_011100110011;
      patterns[47519] = 29'b1_011100110011_111_1_011100110011;
      patterns[47520] = 29'b1_011100110100_000_1_011100110100;
      patterns[47521] = 29'b1_011100110100_001_1_110100011100;
      patterns[47522] = 29'b1_011100110100_010_0_111001101001;
      patterns[47523] = 29'b1_011100110100_011_1_110011010010;
      patterns[47524] = 29'b1_011100110100_100_0_101110011010;
      patterns[47525] = 29'b1_011100110100_101_0_010111001101;
      patterns[47526] = 29'b1_011100110100_110_1_011100110100;
      patterns[47527] = 29'b1_011100110100_111_1_011100110100;
      patterns[47528] = 29'b1_011100110101_000_1_011100110101;
      patterns[47529] = 29'b1_011100110101_001_1_110101011100;
      patterns[47530] = 29'b1_011100110101_010_0_111001101011;
      patterns[47531] = 29'b1_011100110101_011_1_110011010110;
      patterns[47532] = 29'b1_011100110101_100_1_101110011010;
      patterns[47533] = 29'b1_011100110101_101_0_110111001101;
      patterns[47534] = 29'b1_011100110101_110_1_011100110101;
      patterns[47535] = 29'b1_011100110101_111_1_011100110101;
      patterns[47536] = 29'b1_011100110110_000_1_011100110110;
      patterns[47537] = 29'b1_011100110110_001_1_110110011100;
      patterns[47538] = 29'b1_011100110110_010_0_111001101101;
      patterns[47539] = 29'b1_011100110110_011_1_110011011010;
      patterns[47540] = 29'b1_011100110110_100_0_101110011011;
      patterns[47541] = 29'b1_011100110110_101_1_010111001101;
      patterns[47542] = 29'b1_011100110110_110_1_011100110110;
      patterns[47543] = 29'b1_011100110110_111_1_011100110110;
      patterns[47544] = 29'b1_011100110111_000_1_011100110111;
      patterns[47545] = 29'b1_011100110111_001_1_110111011100;
      patterns[47546] = 29'b1_011100110111_010_0_111001101111;
      patterns[47547] = 29'b1_011100110111_011_1_110011011110;
      patterns[47548] = 29'b1_011100110111_100_1_101110011011;
      patterns[47549] = 29'b1_011100110111_101_1_110111001101;
      patterns[47550] = 29'b1_011100110111_110_1_011100110111;
      patterns[47551] = 29'b1_011100110111_111_1_011100110111;
      patterns[47552] = 29'b1_011100111000_000_1_011100111000;
      patterns[47553] = 29'b1_011100111000_001_1_111000011100;
      patterns[47554] = 29'b1_011100111000_010_0_111001110001;
      patterns[47555] = 29'b1_011100111000_011_1_110011100010;
      patterns[47556] = 29'b1_011100111000_100_0_101110011100;
      patterns[47557] = 29'b1_011100111000_101_0_010111001110;
      patterns[47558] = 29'b1_011100111000_110_1_011100111000;
      patterns[47559] = 29'b1_011100111000_111_1_011100111000;
      patterns[47560] = 29'b1_011100111001_000_1_011100111001;
      patterns[47561] = 29'b1_011100111001_001_1_111001011100;
      patterns[47562] = 29'b1_011100111001_010_0_111001110011;
      patterns[47563] = 29'b1_011100111001_011_1_110011100110;
      patterns[47564] = 29'b1_011100111001_100_1_101110011100;
      patterns[47565] = 29'b1_011100111001_101_0_110111001110;
      patterns[47566] = 29'b1_011100111001_110_1_011100111001;
      patterns[47567] = 29'b1_011100111001_111_1_011100111001;
      patterns[47568] = 29'b1_011100111010_000_1_011100111010;
      patterns[47569] = 29'b1_011100111010_001_1_111010011100;
      patterns[47570] = 29'b1_011100111010_010_0_111001110101;
      patterns[47571] = 29'b1_011100111010_011_1_110011101010;
      patterns[47572] = 29'b1_011100111010_100_0_101110011101;
      patterns[47573] = 29'b1_011100111010_101_1_010111001110;
      patterns[47574] = 29'b1_011100111010_110_1_011100111010;
      patterns[47575] = 29'b1_011100111010_111_1_011100111010;
      patterns[47576] = 29'b1_011100111011_000_1_011100111011;
      patterns[47577] = 29'b1_011100111011_001_1_111011011100;
      patterns[47578] = 29'b1_011100111011_010_0_111001110111;
      patterns[47579] = 29'b1_011100111011_011_1_110011101110;
      patterns[47580] = 29'b1_011100111011_100_1_101110011101;
      patterns[47581] = 29'b1_011100111011_101_1_110111001110;
      patterns[47582] = 29'b1_011100111011_110_1_011100111011;
      patterns[47583] = 29'b1_011100111011_111_1_011100111011;
      patterns[47584] = 29'b1_011100111100_000_1_011100111100;
      patterns[47585] = 29'b1_011100111100_001_1_111100011100;
      patterns[47586] = 29'b1_011100111100_010_0_111001111001;
      patterns[47587] = 29'b1_011100111100_011_1_110011110010;
      patterns[47588] = 29'b1_011100111100_100_0_101110011110;
      patterns[47589] = 29'b1_011100111100_101_0_010111001111;
      patterns[47590] = 29'b1_011100111100_110_1_011100111100;
      patterns[47591] = 29'b1_011100111100_111_1_011100111100;
      patterns[47592] = 29'b1_011100111101_000_1_011100111101;
      patterns[47593] = 29'b1_011100111101_001_1_111101011100;
      patterns[47594] = 29'b1_011100111101_010_0_111001111011;
      patterns[47595] = 29'b1_011100111101_011_1_110011110110;
      patterns[47596] = 29'b1_011100111101_100_1_101110011110;
      patterns[47597] = 29'b1_011100111101_101_0_110111001111;
      patterns[47598] = 29'b1_011100111101_110_1_011100111101;
      patterns[47599] = 29'b1_011100111101_111_1_011100111101;
      patterns[47600] = 29'b1_011100111110_000_1_011100111110;
      patterns[47601] = 29'b1_011100111110_001_1_111110011100;
      patterns[47602] = 29'b1_011100111110_010_0_111001111101;
      patterns[47603] = 29'b1_011100111110_011_1_110011111010;
      patterns[47604] = 29'b1_011100111110_100_0_101110011111;
      patterns[47605] = 29'b1_011100111110_101_1_010111001111;
      patterns[47606] = 29'b1_011100111110_110_1_011100111110;
      patterns[47607] = 29'b1_011100111110_111_1_011100111110;
      patterns[47608] = 29'b1_011100111111_000_1_011100111111;
      patterns[47609] = 29'b1_011100111111_001_1_111111011100;
      patterns[47610] = 29'b1_011100111111_010_0_111001111111;
      patterns[47611] = 29'b1_011100111111_011_1_110011111110;
      patterns[47612] = 29'b1_011100111111_100_1_101110011111;
      patterns[47613] = 29'b1_011100111111_101_1_110111001111;
      patterns[47614] = 29'b1_011100111111_110_1_011100111111;
      patterns[47615] = 29'b1_011100111111_111_1_011100111111;
      patterns[47616] = 29'b1_011101000000_000_1_011101000000;
      patterns[47617] = 29'b1_011101000000_001_1_000000011101;
      patterns[47618] = 29'b1_011101000000_010_0_111010000001;
      patterns[47619] = 29'b1_011101000000_011_1_110100000010;
      patterns[47620] = 29'b1_011101000000_100_0_101110100000;
      patterns[47621] = 29'b1_011101000000_101_0_010111010000;
      patterns[47622] = 29'b1_011101000000_110_1_011101000000;
      patterns[47623] = 29'b1_011101000000_111_1_011101000000;
      patterns[47624] = 29'b1_011101000001_000_1_011101000001;
      patterns[47625] = 29'b1_011101000001_001_1_000001011101;
      patterns[47626] = 29'b1_011101000001_010_0_111010000011;
      patterns[47627] = 29'b1_011101000001_011_1_110100000110;
      patterns[47628] = 29'b1_011101000001_100_1_101110100000;
      patterns[47629] = 29'b1_011101000001_101_0_110111010000;
      patterns[47630] = 29'b1_011101000001_110_1_011101000001;
      patterns[47631] = 29'b1_011101000001_111_1_011101000001;
      patterns[47632] = 29'b1_011101000010_000_1_011101000010;
      patterns[47633] = 29'b1_011101000010_001_1_000010011101;
      patterns[47634] = 29'b1_011101000010_010_0_111010000101;
      patterns[47635] = 29'b1_011101000010_011_1_110100001010;
      patterns[47636] = 29'b1_011101000010_100_0_101110100001;
      patterns[47637] = 29'b1_011101000010_101_1_010111010000;
      patterns[47638] = 29'b1_011101000010_110_1_011101000010;
      patterns[47639] = 29'b1_011101000010_111_1_011101000010;
      patterns[47640] = 29'b1_011101000011_000_1_011101000011;
      patterns[47641] = 29'b1_011101000011_001_1_000011011101;
      patterns[47642] = 29'b1_011101000011_010_0_111010000111;
      patterns[47643] = 29'b1_011101000011_011_1_110100001110;
      patterns[47644] = 29'b1_011101000011_100_1_101110100001;
      patterns[47645] = 29'b1_011101000011_101_1_110111010000;
      patterns[47646] = 29'b1_011101000011_110_1_011101000011;
      patterns[47647] = 29'b1_011101000011_111_1_011101000011;
      patterns[47648] = 29'b1_011101000100_000_1_011101000100;
      patterns[47649] = 29'b1_011101000100_001_1_000100011101;
      patterns[47650] = 29'b1_011101000100_010_0_111010001001;
      patterns[47651] = 29'b1_011101000100_011_1_110100010010;
      patterns[47652] = 29'b1_011101000100_100_0_101110100010;
      patterns[47653] = 29'b1_011101000100_101_0_010111010001;
      patterns[47654] = 29'b1_011101000100_110_1_011101000100;
      patterns[47655] = 29'b1_011101000100_111_1_011101000100;
      patterns[47656] = 29'b1_011101000101_000_1_011101000101;
      patterns[47657] = 29'b1_011101000101_001_1_000101011101;
      patterns[47658] = 29'b1_011101000101_010_0_111010001011;
      patterns[47659] = 29'b1_011101000101_011_1_110100010110;
      patterns[47660] = 29'b1_011101000101_100_1_101110100010;
      patterns[47661] = 29'b1_011101000101_101_0_110111010001;
      patterns[47662] = 29'b1_011101000101_110_1_011101000101;
      patterns[47663] = 29'b1_011101000101_111_1_011101000101;
      patterns[47664] = 29'b1_011101000110_000_1_011101000110;
      patterns[47665] = 29'b1_011101000110_001_1_000110011101;
      patterns[47666] = 29'b1_011101000110_010_0_111010001101;
      patterns[47667] = 29'b1_011101000110_011_1_110100011010;
      patterns[47668] = 29'b1_011101000110_100_0_101110100011;
      patterns[47669] = 29'b1_011101000110_101_1_010111010001;
      patterns[47670] = 29'b1_011101000110_110_1_011101000110;
      patterns[47671] = 29'b1_011101000110_111_1_011101000110;
      patterns[47672] = 29'b1_011101000111_000_1_011101000111;
      patterns[47673] = 29'b1_011101000111_001_1_000111011101;
      patterns[47674] = 29'b1_011101000111_010_0_111010001111;
      patterns[47675] = 29'b1_011101000111_011_1_110100011110;
      patterns[47676] = 29'b1_011101000111_100_1_101110100011;
      patterns[47677] = 29'b1_011101000111_101_1_110111010001;
      patterns[47678] = 29'b1_011101000111_110_1_011101000111;
      patterns[47679] = 29'b1_011101000111_111_1_011101000111;
      patterns[47680] = 29'b1_011101001000_000_1_011101001000;
      patterns[47681] = 29'b1_011101001000_001_1_001000011101;
      patterns[47682] = 29'b1_011101001000_010_0_111010010001;
      patterns[47683] = 29'b1_011101001000_011_1_110100100010;
      patterns[47684] = 29'b1_011101001000_100_0_101110100100;
      patterns[47685] = 29'b1_011101001000_101_0_010111010010;
      patterns[47686] = 29'b1_011101001000_110_1_011101001000;
      patterns[47687] = 29'b1_011101001000_111_1_011101001000;
      patterns[47688] = 29'b1_011101001001_000_1_011101001001;
      patterns[47689] = 29'b1_011101001001_001_1_001001011101;
      patterns[47690] = 29'b1_011101001001_010_0_111010010011;
      patterns[47691] = 29'b1_011101001001_011_1_110100100110;
      patterns[47692] = 29'b1_011101001001_100_1_101110100100;
      patterns[47693] = 29'b1_011101001001_101_0_110111010010;
      patterns[47694] = 29'b1_011101001001_110_1_011101001001;
      patterns[47695] = 29'b1_011101001001_111_1_011101001001;
      patterns[47696] = 29'b1_011101001010_000_1_011101001010;
      patterns[47697] = 29'b1_011101001010_001_1_001010011101;
      patterns[47698] = 29'b1_011101001010_010_0_111010010101;
      patterns[47699] = 29'b1_011101001010_011_1_110100101010;
      patterns[47700] = 29'b1_011101001010_100_0_101110100101;
      patterns[47701] = 29'b1_011101001010_101_1_010111010010;
      patterns[47702] = 29'b1_011101001010_110_1_011101001010;
      patterns[47703] = 29'b1_011101001010_111_1_011101001010;
      patterns[47704] = 29'b1_011101001011_000_1_011101001011;
      patterns[47705] = 29'b1_011101001011_001_1_001011011101;
      patterns[47706] = 29'b1_011101001011_010_0_111010010111;
      patterns[47707] = 29'b1_011101001011_011_1_110100101110;
      patterns[47708] = 29'b1_011101001011_100_1_101110100101;
      patterns[47709] = 29'b1_011101001011_101_1_110111010010;
      patterns[47710] = 29'b1_011101001011_110_1_011101001011;
      patterns[47711] = 29'b1_011101001011_111_1_011101001011;
      patterns[47712] = 29'b1_011101001100_000_1_011101001100;
      patterns[47713] = 29'b1_011101001100_001_1_001100011101;
      patterns[47714] = 29'b1_011101001100_010_0_111010011001;
      patterns[47715] = 29'b1_011101001100_011_1_110100110010;
      patterns[47716] = 29'b1_011101001100_100_0_101110100110;
      patterns[47717] = 29'b1_011101001100_101_0_010111010011;
      patterns[47718] = 29'b1_011101001100_110_1_011101001100;
      patterns[47719] = 29'b1_011101001100_111_1_011101001100;
      patterns[47720] = 29'b1_011101001101_000_1_011101001101;
      patterns[47721] = 29'b1_011101001101_001_1_001101011101;
      patterns[47722] = 29'b1_011101001101_010_0_111010011011;
      patterns[47723] = 29'b1_011101001101_011_1_110100110110;
      patterns[47724] = 29'b1_011101001101_100_1_101110100110;
      patterns[47725] = 29'b1_011101001101_101_0_110111010011;
      patterns[47726] = 29'b1_011101001101_110_1_011101001101;
      patterns[47727] = 29'b1_011101001101_111_1_011101001101;
      patterns[47728] = 29'b1_011101001110_000_1_011101001110;
      patterns[47729] = 29'b1_011101001110_001_1_001110011101;
      patterns[47730] = 29'b1_011101001110_010_0_111010011101;
      patterns[47731] = 29'b1_011101001110_011_1_110100111010;
      patterns[47732] = 29'b1_011101001110_100_0_101110100111;
      patterns[47733] = 29'b1_011101001110_101_1_010111010011;
      patterns[47734] = 29'b1_011101001110_110_1_011101001110;
      patterns[47735] = 29'b1_011101001110_111_1_011101001110;
      patterns[47736] = 29'b1_011101001111_000_1_011101001111;
      patterns[47737] = 29'b1_011101001111_001_1_001111011101;
      patterns[47738] = 29'b1_011101001111_010_0_111010011111;
      patterns[47739] = 29'b1_011101001111_011_1_110100111110;
      patterns[47740] = 29'b1_011101001111_100_1_101110100111;
      patterns[47741] = 29'b1_011101001111_101_1_110111010011;
      patterns[47742] = 29'b1_011101001111_110_1_011101001111;
      patterns[47743] = 29'b1_011101001111_111_1_011101001111;
      patterns[47744] = 29'b1_011101010000_000_1_011101010000;
      patterns[47745] = 29'b1_011101010000_001_1_010000011101;
      patterns[47746] = 29'b1_011101010000_010_0_111010100001;
      patterns[47747] = 29'b1_011101010000_011_1_110101000010;
      patterns[47748] = 29'b1_011101010000_100_0_101110101000;
      patterns[47749] = 29'b1_011101010000_101_0_010111010100;
      patterns[47750] = 29'b1_011101010000_110_1_011101010000;
      patterns[47751] = 29'b1_011101010000_111_1_011101010000;
      patterns[47752] = 29'b1_011101010001_000_1_011101010001;
      patterns[47753] = 29'b1_011101010001_001_1_010001011101;
      patterns[47754] = 29'b1_011101010001_010_0_111010100011;
      patterns[47755] = 29'b1_011101010001_011_1_110101000110;
      patterns[47756] = 29'b1_011101010001_100_1_101110101000;
      patterns[47757] = 29'b1_011101010001_101_0_110111010100;
      patterns[47758] = 29'b1_011101010001_110_1_011101010001;
      patterns[47759] = 29'b1_011101010001_111_1_011101010001;
      patterns[47760] = 29'b1_011101010010_000_1_011101010010;
      patterns[47761] = 29'b1_011101010010_001_1_010010011101;
      patterns[47762] = 29'b1_011101010010_010_0_111010100101;
      patterns[47763] = 29'b1_011101010010_011_1_110101001010;
      patterns[47764] = 29'b1_011101010010_100_0_101110101001;
      patterns[47765] = 29'b1_011101010010_101_1_010111010100;
      patterns[47766] = 29'b1_011101010010_110_1_011101010010;
      patterns[47767] = 29'b1_011101010010_111_1_011101010010;
      patterns[47768] = 29'b1_011101010011_000_1_011101010011;
      patterns[47769] = 29'b1_011101010011_001_1_010011011101;
      patterns[47770] = 29'b1_011101010011_010_0_111010100111;
      patterns[47771] = 29'b1_011101010011_011_1_110101001110;
      patterns[47772] = 29'b1_011101010011_100_1_101110101001;
      patterns[47773] = 29'b1_011101010011_101_1_110111010100;
      patterns[47774] = 29'b1_011101010011_110_1_011101010011;
      patterns[47775] = 29'b1_011101010011_111_1_011101010011;
      patterns[47776] = 29'b1_011101010100_000_1_011101010100;
      patterns[47777] = 29'b1_011101010100_001_1_010100011101;
      patterns[47778] = 29'b1_011101010100_010_0_111010101001;
      patterns[47779] = 29'b1_011101010100_011_1_110101010010;
      patterns[47780] = 29'b1_011101010100_100_0_101110101010;
      patterns[47781] = 29'b1_011101010100_101_0_010111010101;
      patterns[47782] = 29'b1_011101010100_110_1_011101010100;
      patterns[47783] = 29'b1_011101010100_111_1_011101010100;
      patterns[47784] = 29'b1_011101010101_000_1_011101010101;
      patterns[47785] = 29'b1_011101010101_001_1_010101011101;
      patterns[47786] = 29'b1_011101010101_010_0_111010101011;
      patterns[47787] = 29'b1_011101010101_011_1_110101010110;
      patterns[47788] = 29'b1_011101010101_100_1_101110101010;
      patterns[47789] = 29'b1_011101010101_101_0_110111010101;
      patterns[47790] = 29'b1_011101010101_110_1_011101010101;
      patterns[47791] = 29'b1_011101010101_111_1_011101010101;
      patterns[47792] = 29'b1_011101010110_000_1_011101010110;
      patterns[47793] = 29'b1_011101010110_001_1_010110011101;
      patterns[47794] = 29'b1_011101010110_010_0_111010101101;
      patterns[47795] = 29'b1_011101010110_011_1_110101011010;
      patterns[47796] = 29'b1_011101010110_100_0_101110101011;
      patterns[47797] = 29'b1_011101010110_101_1_010111010101;
      patterns[47798] = 29'b1_011101010110_110_1_011101010110;
      patterns[47799] = 29'b1_011101010110_111_1_011101010110;
      patterns[47800] = 29'b1_011101010111_000_1_011101010111;
      patterns[47801] = 29'b1_011101010111_001_1_010111011101;
      patterns[47802] = 29'b1_011101010111_010_0_111010101111;
      patterns[47803] = 29'b1_011101010111_011_1_110101011110;
      patterns[47804] = 29'b1_011101010111_100_1_101110101011;
      patterns[47805] = 29'b1_011101010111_101_1_110111010101;
      patterns[47806] = 29'b1_011101010111_110_1_011101010111;
      patterns[47807] = 29'b1_011101010111_111_1_011101010111;
      patterns[47808] = 29'b1_011101011000_000_1_011101011000;
      patterns[47809] = 29'b1_011101011000_001_1_011000011101;
      patterns[47810] = 29'b1_011101011000_010_0_111010110001;
      patterns[47811] = 29'b1_011101011000_011_1_110101100010;
      patterns[47812] = 29'b1_011101011000_100_0_101110101100;
      patterns[47813] = 29'b1_011101011000_101_0_010111010110;
      patterns[47814] = 29'b1_011101011000_110_1_011101011000;
      patterns[47815] = 29'b1_011101011000_111_1_011101011000;
      patterns[47816] = 29'b1_011101011001_000_1_011101011001;
      patterns[47817] = 29'b1_011101011001_001_1_011001011101;
      patterns[47818] = 29'b1_011101011001_010_0_111010110011;
      patterns[47819] = 29'b1_011101011001_011_1_110101100110;
      patterns[47820] = 29'b1_011101011001_100_1_101110101100;
      patterns[47821] = 29'b1_011101011001_101_0_110111010110;
      patterns[47822] = 29'b1_011101011001_110_1_011101011001;
      patterns[47823] = 29'b1_011101011001_111_1_011101011001;
      patterns[47824] = 29'b1_011101011010_000_1_011101011010;
      patterns[47825] = 29'b1_011101011010_001_1_011010011101;
      patterns[47826] = 29'b1_011101011010_010_0_111010110101;
      patterns[47827] = 29'b1_011101011010_011_1_110101101010;
      patterns[47828] = 29'b1_011101011010_100_0_101110101101;
      patterns[47829] = 29'b1_011101011010_101_1_010111010110;
      patterns[47830] = 29'b1_011101011010_110_1_011101011010;
      patterns[47831] = 29'b1_011101011010_111_1_011101011010;
      patterns[47832] = 29'b1_011101011011_000_1_011101011011;
      patterns[47833] = 29'b1_011101011011_001_1_011011011101;
      patterns[47834] = 29'b1_011101011011_010_0_111010110111;
      patterns[47835] = 29'b1_011101011011_011_1_110101101110;
      patterns[47836] = 29'b1_011101011011_100_1_101110101101;
      patterns[47837] = 29'b1_011101011011_101_1_110111010110;
      patterns[47838] = 29'b1_011101011011_110_1_011101011011;
      patterns[47839] = 29'b1_011101011011_111_1_011101011011;
      patterns[47840] = 29'b1_011101011100_000_1_011101011100;
      patterns[47841] = 29'b1_011101011100_001_1_011100011101;
      patterns[47842] = 29'b1_011101011100_010_0_111010111001;
      patterns[47843] = 29'b1_011101011100_011_1_110101110010;
      patterns[47844] = 29'b1_011101011100_100_0_101110101110;
      patterns[47845] = 29'b1_011101011100_101_0_010111010111;
      patterns[47846] = 29'b1_011101011100_110_1_011101011100;
      patterns[47847] = 29'b1_011101011100_111_1_011101011100;
      patterns[47848] = 29'b1_011101011101_000_1_011101011101;
      patterns[47849] = 29'b1_011101011101_001_1_011101011101;
      patterns[47850] = 29'b1_011101011101_010_0_111010111011;
      patterns[47851] = 29'b1_011101011101_011_1_110101110110;
      patterns[47852] = 29'b1_011101011101_100_1_101110101110;
      patterns[47853] = 29'b1_011101011101_101_0_110111010111;
      patterns[47854] = 29'b1_011101011101_110_1_011101011101;
      patterns[47855] = 29'b1_011101011101_111_1_011101011101;
      patterns[47856] = 29'b1_011101011110_000_1_011101011110;
      patterns[47857] = 29'b1_011101011110_001_1_011110011101;
      patterns[47858] = 29'b1_011101011110_010_0_111010111101;
      patterns[47859] = 29'b1_011101011110_011_1_110101111010;
      patterns[47860] = 29'b1_011101011110_100_0_101110101111;
      patterns[47861] = 29'b1_011101011110_101_1_010111010111;
      patterns[47862] = 29'b1_011101011110_110_1_011101011110;
      patterns[47863] = 29'b1_011101011110_111_1_011101011110;
      patterns[47864] = 29'b1_011101011111_000_1_011101011111;
      patterns[47865] = 29'b1_011101011111_001_1_011111011101;
      patterns[47866] = 29'b1_011101011111_010_0_111010111111;
      patterns[47867] = 29'b1_011101011111_011_1_110101111110;
      patterns[47868] = 29'b1_011101011111_100_1_101110101111;
      patterns[47869] = 29'b1_011101011111_101_1_110111010111;
      patterns[47870] = 29'b1_011101011111_110_1_011101011111;
      patterns[47871] = 29'b1_011101011111_111_1_011101011111;
      patterns[47872] = 29'b1_011101100000_000_1_011101100000;
      patterns[47873] = 29'b1_011101100000_001_1_100000011101;
      patterns[47874] = 29'b1_011101100000_010_0_111011000001;
      patterns[47875] = 29'b1_011101100000_011_1_110110000010;
      patterns[47876] = 29'b1_011101100000_100_0_101110110000;
      patterns[47877] = 29'b1_011101100000_101_0_010111011000;
      patterns[47878] = 29'b1_011101100000_110_1_011101100000;
      patterns[47879] = 29'b1_011101100000_111_1_011101100000;
      patterns[47880] = 29'b1_011101100001_000_1_011101100001;
      patterns[47881] = 29'b1_011101100001_001_1_100001011101;
      patterns[47882] = 29'b1_011101100001_010_0_111011000011;
      patterns[47883] = 29'b1_011101100001_011_1_110110000110;
      patterns[47884] = 29'b1_011101100001_100_1_101110110000;
      patterns[47885] = 29'b1_011101100001_101_0_110111011000;
      patterns[47886] = 29'b1_011101100001_110_1_011101100001;
      patterns[47887] = 29'b1_011101100001_111_1_011101100001;
      patterns[47888] = 29'b1_011101100010_000_1_011101100010;
      patterns[47889] = 29'b1_011101100010_001_1_100010011101;
      patterns[47890] = 29'b1_011101100010_010_0_111011000101;
      patterns[47891] = 29'b1_011101100010_011_1_110110001010;
      patterns[47892] = 29'b1_011101100010_100_0_101110110001;
      patterns[47893] = 29'b1_011101100010_101_1_010111011000;
      patterns[47894] = 29'b1_011101100010_110_1_011101100010;
      patterns[47895] = 29'b1_011101100010_111_1_011101100010;
      patterns[47896] = 29'b1_011101100011_000_1_011101100011;
      patterns[47897] = 29'b1_011101100011_001_1_100011011101;
      patterns[47898] = 29'b1_011101100011_010_0_111011000111;
      patterns[47899] = 29'b1_011101100011_011_1_110110001110;
      patterns[47900] = 29'b1_011101100011_100_1_101110110001;
      patterns[47901] = 29'b1_011101100011_101_1_110111011000;
      patterns[47902] = 29'b1_011101100011_110_1_011101100011;
      patterns[47903] = 29'b1_011101100011_111_1_011101100011;
      patterns[47904] = 29'b1_011101100100_000_1_011101100100;
      patterns[47905] = 29'b1_011101100100_001_1_100100011101;
      patterns[47906] = 29'b1_011101100100_010_0_111011001001;
      patterns[47907] = 29'b1_011101100100_011_1_110110010010;
      patterns[47908] = 29'b1_011101100100_100_0_101110110010;
      patterns[47909] = 29'b1_011101100100_101_0_010111011001;
      patterns[47910] = 29'b1_011101100100_110_1_011101100100;
      patterns[47911] = 29'b1_011101100100_111_1_011101100100;
      patterns[47912] = 29'b1_011101100101_000_1_011101100101;
      patterns[47913] = 29'b1_011101100101_001_1_100101011101;
      patterns[47914] = 29'b1_011101100101_010_0_111011001011;
      patterns[47915] = 29'b1_011101100101_011_1_110110010110;
      patterns[47916] = 29'b1_011101100101_100_1_101110110010;
      patterns[47917] = 29'b1_011101100101_101_0_110111011001;
      patterns[47918] = 29'b1_011101100101_110_1_011101100101;
      patterns[47919] = 29'b1_011101100101_111_1_011101100101;
      patterns[47920] = 29'b1_011101100110_000_1_011101100110;
      patterns[47921] = 29'b1_011101100110_001_1_100110011101;
      patterns[47922] = 29'b1_011101100110_010_0_111011001101;
      patterns[47923] = 29'b1_011101100110_011_1_110110011010;
      patterns[47924] = 29'b1_011101100110_100_0_101110110011;
      patterns[47925] = 29'b1_011101100110_101_1_010111011001;
      patterns[47926] = 29'b1_011101100110_110_1_011101100110;
      patterns[47927] = 29'b1_011101100110_111_1_011101100110;
      patterns[47928] = 29'b1_011101100111_000_1_011101100111;
      patterns[47929] = 29'b1_011101100111_001_1_100111011101;
      patterns[47930] = 29'b1_011101100111_010_0_111011001111;
      patterns[47931] = 29'b1_011101100111_011_1_110110011110;
      patterns[47932] = 29'b1_011101100111_100_1_101110110011;
      patterns[47933] = 29'b1_011101100111_101_1_110111011001;
      patterns[47934] = 29'b1_011101100111_110_1_011101100111;
      patterns[47935] = 29'b1_011101100111_111_1_011101100111;
      patterns[47936] = 29'b1_011101101000_000_1_011101101000;
      patterns[47937] = 29'b1_011101101000_001_1_101000011101;
      patterns[47938] = 29'b1_011101101000_010_0_111011010001;
      patterns[47939] = 29'b1_011101101000_011_1_110110100010;
      patterns[47940] = 29'b1_011101101000_100_0_101110110100;
      patterns[47941] = 29'b1_011101101000_101_0_010111011010;
      patterns[47942] = 29'b1_011101101000_110_1_011101101000;
      patterns[47943] = 29'b1_011101101000_111_1_011101101000;
      patterns[47944] = 29'b1_011101101001_000_1_011101101001;
      patterns[47945] = 29'b1_011101101001_001_1_101001011101;
      patterns[47946] = 29'b1_011101101001_010_0_111011010011;
      patterns[47947] = 29'b1_011101101001_011_1_110110100110;
      patterns[47948] = 29'b1_011101101001_100_1_101110110100;
      patterns[47949] = 29'b1_011101101001_101_0_110111011010;
      patterns[47950] = 29'b1_011101101001_110_1_011101101001;
      patterns[47951] = 29'b1_011101101001_111_1_011101101001;
      patterns[47952] = 29'b1_011101101010_000_1_011101101010;
      patterns[47953] = 29'b1_011101101010_001_1_101010011101;
      patterns[47954] = 29'b1_011101101010_010_0_111011010101;
      patterns[47955] = 29'b1_011101101010_011_1_110110101010;
      patterns[47956] = 29'b1_011101101010_100_0_101110110101;
      patterns[47957] = 29'b1_011101101010_101_1_010111011010;
      patterns[47958] = 29'b1_011101101010_110_1_011101101010;
      patterns[47959] = 29'b1_011101101010_111_1_011101101010;
      patterns[47960] = 29'b1_011101101011_000_1_011101101011;
      patterns[47961] = 29'b1_011101101011_001_1_101011011101;
      patterns[47962] = 29'b1_011101101011_010_0_111011010111;
      patterns[47963] = 29'b1_011101101011_011_1_110110101110;
      patterns[47964] = 29'b1_011101101011_100_1_101110110101;
      patterns[47965] = 29'b1_011101101011_101_1_110111011010;
      patterns[47966] = 29'b1_011101101011_110_1_011101101011;
      patterns[47967] = 29'b1_011101101011_111_1_011101101011;
      patterns[47968] = 29'b1_011101101100_000_1_011101101100;
      patterns[47969] = 29'b1_011101101100_001_1_101100011101;
      patterns[47970] = 29'b1_011101101100_010_0_111011011001;
      patterns[47971] = 29'b1_011101101100_011_1_110110110010;
      patterns[47972] = 29'b1_011101101100_100_0_101110110110;
      patterns[47973] = 29'b1_011101101100_101_0_010111011011;
      patterns[47974] = 29'b1_011101101100_110_1_011101101100;
      patterns[47975] = 29'b1_011101101100_111_1_011101101100;
      patterns[47976] = 29'b1_011101101101_000_1_011101101101;
      patterns[47977] = 29'b1_011101101101_001_1_101101011101;
      patterns[47978] = 29'b1_011101101101_010_0_111011011011;
      patterns[47979] = 29'b1_011101101101_011_1_110110110110;
      patterns[47980] = 29'b1_011101101101_100_1_101110110110;
      patterns[47981] = 29'b1_011101101101_101_0_110111011011;
      patterns[47982] = 29'b1_011101101101_110_1_011101101101;
      patterns[47983] = 29'b1_011101101101_111_1_011101101101;
      patterns[47984] = 29'b1_011101101110_000_1_011101101110;
      patterns[47985] = 29'b1_011101101110_001_1_101110011101;
      patterns[47986] = 29'b1_011101101110_010_0_111011011101;
      patterns[47987] = 29'b1_011101101110_011_1_110110111010;
      patterns[47988] = 29'b1_011101101110_100_0_101110110111;
      patterns[47989] = 29'b1_011101101110_101_1_010111011011;
      patterns[47990] = 29'b1_011101101110_110_1_011101101110;
      patterns[47991] = 29'b1_011101101110_111_1_011101101110;
      patterns[47992] = 29'b1_011101101111_000_1_011101101111;
      patterns[47993] = 29'b1_011101101111_001_1_101111011101;
      patterns[47994] = 29'b1_011101101111_010_0_111011011111;
      patterns[47995] = 29'b1_011101101111_011_1_110110111110;
      patterns[47996] = 29'b1_011101101111_100_1_101110110111;
      patterns[47997] = 29'b1_011101101111_101_1_110111011011;
      patterns[47998] = 29'b1_011101101111_110_1_011101101111;
      patterns[47999] = 29'b1_011101101111_111_1_011101101111;
      patterns[48000] = 29'b1_011101110000_000_1_011101110000;
      patterns[48001] = 29'b1_011101110000_001_1_110000011101;
      patterns[48002] = 29'b1_011101110000_010_0_111011100001;
      patterns[48003] = 29'b1_011101110000_011_1_110111000010;
      patterns[48004] = 29'b1_011101110000_100_0_101110111000;
      patterns[48005] = 29'b1_011101110000_101_0_010111011100;
      patterns[48006] = 29'b1_011101110000_110_1_011101110000;
      patterns[48007] = 29'b1_011101110000_111_1_011101110000;
      patterns[48008] = 29'b1_011101110001_000_1_011101110001;
      patterns[48009] = 29'b1_011101110001_001_1_110001011101;
      patterns[48010] = 29'b1_011101110001_010_0_111011100011;
      patterns[48011] = 29'b1_011101110001_011_1_110111000110;
      patterns[48012] = 29'b1_011101110001_100_1_101110111000;
      patterns[48013] = 29'b1_011101110001_101_0_110111011100;
      patterns[48014] = 29'b1_011101110001_110_1_011101110001;
      patterns[48015] = 29'b1_011101110001_111_1_011101110001;
      patterns[48016] = 29'b1_011101110010_000_1_011101110010;
      patterns[48017] = 29'b1_011101110010_001_1_110010011101;
      patterns[48018] = 29'b1_011101110010_010_0_111011100101;
      patterns[48019] = 29'b1_011101110010_011_1_110111001010;
      patterns[48020] = 29'b1_011101110010_100_0_101110111001;
      patterns[48021] = 29'b1_011101110010_101_1_010111011100;
      patterns[48022] = 29'b1_011101110010_110_1_011101110010;
      patterns[48023] = 29'b1_011101110010_111_1_011101110010;
      patterns[48024] = 29'b1_011101110011_000_1_011101110011;
      patterns[48025] = 29'b1_011101110011_001_1_110011011101;
      patterns[48026] = 29'b1_011101110011_010_0_111011100111;
      patterns[48027] = 29'b1_011101110011_011_1_110111001110;
      patterns[48028] = 29'b1_011101110011_100_1_101110111001;
      patterns[48029] = 29'b1_011101110011_101_1_110111011100;
      patterns[48030] = 29'b1_011101110011_110_1_011101110011;
      patterns[48031] = 29'b1_011101110011_111_1_011101110011;
      patterns[48032] = 29'b1_011101110100_000_1_011101110100;
      patterns[48033] = 29'b1_011101110100_001_1_110100011101;
      patterns[48034] = 29'b1_011101110100_010_0_111011101001;
      patterns[48035] = 29'b1_011101110100_011_1_110111010010;
      patterns[48036] = 29'b1_011101110100_100_0_101110111010;
      patterns[48037] = 29'b1_011101110100_101_0_010111011101;
      patterns[48038] = 29'b1_011101110100_110_1_011101110100;
      patterns[48039] = 29'b1_011101110100_111_1_011101110100;
      patterns[48040] = 29'b1_011101110101_000_1_011101110101;
      patterns[48041] = 29'b1_011101110101_001_1_110101011101;
      patterns[48042] = 29'b1_011101110101_010_0_111011101011;
      patterns[48043] = 29'b1_011101110101_011_1_110111010110;
      patterns[48044] = 29'b1_011101110101_100_1_101110111010;
      patterns[48045] = 29'b1_011101110101_101_0_110111011101;
      patterns[48046] = 29'b1_011101110101_110_1_011101110101;
      patterns[48047] = 29'b1_011101110101_111_1_011101110101;
      patterns[48048] = 29'b1_011101110110_000_1_011101110110;
      patterns[48049] = 29'b1_011101110110_001_1_110110011101;
      patterns[48050] = 29'b1_011101110110_010_0_111011101101;
      patterns[48051] = 29'b1_011101110110_011_1_110111011010;
      patterns[48052] = 29'b1_011101110110_100_0_101110111011;
      patterns[48053] = 29'b1_011101110110_101_1_010111011101;
      patterns[48054] = 29'b1_011101110110_110_1_011101110110;
      patterns[48055] = 29'b1_011101110110_111_1_011101110110;
      patterns[48056] = 29'b1_011101110111_000_1_011101110111;
      patterns[48057] = 29'b1_011101110111_001_1_110111011101;
      patterns[48058] = 29'b1_011101110111_010_0_111011101111;
      patterns[48059] = 29'b1_011101110111_011_1_110111011110;
      patterns[48060] = 29'b1_011101110111_100_1_101110111011;
      patterns[48061] = 29'b1_011101110111_101_1_110111011101;
      patterns[48062] = 29'b1_011101110111_110_1_011101110111;
      patterns[48063] = 29'b1_011101110111_111_1_011101110111;
      patterns[48064] = 29'b1_011101111000_000_1_011101111000;
      patterns[48065] = 29'b1_011101111000_001_1_111000011101;
      patterns[48066] = 29'b1_011101111000_010_0_111011110001;
      patterns[48067] = 29'b1_011101111000_011_1_110111100010;
      patterns[48068] = 29'b1_011101111000_100_0_101110111100;
      patterns[48069] = 29'b1_011101111000_101_0_010111011110;
      patterns[48070] = 29'b1_011101111000_110_1_011101111000;
      patterns[48071] = 29'b1_011101111000_111_1_011101111000;
      patterns[48072] = 29'b1_011101111001_000_1_011101111001;
      patterns[48073] = 29'b1_011101111001_001_1_111001011101;
      patterns[48074] = 29'b1_011101111001_010_0_111011110011;
      patterns[48075] = 29'b1_011101111001_011_1_110111100110;
      patterns[48076] = 29'b1_011101111001_100_1_101110111100;
      patterns[48077] = 29'b1_011101111001_101_0_110111011110;
      patterns[48078] = 29'b1_011101111001_110_1_011101111001;
      patterns[48079] = 29'b1_011101111001_111_1_011101111001;
      patterns[48080] = 29'b1_011101111010_000_1_011101111010;
      patterns[48081] = 29'b1_011101111010_001_1_111010011101;
      patterns[48082] = 29'b1_011101111010_010_0_111011110101;
      patterns[48083] = 29'b1_011101111010_011_1_110111101010;
      patterns[48084] = 29'b1_011101111010_100_0_101110111101;
      patterns[48085] = 29'b1_011101111010_101_1_010111011110;
      patterns[48086] = 29'b1_011101111010_110_1_011101111010;
      patterns[48087] = 29'b1_011101111010_111_1_011101111010;
      patterns[48088] = 29'b1_011101111011_000_1_011101111011;
      patterns[48089] = 29'b1_011101111011_001_1_111011011101;
      patterns[48090] = 29'b1_011101111011_010_0_111011110111;
      patterns[48091] = 29'b1_011101111011_011_1_110111101110;
      patterns[48092] = 29'b1_011101111011_100_1_101110111101;
      patterns[48093] = 29'b1_011101111011_101_1_110111011110;
      patterns[48094] = 29'b1_011101111011_110_1_011101111011;
      patterns[48095] = 29'b1_011101111011_111_1_011101111011;
      patterns[48096] = 29'b1_011101111100_000_1_011101111100;
      patterns[48097] = 29'b1_011101111100_001_1_111100011101;
      patterns[48098] = 29'b1_011101111100_010_0_111011111001;
      patterns[48099] = 29'b1_011101111100_011_1_110111110010;
      patterns[48100] = 29'b1_011101111100_100_0_101110111110;
      patterns[48101] = 29'b1_011101111100_101_0_010111011111;
      patterns[48102] = 29'b1_011101111100_110_1_011101111100;
      patterns[48103] = 29'b1_011101111100_111_1_011101111100;
      patterns[48104] = 29'b1_011101111101_000_1_011101111101;
      patterns[48105] = 29'b1_011101111101_001_1_111101011101;
      patterns[48106] = 29'b1_011101111101_010_0_111011111011;
      patterns[48107] = 29'b1_011101111101_011_1_110111110110;
      patterns[48108] = 29'b1_011101111101_100_1_101110111110;
      patterns[48109] = 29'b1_011101111101_101_0_110111011111;
      patterns[48110] = 29'b1_011101111101_110_1_011101111101;
      patterns[48111] = 29'b1_011101111101_111_1_011101111101;
      patterns[48112] = 29'b1_011101111110_000_1_011101111110;
      patterns[48113] = 29'b1_011101111110_001_1_111110011101;
      patterns[48114] = 29'b1_011101111110_010_0_111011111101;
      patterns[48115] = 29'b1_011101111110_011_1_110111111010;
      patterns[48116] = 29'b1_011101111110_100_0_101110111111;
      patterns[48117] = 29'b1_011101111110_101_1_010111011111;
      patterns[48118] = 29'b1_011101111110_110_1_011101111110;
      patterns[48119] = 29'b1_011101111110_111_1_011101111110;
      patterns[48120] = 29'b1_011101111111_000_1_011101111111;
      patterns[48121] = 29'b1_011101111111_001_1_111111011101;
      patterns[48122] = 29'b1_011101111111_010_0_111011111111;
      patterns[48123] = 29'b1_011101111111_011_1_110111111110;
      patterns[48124] = 29'b1_011101111111_100_1_101110111111;
      patterns[48125] = 29'b1_011101111111_101_1_110111011111;
      patterns[48126] = 29'b1_011101111111_110_1_011101111111;
      patterns[48127] = 29'b1_011101111111_111_1_011101111111;
      patterns[48128] = 29'b1_011110000000_000_1_011110000000;
      patterns[48129] = 29'b1_011110000000_001_1_000000011110;
      patterns[48130] = 29'b1_011110000000_010_0_111100000001;
      patterns[48131] = 29'b1_011110000000_011_1_111000000010;
      patterns[48132] = 29'b1_011110000000_100_0_101111000000;
      patterns[48133] = 29'b1_011110000000_101_0_010111100000;
      patterns[48134] = 29'b1_011110000000_110_1_011110000000;
      patterns[48135] = 29'b1_011110000000_111_1_011110000000;
      patterns[48136] = 29'b1_011110000001_000_1_011110000001;
      patterns[48137] = 29'b1_011110000001_001_1_000001011110;
      patterns[48138] = 29'b1_011110000001_010_0_111100000011;
      patterns[48139] = 29'b1_011110000001_011_1_111000000110;
      patterns[48140] = 29'b1_011110000001_100_1_101111000000;
      patterns[48141] = 29'b1_011110000001_101_0_110111100000;
      patterns[48142] = 29'b1_011110000001_110_1_011110000001;
      patterns[48143] = 29'b1_011110000001_111_1_011110000001;
      patterns[48144] = 29'b1_011110000010_000_1_011110000010;
      patterns[48145] = 29'b1_011110000010_001_1_000010011110;
      patterns[48146] = 29'b1_011110000010_010_0_111100000101;
      patterns[48147] = 29'b1_011110000010_011_1_111000001010;
      patterns[48148] = 29'b1_011110000010_100_0_101111000001;
      patterns[48149] = 29'b1_011110000010_101_1_010111100000;
      patterns[48150] = 29'b1_011110000010_110_1_011110000010;
      patterns[48151] = 29'b1_011110000010_111_1_011110000010;
      patterns[48152] = 29'b1_011110000011_000_1_011110000011;
      patterns[48153] = 29'b1_011110000011_001_1_000011011110;
      patterns[48154] = 29'b1_011110000011_010_0_111100000111;
      patterns[48155] = 29'b1_011110000011_011_1_111000001110;
      patterns[48156] = 29'b1_011110000011_100_1_101111000001;
      patterns[48157] = 29'b1_011110000011_101_1_110111100000;
      patterns[48158] = 29'b1_011110000011_110_1_011110000011;
      patterns[48159] = 29'b1_011110000011_111_1_011110000011;
      patterns[48160] = 29'b1_011110000100_000_1_011110000100;
      patterns[48161] = 29'b1_011110000100_001_1_000100011110;
      patterns[48162] = 29'b1_011110000100_010_0_111100001001;
      patterns[48163] = 29'b1_011110000100_011_1_111000010010;
      patterns[48164] = 29'b1_011110000100_100_0_101111000010;
      patterns[48165] = 29'b1_011110000100_101_0_010111100001;
      patterns[48166] = 29'b1_011110000100_110_1_011110000100;
      patterns[48167] = 29'b1_011110000100_111_1_011110000100;
      patterns[48168] = 29'b1_011110000101_000_1_011110000101;
      patterns[48169] = 29'b1_011110000101_001_1_000101011110;
      patterns[48170] = 29'b1_011110000101_010_0_111100001011;
      patterns[48171] = 29'b1_011110000101_011_1_111000010110;
      patterns[48172] = 29'b1_011110000101_100_1_101111000010;
      patterns[48173] = 29'b1_011110000101_101_0_110111100001;
      patterns[48174] = 29'b1_011110000101_110_1_011110000101;
      patterns[48175] = 29'b1_011110000101_111_1_011110000101;
      patterns[48176] = 29'b1_011110000110_000_1_011110000110;
      patterns[48177] = 29'b1_011110000110_001_1_000110011110;
      patterns[48178] = 29'b1_011110000110_010_0_111100001101;
      patterns[48179] = 29'b1_011110000110_011_1_111000011010;
      patterns[48180] = 29'b1_011110000110_100_0_101111000011;
      patterns[48181] = 29'b1_011110000110_101_1_010111100001;
      patterns[48182] = 29'b1_011110000110_110_1_011110000110;
      patterns[48183] = 29'b1_011110000110_111_1_011110000110;
      patterns[48184] = 29'b1_011110000111_000_1_011110000111;
      patterns[48185] = 29'b1_011110000111_001_1_000111011110;
      patterns[48186] = 29'b1_011110000111_010_0_111100001111;
      patterns[48187] = 29'b1_011110000111_011_1_111000011110;
      patterns[48188] = 29'b1_011110000111_100_1_101111000011;
      patterns[48189] = 29'b1_011110000111_101_1_110111100001;
      patterns[48190] = 29'b1_011110000111_110_1_011110000111;
      patterns[48191] = 29'b1_011110000111_111_1_011110000111;
      patterns[48192] = 29'b1_011110001000_000_1_011110001000;
      patterns[48193] = 29'b1_011110001000_001_1_001000011110;
      patterns[48194] = 29'b1_011110001000_010_0_111100010001;
      patterns[48195] = 29'b1_011110001000_011_1_111000100010;
      patterns[48196] = 29'b1_011110001000_100_0_101111000100;
      patterns[48197] = 29'b1_011110001000_101_0_010111100010;
      patterns[48198] = 29'b1_011110001000_110_1_011110001000;
      patterns[48199] = 29'b1_011110001000_111_1_011110001000;
      patterns[48200] = 29'b1_011110001001_000_1_011110001001;
      patterns[48201] = 29'b1_011110001001_001_1_001001011110;
      patterns[48202] = 29'b1_011110001001_010_0_111100010011;
      patterns[48203] = 29'b1_011110001001_011_1_111000100110;
      patterns[48204] = 29'b1_011110001001_100_1_101111000100;
      patterns[48205] = 29'b1_011110001001_101_0_110111100010;
      patterns[48206] = 29'b1_011110001001_110_1_011110001001;
      patterns[48207] = 29'b1_011110001001_111_1_011110001001;
      patterns[48208] = 29'b1_011110001010_000_1_011110001010;
      patterns[48209] = 29'b1_011110001010_001_1_001010011110;
      patterns[48210] = 29'b1_011110001010_010_0_111100010101;
      patterns[48211] = 29'b1_011110001010_011_1_111000101010;
      patterns[48212] = 29'b1_011110001010_100_0_101111000101;
      patterns[48213] = 29'b1_011110001010_101_1_010111100010;
      patterns[48214] = 29'b1_011110001010_110_1_011110001010;
      patterns[48215] = 29'b1_011110001010_111_1_011110001010;
      patterns[48216] = 29'b1_011110001011_000_1_011110001011;
      patterns[48217] = 29'b1_011110001011_001_1_001011011110;
      patterns[48218] = 29'b1_011110001011_010_0_111100010111;
      patterns[48219] = 29'b1_011110001011_011_1_111000101110;
      patterns[48220] = 29'b1_011110001011_100_1_101111000101;
      patterns[48221] = 29'b1_011110001011_101_1_110111100010;
      patterns[48222] = 29'b1_011110001011_110_1_011110001011;
      patterns[48223] = 29'b1_011110001011_111_1_011110001011;
      patterns[48224] = 29'b1_011110001100_000_1_011110001100;
      patterns[48225] = 29'b1_011110001100_001_1_001100011110;
      patterns[48226] = 29'b1_011110001100_010_0_111100011001;
      patterns[48227] = 29'b1_011110001100_011_1_111000110010;
      patterns[48228] = 29'b1_011110001100_100_0_101111000110;
      patterns[48229] = 29'b1_011110001100_101_0_010111100011;
      patterns[48230] = 29'b1_011110001100_110_1_011110001100;
      patterns[48231] = 29'b1_011110001100_111_1_011110001100;
      patterns[48232] = 29'b1_011110001101_000_1_011110001101;
      patterns[48233] = 29'b1_011110001101_001_1_001101011110;
      patterns[48234] = 29'b1_011110001101_010_0_111100011011;
      patterns[48235] = 29'b1_011110001101_011_1_111000110110;
      patterns[48236] = 29'b1_011110001101_100_1_101111000110;
      patterns[48237] = 29'b1_011110001101_101_0_110111100011;
      patterns[48238] = 29'b1_011110001101_110_1_011110001101;
      patterns[48239] = 29'b1_011110001101_111_1_011110001101;
      patterns[48240] = 29'b1_011110001110_000_1_011110001110;
      patterns[48241] = 29'b1_011110001110_001_1_001110011110;
      patterns[48242] = 29'b1_011110001110_010_0_111100011101;
      patterns[48243] = 29'b1_011110001110_011_1_111000111010;
      patterns[48244] = 29'b1_011110001110_100_0_101111000111;
      patterns[48245] = 29'b1_011110001110_101_1_010111100011;
      patterns[48246] = 29'b1_011110001110_110_1_011110001110;
      patterns[48247] = 29'b1_011110001110_111_1_011110001110;
      patterns[48248] = 29'b1_011110001111_000_1_011110001111;
      patterns[48249] = 29'b1_011110001111_001_1_001111011110;
      patterns[48250] = 29'b1_011110001111_010_0_111100011111;
      patterns[48251] = 29'b1_011110001111_011_1_111000111110;
      patterns[48252] = 29'b1_011110001111_100_1_101111000111;
      patterns[48253] = 29'b1_011110001111_101_1_110111100011;
      patterns[48254] = 29'b1_011110001111_110_1_011110001111;
      patterns[48255] = 29'b1_011110001111_111_1_011110001111;
      patterns[48256] = 29'b1_011110010000_000_1_011110010000;
      patterns[48257] = 29'b1_011110010000_001_1_010000011110;
      patterns[48258] = 29'b1_011110010000_010_0_111100100001;
      patterns[48259] = 29'b1_011110010000_011_1_111001000010;
      patterns[48260] = 29'b1_011110010000_100_0_101111001000;
      patterns[48261] = 29'b1_011110010000_101_0_010111100100;
      patterns[48262] = 29'b1_011110010000_110_1_011110010000;
      patterns[48263] = 29'b1_011110010000_111_1_011110010000;
      patterns[48264] = 29'b1_011110010001_000_1_011110010001;
      patterns[48265] = 29'b1_011110010001_001_1_010001011110;
      patterns[48266] = 29'b1_011110010001_010_0_111100100011;
      patterns[48267] = 29'b1_011110010001_011_1_111001000110;
      patterns[48268] = 29'b1_011110010001_100_1_101111001000;
      patterns[48269] = 29'b1_011110010001_101_0_110111100100;
      patterns[48270] = 29'b1_011110010001_110_1_011110010001;
      patterns[48271] = 29'b1_011110010001_111_1_011110010001;
      patterns[48272] = 29'b1_011110010010_000_1_011110010010;
      patterns[48273] = 29'b1_011110010010_001_1_010010011110;
      patterns[48274] = 29'b1_011110010010_010_0_111100100101;
      patterns[48275] = 29'b1_011110010010_011_1_111001001010;
      patterns[48276] = 29'b1_011110010010_100_0_101111001001;
      patterns[48277] = 29'b1_011110010010_101_1_010111100100;
      patterns[48278] = 29'b1_011110010010_110_1_011110010010;
      patterns[48279] = 29'b1_011110010010_111_1_011110010010;
      patterns[48280] = 29'b1_011110010011_000_1_011110010011;
      patterns[48281] = 29'b1_011110010011_001_1_010011011110;
      patterns[48282] = 29'b1_011110010011_010_0_111100100111;
      patterns[48283] = 29'b1_011110010011_011_1_111001001110;
      patterns[48284] = 29'b1_011110010011_100_1_101111001001;
      patterns[48285] = 29'b1_011110010011_101_1_110111100100;
      patterns[48286] = 29'b1_011110010011_110_1_011110010011;
      patterns[48287] = 29'b1_011110010011_111_1_011110010011;
      patterns[48288] = 29'b1_011110010100_000_1_011110010100;
      patterns[48289] = 29'b1_011110010100_001_1_010100011110;
      patterns[48290] = 29'b1_011110010100_010_0_111100101001;
      patterns[48291] = 29'b1_011110010100_011_1_111001010010;
      patterns[48292] = 29'b1_011110010100_100_0_101111001010;
      patterns[48293] = 29'b1_011110010100_101_0_010111100101;
      patterns[48294] = 29'b1_011110010100_110_1_011110010100;
      patterns[48295] = 29'b1_011110010100_111_1_011110010100;
      patterns[48296] = 29'b1_011110010101_000_1_011110010101;
      patterns[48297] = 29'b1_011110010101_001_1_010101011110;
      patterns[48298] = 29'b1_011110010101_010_0_111100101011;
      patterns[48299] = 29'b1_011110010101_011_1_111001010110;
      patterns[48300] = 29'b1_011110010101_100_1_101111001010;
      patterns[48301] = 29'b1_011110010101_101_0_110111100101;
      patterns[48302] = 29'b1_011110010101_110_1_011110010101;
      patterns[48303] = 29'b1_011110010101_111_1_011110010101;
      patterns[48304] = 29'b1_011110010110_000_1_011110010110;
      patterns[48305] = 29'b1_011110010110_001_1_010110011110;
      patterns[48306] = 29'b1_011110010110_010_0_111100101101;
      patterns[48307] = 29'b1_011110010110_011_1_111001011010;
      patterns[48308] = 29'b1_011110010110_100_0_101111001011;
      patterns[48309] = 29'b1_011110010110_101_1_010111100101;
      patterns[48310] = 29'b1_011110010110_110_1_011110010110;
      patterns[48311] = 29'b1_011110010110_111_1_011110010110;
      patterns[48312] = 29'b1_011110010111_000_1_011110010111;
      patterns[48313] = 29'b1_011110010111_001_1_010111011110;
      patterns[48314] = 29'b1_011110010111_010_0_111100101111;
      patterns[48315] = 29'b1_011110010111_011_1_111001011110;
      patterns[48316] = 29'b1_011110010111_100_1_101111001011;
      patterns[48317] = 29'b1_011110010111_101_1_110111100101;
      patterns[48318] = 29'b1_011110010111_110_1_011110010111;
      patterns[48319] = 29'b1_011110010111_111_1_011110010111;
      patterns[48320] = 29'b1_011110011000_000_1_011110011000;
      patterns[48321] = 29'b1_011110011000_001_1_011000011110;
      patterns[48322] = 29'b1_011110011000_010_0_111100110001;
      patterns[48323] = 29'b1_011110011000_011_1_111001100010;
      patterns[48324] = 29'b1_011110011000_100_0_101111001100;
      patterns[48325] = 29'b1_011110011000_101_0_010111100110;
      patterns[48326] = 29'b1_011110011000_110_1_011110011000;
      patterns[48327] = 29'b1_011110011000_111_1_011110011000;
      patterns[48328] = 29'b1_011110011001_000_1_011110011001;
      patterns[48329] = 29'b1_011110011001_001_1_011001011110;
      patterns[48330] = 29'b1_011110011001_010_0_111100110011;
      patterns[48331] = 29'b1_011110011001_011_1_111001100110;
      patterns[48332] = 29'b1_011110011001_100_1_101111001100;
      patterns[48333] = 29'b1_011110011001_101_0_110111100110;
      patterns[48334] = 29'b1_011110011001_110_1_011110011001;
      patterns[48335] = 29'b1_011110011001_111_1_011110011001;
      patterns[48336] = 29'b1_011110011010_000_1_011110011010;
      patterns[48337] = 29'b1_011110011010_001_1_011010011110;
      patterns[48338] = 29'b1_011110011010_010_0_111100110101;
      patterns[48339] = 29'b1_011110011010_011_1_111001101010;
      patterns[48340] = 29'b1_011110011010_100_0_101111001101;
      patterns[48341] = 29'b1_011110011010_101_1_010111100110;
      patterns[48342] = 29'b1_011110011010_110_1_011110011010;
      patterns[48343] = 29'b1_011110011010_111_1_011110011010;
      patterns[48344] = 29'b1_011110011011_000_1_011110011011;
      patterns[48345] = 29'b1_011110011011_001_1_011011011110;
      patterns[48346] = 29'b1_011110011011_010_0_111100110111;
      patterns[48347] = 29'b1_011110011011_011_1_111001101110;
      patterns[48348] = 29'b1_011110011011_100_1_101111001101;
      patterns[48349] = 29'b1_011110011011_101_1_110111100110;
      patterns[48350] = 29'b1_011110011011_110_1_011110011011;
      patterns[48351] = 29'b1_011110011011_111_1_011110011011;
      patterns[48352] = 29'b1_011110011100_000_1_011110011100;
      patterns[48353] = 29'b1_011110011100_001_1_011100011110;
      patterns[48354] = 29'b1_011110011100_010_0_111100111001;
      patterns[48355] = 29'b1_011110011100_011_1_111001110010;
      patterns[48356] = 29'b1_011110011100_100_0_101111001110;
      patterns[48357] = 29'b1_011110011100_101_0_010111100111;
      patterns[48358] = 29'b1_011110011100_110_1_011110011100;
      patterns[48359] = 29'b1_011110011100_111_1_011110011100;
      patterns[48360] = 29'b1_011110011101_000_1_011110011101;
      patterns[48361] = 29'b1_011110011101_001_1_011101011110;
      patterns[48362] = 29'b1_011110011101_010_0_111100111011;
      patterns[48363] = 29'b1_011110011101_011_1_111001110110;
      patterns[48364] = 29'b1_011110011101_100_1_101111001110;
      patterns[48365] = 29'b1_011110011101_101_0_110111100111;
      patterns[48366] = 29'b1_011110011101_110_1_011110011101;
      patterns[48367] = 29'b1_011110011101_111_1_011110011101;
      patterns[48368] = 29'b1_011110011110_000_1_011110011110;
      patterns[48369] = 29'b1_011110011110_001_1_011110011110;
      patterns[48370] = 29'b1_011110011110_010_0_111100111101;
      patterns[48371] = 29'b1_011110011110_011_1_111001111010;
      patterns[48372] = 29'b1_011110011110_100_0_101111001111;
      patterns[48373] = 29'b1_011110011110_101_1_010111100111;
      patterns[48374] = 29'b1_011110011110_110_1_011110011110;
      patterns[48375] = 29'b1_011110011110_111_1_011110011110;
      patterns[48376] = 29'b1_011110011111_000_1_011110011111;
      patterns[48377] = 29'b1_011110011111_001_1_011111011110;
      patterns[48378] = 29'b1_011110011111_010_0_111100111111;
      patterns[48379] = 29'b1_011110011111_011_1_111001111110;
      patterns[48380] = 29'b1_011110011111_100_1_101111001111;
      patterns[48381] = 29'b1_011110011111_101_1_110111100111;
      patterns[48382] = 29'b1_011110011111_110_1_011110011111;
      patterns[48383] = 29'b1_011110011111_111_1_011110011111;
      patterns[48384] = 29'b1_011110100000_000_1_011110100000;
      patterns[48385] = 29'b1_011110100000_001_1_100000011110;
      patterns[48386] = 29'b1_011110100000_010_0_111101000001;
      patterns[48387] = 29'b1_011110100000_011_1_111010000010;
      patterns[48388] = 29'b1_011110100000_100_0_101111010000;
      patterns[48389] = 29'b1_011110100000_101_0_010111101000;
      patterns[48390] = 29'b1_011110100000_110_1_011110100000;
      patterns[48391] = 29'b1_011110100000_111_1_011110100000;
      patterns[48392] = 29'b1_011110100001_000_1_011110100001;
      patterns[48393] = 29'b1_011110100001_001_1_100001011110;
      patterns[48394] = 29'b1_011110100001_010_0_111101000011;
      patterns[48395] = 29'b1_011110100001_011_1_111010000110;
      patterns[48396] = 29'b1_011110100001_100_1_101111010000;
      patterns[48397] = 29'b1_011110100001_101_0_110111101000;
      patterns[48398] = 29'b1_011110100001_110_1_011110100001;
      patterns[48399] = 29'b1_011110100001_111_1_011110100001;
      patterns[48400] = 29'b1_011110100010_000_1_011110100010;
      patterns[48401] = 29'b1_011110100010_001_1_100010011110;
      patterns[48402] = 29'b1_011110100010_010_0_111101000101;
      patterns[48403] = 29'b1_011110100010_011_1_111010001010;
      patterns[48404] = 29'b1_011110100010_100_0_101111010001;
      patterns[48405] = 29'b1_011110100010_101_1_010111101000;
      patterns[48406] = 29'b1_011110100010_110_1_011110100010;
      patterns[48407] = 29'b1_011110100010_111_1_011110100010;
      patterns[48408] = 29'b1_011110100011_000_1_011110100011;
      patterns[48409] = 29'b1_011110100011_001_1_100011011110;
      patterns[48410] = 29'b1_011110100011_010_0_111101000111;
      patterns[48411] = 29'b1_011110100011_011_1_111010001110;
      patterns[48412] = 29'b1_011110100011_100_1_101111010001;
      patterns[48413] = 29'b1_011110100011_101_1_110111101000;
      patterns[48414] = 29'b1_011110100011_110_1_011110100011;
      patterns[48415] = 29'b1_011110100011_111_1_011110100011;
      patterns[48416] = 29'b1_011110100100_000_1_011110100100;
      patterns[48417] = 29'b1_011110100100_001_1_100100011110;
      patterns[48418] = 29'b1_011110100100_010_0_111101001001;
      patterns[48419] = 29'b1_011110100100_011_1_111010010010;
      patterns[48420] = 29'b1_011110100100_100_0_101111010010;
      patterns[48421] = 29'b1_011110100100_101_0_010111101001;
      patterns[48422] = 29'b1_011110100100_110_1_011110100100;
      patterns[48423] = 29'b1_011110100100_111_1_011110100100;
      patterns[48424] = 29'b1_011110100101_000_1_011110100101;
      patterns[48425] = 29'b1_011110100101_001_1_100101011110;
      patterns[48426] = 29'b1_011110100101_010_0_111101001011;
      patterns[48427] = 29'b1_011110100101_011_1_111010010110;
      patterns[48428] = 29'b1_011110100101_100_1_101111010010;
      patterns[48429] = 29'b1_011110100101_101_0_110111101001;
      patterns[48430] = 29'b1_011110100101_110_1_011110100101;
      patterns[48431] = 29'b1_011110100101_111_1_011110100101;
      patterns[48432] = 29'b1_011110100110_000_1_011110100110;
      patterns[48433] = 29'b1_011110100110_001_1_100110011110;
      patterns[48434] = 29'b1_011110100110_010_0_111101001101;
      patterns[48435] = 29'b1_011110100110_011_1_111010011010;
      patterns[48436] = 29'b1_011110100110_100_0_101111010011;
      patterns[48437] = 29'b1_011110100110_101_1_010111101001;
      patterns[48438] = 29'b1_011110100110_110_1_011110100110;
      patterns[48439] = 29'b1_011110100110_111_1_011110100110;
      patterns[48440] = 29'b1_011110100111_000_1_011110100111;
      patterns[48441] = 29'b1_011110100111_001_1_100111011110;
      patterns[48442] = 29'b1_011110100111_010_0_111101001111;
      patterns[48443] = 29'b1_011110100111_011_1_111010011110;
      patterns[48444] = 29'b1_011110100111_100_1_101111010011;
      patterns[48445] = 29'b1_011110100111_101_1_110111101001;
      patterns[48446] = 29'b1_011110100111_110_1_011110100111;
      patterns[48447] = 29'b1_011110100111_111_1_011110100111;
      patterns[48448] = 29'b1_011110101000_000_1_011110101000;
      patterns[48449] = 29'b1_011110101000_001_1_101000011110;
      patterns[48450] = 29'b1_011110101000_010_0_111101010001;
      patterns[48451] = 29'b1_011110101000_011_1_111010100010;
      patterns[48452] = 29'b1_011110101000_100_0_101111010100;
      patterns[48453] = 29'b1_011110101000_101_0_010111101010;
      patterns[48454] = 29'b1_011110101000_110_1_011110101000;
      patterns[48455] = 29'b1_011110101000_111_1_011110101000;
      patterns[48456] = 29'b1_011110101001_000_1_011110101001;
      patterns[48457] = 29'b1_011110101001_001_1_101001011110;
      patterns[48458] = 29'b1_011110101001_010_0_111101010011;
      patterns[48459] = 29'b1_011110101001_011_1_111010100110;
      patterns[48460] = 29'b1_011110101001_100_1_101111010100;
      patterns[48461] = 29'b1_011110101001_101_0_110111101010;
      patterns[48462] = 29'b1_011110101001_110_1_011110101001;
      patterns[48463] = 29'b1_011110101001_111_1_011110101001;
      patterns[48464] = 29'b1_011110101010_000_1_011110101010;
      patterns[48465] = 29'b1_011110101010_001_1_101010011110;
      patterns[48466] = 29'b1_011110101010_010_0_111101010101;
      patterns[48467] = 29'b1_011110101010_011_1_111010101010;
      patterns[48468] = 29'b1_011110101010_100_0_101111010101;
      patterns[48469] = 29'b1_011110101010_101_1_010111101010;
      patterns[48470] = 29'b1_011110101010_110_1_011110101010;
      patterns[48471] = 29'b1_011110101010_111_1_011110101010;
      patterns[48472] = 29'b1_011110101011_000_1_011110101011;
      patterns[48473] = 29'b1_011110101011_001_1_101011011110;
      patterns[48474] = 29'b1_011110101011_010_0_111101010111;
      patterns[48475] = 29'b1_011110101011_011_1_111010101110;
      patterns[48476] = 29'b1_011110101011_100_1_101111010101;
      patterns[48477] = 29'b1_011110101011_101_1_110111101010;
      patterns[48478] = 29'b1_011110101011_110_1_011110101011;
      patterns[48479] = 29'b1_011110101011_111_1_011110101011;
      patterns[48480] = 29'b1_011110101100_000_1_011110101100;
      patterns[48481] = 29'b1_011110101100_001_1_101100011110;
      patterns[48482] = 29'b1_011110101100_010_0_111101011001;
      patterns[48483] = 29'b1_011110101100_011_1_111010110010;
      patterns[48484] = 29'b1_011110101100_100_0_101111010110;
      patterns[48485] = 29'b1_011110101100_101_0_010111101011;
      patterns[48486] = 29'b1_011110101100_110_1_011110101100;
      patterns[48487] = 29'b1_011110101100_111_1_011110101100;
      patterns[48488] = 29'b1_011110101101_000_1_011110101101;
      patterns[48489] = 29'b1_011110101101_001_1_101101011110;
      patterns[48490] = 29'b1_011110101101_010_0_111101011011;
      patterns[48491] = 29'b1_011110101101_011_1_111010110110;
      patterns[48492] = 29'b1_011110101101_100_1_101111010110;
      patterns[48493] = 29'b1_011110101101_101_0_110111101011;
      patterns[48494] = 29'b1_011110101101_110_1_011110101101;
      patterns[48495] = 29'b1_011110101101_111_1_011110101101;
      patterns[48496] = 29'b1_011110101110_000_1_011110101110;
      patterns[48497] = 29'b1_011110101110_001_1_101110011110;
      patterns[48498] = 29'b1_011110101110_010_0_111101011101;
      patterns[48499] = 29'b1_011110101110_011_1_111010111010;
      patterns[48500] = 29'b1_011110101110_100_0_101111010111;
      patterns[48501] = 29'b1_011110101110_101_1_010111101011;
      patterns[48502] = 29'b1_011110101110_110_1_011110101110;
      patterns[48503] = 29'b1_011110101110_111_1_011110101110;
      patterns[48504] = 29'b1_011110101111_000_1_011110101111;
      patterns[48505] = 29'b1_011110101111_001_1_101111011110;
      patterns[48506] = 29'b1_011110101111_010_0_111101011111;
      patterns[48507] = 29'b1_011110101111_011_1_111010111110;
      patterns[48508] = 29'b1_011110101111_100_1_101111010111;
      patterns[48509] = 29'b1_011110101111_101_1_110111101011;
      patterns[48510] = 29'b1_011110101111_110_1_011110101111;
      patterns[48511] = 29'b1_011110101111_111_1_011110101111;
      patterns[48512] = 29'b1_011110110000_000_1_011110110000;
      patterns[48513] = 29'b1_011110110000_001_1_110000011110;
      patterns[48514] = 29'b1_011110110000_010_0_111101100001;
      patterns[48515] = 29'b1_011110110000_011_1_111011000010;
      patterns[48516] = 29'b1_011110110000_100_0_101111011000;
      patterns[48517] = 29'b1_011110110000_101_0_010111101100;
      patterns[48518] = 29'b1_011110110000_110_1_011110110000;
      patterns[48519] = 29'b1_011110110000_111_1_011110110000;
      patterns[48520] = 29'b1_011110110001_000_1_011110110001;
      patterns[48521] = 29'b1_011110110001_001_1_110001011110;
      patterns[48522] = 29'b1_011110110001_010_0_111101100011;
      patterns[48523] = 29'b1_011110110001_011_1_111011000110;
      patterns[48524] = 29'b1_011110110001_100_1_101111011000;
      patterns[48525] = 29'b1_011110110001_101_0_110111101100;
      patterns[48526] = 29'b1_011110110001_110_1_011110110001;
      patterns[48527] = 29'b1_011110110001_111_1_011110110001;
      patterns[48528] = 29'b1_011110110010_000_1_011110110010;
      patterns[48529] = 29'b1_011110110010_001_1_110010011110;
      patterns[48530] = 29'b1_011110110010_010_0_111101100101;
      patterns[48531] = 29'b1_011110110010_011_1_111011001010;
      patterns[48532] = 29'b1_011110110010_100_0_101111011001;
      patterns[48533] = 29'b1_011110110010_101_1_010111101100;
      patterns[48534] = 29'b1_011110110010_110_1_011110110010;
      patterns[48535] = 29'b1_011110110010_111_1_011110110010;
      patterns[48536] = 29'b1_011110110011_000_1_011110110011;
      patterns[48537] = 29'b1_011110110011_001_1_110011011110;
      patterns[48538] = 29'b1_011110110011_010_0_111101100111;
      patterns[48539] = 29'b1_011110110011_011_1_111011001110;
      patterns[48540] = 29'b1_011110110011_100_1_101111011001;
      patterns[48541] = 29'b1_011110110011_101_1_110111101100;
      patterns[48542] = 29'b1_011110110011_110_1_011110110011;
      patterns[48543] = 29'b1_011110110011_111_1_011110110011;
      patterns[48544] = 29'b1_011110110100_000_1_011110110100;
      patterns[48545] = 29'b1_011110110100_001_1_110100011110;
      patterns[48546] = 29'b1_011110110100_010_0_111101101001;
      patterns[48547] = 29'b1_011110110100_011_1_111011010010;
      patterns[48548] = 29'b1_011110110100_100_0_101111011010;
      patterns[48549] = 29'b1_011110110100_101_0_010111101101;
      patterns[48550] = 29'b1_011110110100_110_1_011110110100;
      patterns[48551] = 29'b1_011110110100_111_1_011110110100;
      patterns[48552] = 29'b1_011110110101_000_1_011110110101;
      patterns[48553] = 29'b1_011110110101_001_1_110101011110;
      patterns[48554] = 29'b1_011110110101_010_0_111101101011;
      patterns[48555] = 29'b1_011110110101_011_1_111011010110;
      patterns[48556] = 29'b1_011110110101_100_1_101111011010;
      patterns[48557] = 29'b1_011110110101_101_0_110111101101;
      patterns[48558] = 29'b1_011110110101_110_1_011110110101;
      patterns[48559] = 29'b1_011110110101_111_1_011110110101;
      patterns[48560] = 29'b1_011110110110_000_1_011110110110;
      patterns[48561] = 29'b1_011110110110_001_1_110110011110;
      patterns[48562] = 29'b1_011110110110_010_0_111101101101;
      patterns[48563] = 29'b1_011110110110_011_1_111011011010;
      patterns[48564] = 29'b1_011110110110_100_0_101111011011;
      patterns[48565] = 29'b1_011110110110_101_1_010111101101;
      patterns[48566] = 29'b1_011110110110_110_1_011110110110;
      patterns[48567] = 29'b1_011110110110_111_1_011110110110;
      patterns[48568] = 29'b1_011110110111_000_1_011110110111;
      patterns[48569] = 29'b1_011110110111_001_1_110111011110;
      patterns[48570] = 29'b1_011110110111_010_0_111101101111;
      patterns[48571] = 29'b1_011110110111_011_1_111011011110;
      patterns[48572] = 29'b1_011110110111_100_1_101111011011;
      patterns[48573] = 29'b1_011110110111_101_1_110111101101;
      patterns[48574] = 29'b1_011110110111_110_1_011110110111;
      patterns[48575] = 29'b1_011110110111_111_1_011110110111;
      patterns[48576] = 29'b1_011110111000_000_1_011110111000;
      patterns[48577] = 29'b1_011110111000_001_1_111000011110;
      patterns[48578] = 29'b1_011110111000_010_0_111101110001;
      patterns[48579] = 29'b1_011110111000_011_1_111011100010;
      patterns[48580] = 29'b1_011110111000_100_0_101111011100;
      patterns[48581] = 29'b1_011110111000_101_0_010111101110;
      patterns[48582] = 29'b1_011110111000_110_1_011110111000;
      patterns[48583] = 29'b1_011110111000_111_1_011110111000;
      patterns[48584] = 29'b1_011110111001_000_1_011110111001;
      patterns[48585] = 29'b1_011110111001_001_1_111001011110;
      patterns[48586] = 29'b1_011110111001_010_0_111101110011;
      patterns[48587] = 29'b1_011110111001_011_1_111011100110;
      patterns[48588] = 29'b1_011110111001_100_1_101111011100;
      patterns[48589] = 29'b1_011110111001_101_0_110111101110;
      patterns[48590] = 29'b1_011110111001_110_1_011110111001;
      patterns[48591] = 29'b1_011110111001_111_1_011110111001;
      patterns[48592] = 29'b1_011110111010_000_1_011110111010;
      patterns[48593] = 29'b1_011110111010_001_1_111010011110;
      patterns[48594] = 29'b1_011110111010_010_0_111101110101;
      patterns[48595] = 29'b1_011110111010_011_1_111011101010;
      patterns[48596] = 29'b1_011110111010_100_0_101111011101;
      patterns[48597] = 29'b1_011110111010_101_1_010111101110;
      patterns[48598] = 29'b1_011110111010_110_1_011110111010;
      patterns[48599] = 29'b1_011110111010_111_1_011110111010;
      patterns[48600] = 29'b1_011110111011_000_1_011110111011;
      patterns[48601] = 29'b1_011110111011_001_1_111011011110;
      patterns[48602] = 29'b1_011110111011_010_0_111101110111;
      patterns[48603] = 29'b1_011110111011_011_1_111011101110;
      patterns[48604] = 29'b1_011110111011_100_1_101111011101;
      patterns[48605] = 29'b1_011110111011_101_1_110111101110;
      patterns[48606] = 29'b1_011110111011_110_1_011110111011;
      patterns[48607] = 29'b1_011110111011_111_1_011110111011;
      patterns[48608] = 29'b1_011110111100_000_1_011110111100;
      patterns[48609] = 29'b1_011110111100_001_1_111100011110;
      patterns[48610] = 29'b1_011110111100_010_0_111101111001;
      patterns[48611] = 29'b1_011110111100_011_1_111011110010;
      patterns[48612] = 29'b1_011110111100_100_0_101111011110;
      patterns[48613] = 29'b1_011110111100_101_0_010111101111;
      patterns[48614] = 29'b1_011110111100_110_1_011110111100;
      patterns[48615] = 29'b1_011110111100_111_1_011110111100;
      patterns[48616] = 29'b1_011110111101_000_1_011110111101;
      patterns[48617] = 29'b1_011110111101_001_1_111101011110;
      patterns[48618] = 29'b1_011110111101_010_0_111101111011;
      patterns[48619] = 29'b1_011110111101_011_1_111011110110;
      patterns[48620] = 29'b1_011110111101_100_1_101111011110;
      patterns[48621] = 29'b1_011110111101_101_0_110111101111;
      patterns[48622] = 29'b1_011110111101_110_1_011110111101;
      patterns[48623] = 29'b1_011110111101_111_1_011110111101;
      patterns[48624] = 29'b1_011110111110_000_1_011110111110;
      patterns[48625] = 29'b1_011110111110_001_1_111110011110;
      patterns[48626] = 29'b1_011110111110_010_0_111101111101;
      patterns[48627] = 29'b1_011110111110_011_1_111011111010;
      patterns[48628] = 29'b1_011110111110_100_0_101111011111;
      patterns[48629] = 29'b1_011110111110_101_1_010111101111;
      patterns[48630] = 29'b1_011110111110_110_1_011110111110;
      patterns[48631] = 29'b1_011110111110_111_1_011110111110;
      patterns[48632] = 29'b1_011110111111_000_1_011110111111;
      patterns[48633] = 29'b1_011110111111_001_1_111111011110;
      patterns[48634] = 29'b1_011110111111_010_0_111101111111;
      patterns[48635] = 29'b1_011110111111_011_1_111011111110;
      patterns[48636] = 29'b1_011110111111_100_1_101111011111;
      patterns[48637] = 29'b1_011110111111_101_1_110111101111;
      patterns[48638] = 29'b1_011110111111_110_1_011110111111;
      patterns[48639] = 29'b1_011110111111_111_1_011110111111;
      patterns[48640] = 29'b1_011111000000_000_1_011111000000;
      patterns[48641] = 29'b1_011111000000_001_1_000000011111;
      patterns[48642] = 29'b1_011111000000_010_0_111110000001;
      patterns[48643] = 29'b1_011111000000_011_1_111100000010;
      patterns[48644] = 29'b1_011111000000_100_0_101111100000;
      patterns[48645] = 29'b1_011111000000_101_0_010111110000;
      patterns[48646] = 29'b1_011111000000_110_1_011111000000;
      patterns[48647] = 29'b1_011111000000_111_1_011111000000;
      patterns[48648] = 29'b1_011111000001_000_1_011111000001;
      patterns[48649] = 29'b1_011111000001_001_1_000001011111;
      patterns[48650] = 29'b1_011111000001_010_0_111110000011;
      patterns[48651] = 29'b1_011111000001_011_1_111100000110;
      patterns[48652] = 29'b1_011111000001_100_1_101111100000;
      patterns[48653] = 29'b1_011111000001_101_0_110111110000;
      patterns[48654] = 29'b1_011111000001_110_1_011111000001;
      patterns[48655] = 29'b1_011111000001_111_1_011111000001;
      patterns[48656] = 29'b1_011111000010_000_1_011111000010;
      patterns[48657] = 29'b1_011111000010_001_1_000010011111;
      patterns[48658] = 29'b1_011111000010_010_0_111110000101;
      patterns[48659] = 29'b1_011111000010_011_1_111100001010;
      patterns[48660] = 29'b1_011111000010_100_0_101111100001;
      patterns[48661] = 29'b1_011111000010_101_1_010111110000;
      patterns[48662] = 29'b1_011111000010_110_1_011111000010;
      patterns[48663] = 29'b1_011111000010_111_1_011111000010;
      patterns[48664] = 29'b1_011111000011_000_1_011111000011;
      patterns[48665] = 29'b1_011111000011_001_1_000011011111;
      patterns[48666] = 29'b1_011111000011_010_0_111110000111;
      patterns[48667] = 29'b1_011111000011_011_1_111100001110;
      patterns[48668] = 29'b1_011111000011_100_1_101111100001;
      patterns[48669] = 29'b1_011111000011_101_1_110111110000;
      patterns[48670] = 29'b1_011111000011_110_1_011111000011;
      patterns[48671] = 29'b1_011111000011_111_1_011111000011;
      patterns[48672] = 29'b1_011111000100_000_1_011111000100;
      patterns[48673] = 29'b1_011111000100_001_1_000100011111;
      patterns[48674] = 29'b1_011111000100_010_0_111110001001;
      patterns[48675] = 29'b1_011111000100_011_1_111100010010;
      patterns[48676] = 29'b1_011111000100_100_0_101111100010;
      patterns[48677] = 29'b1_011111000100_101_0_010111110001;
      patterns[48678] = 29'b1_011111000100_110_1_011111000100;
      patterns[48679] = 29'b1_011111000100_111_1_011111000100;
      patterns[48680] = 29'b1_011111000101_000_1_011111000101;
      patterns[48681] = 29'b1_011111000101_001_1_000101011111;
      patterns[48682] = 29'b1_011111000101_010_0_111110001011;
      patterns[48683] = 29'b1_011111000101_011_1_111100010110;
      patterns[48684] = 29'b1_011111000101_100_1_101111100010;
      patterns[48685] = 29'b1_011111000101_101_0_110111110001;
      patterns[48686] = 29'b1_011111000101_110_1_011111000101;
      patterns[48687] = 29'b1_011111000101_111_1_011111000101;
      patterns[48688] = 29'b1_011111000110_000_1_011111000110;
      patterns[48689] = 29'b1_011111000110_001_1_000110011111;
      patterns[48690] = 29'b1_011111000110_010_0_111110001101;
      patterns[48691] = 29'b1_011111000110_011_1_111100011010;
      patterns[48692] = 29'b1_011111000110_100_0_101111100011;
      patterns[48693] = 29'b1_011111000110_101_1_010111110001;
      patterns[48694] = 29'b1_011111000110_110_1_011111000110;
      patterns[48695] = 29'b1_011111000110_111_1_011111000110;
      patterns[48696] = 29'b1_011111000111_000_1_011111000111;
      patterns[48697] = 29'b1_011111000111_001_1_000111011111;
      patterns[48698] = 29'b1_011111000111_010_0_111110001111;
      patterns[48699] = 29'b1_011111000111_011_1_111100011110;
      patterns[48700] = 29'b1_011111000111_100_1_101111100011;
      patterns[48701] = 29'b1_011111000111_101_1_110111110001;
      patterns[48702] = 29'b1_011111000111_110_1_011111000111;
      patterns[48703] = 29'b1_011111000111_111_1_011111000111;
      patterns[48704] = 29'b1_011111001000_000_1_011111001000;
      patterns[48705] = 29'b1_011111001000_001_1_001000011111;
      patterns[48706] = 29'b1_011111001000_010_0_111110010001;
      patterns[48707] = 29'b1_011111001000_011_1_111100100010;
      patterns[48708] = 29'b1_011111001000_100_0_101111100100;
      patterns[48709] = 29'b1_011111001000_101_0_010111110010;
      patterns[48710] = 29'b1_011111001000_110_1_011111001000;
      patterns[48711] = 29'b1_011111001000_111_1_011111001000;
      patterns[48712] = 29'b1_011111001001_000_1_011111001001;
      patterns[48713] = 29'b1_011111001001_001_1_001001011111;
      patterns[48714] = 29'b1_011111001001_010_0_111110010011;
      patterns[48715] = 29'b1_011111001001_011_1_111100100110;
      patterns[48716] = 29'b1_011111001001_100_1_101111100100;
      patterns[48717] = 29'b1_011111001001_101_0_110111110010;
      patterns[48718] = 29'b1_011111001001_110_1_011111001001;
      patterns[48719] = 29'b1_011111001001_111_1_011111001001;
      patterns[48720] = 29'b1_011111001010_000_1_011111001010;
      patterns[48721] = 29'b1_011111001010_001_1_001010011111;
      patterns[48722] = 29'b1_011111001010_010_0_111110010101;
      patterns[48723] = 29'b1_011111001010_011_1_111100101010;
      patterns[48724] = 29'b1_011111001010_100_0_101111100101;
      patterns[48725] = 29'b1_011111001010_101_1_010111110010;
      patterns[48726] = 29'b1_011111001010_110_1_011111001010;
      patterns[48727] = 29'b1_011111001010_111_1_011111001010;
      patterns[48728] = 29'b1_011111001011_000_1_011111001011;
      patterns[48729] = 29'b1_011111001011_001_1_001011011111;
      patterns[48730] = 29'b1_011111001011_010_0_111110010111;
      patterns[48731] = 29'b1_011111001011_011_1_111100101110;
      patterns[48732] = 29'b1_011111001011_100_1_101111100101;
      patterns[48733] = 29'b1_011111001011_101_1_110111110010;
      patterns[48734] = 29'b1_011111001011_110_1_011111001011;
      patterns[48735] = 29'b1_011111001011_111_1_011111001011;
      patterns[48736] = 29'b1_011111001100_000_1_011111001100;
      patterns[48737] = 29'b1_011111001100_001_1_001100011111;
      patterns[48738] = 29'b1_011111001100_010_0_111110011001;
      patterns[48739] = 29'b1_011111001100_011_1_111100110010;
      patterns[48740] = 29'b1_011111001100_100_0_101111100110;
      patterns[48741] = 29'b1_011111001100_101_0_010111110011;
      patterns[48742] = 29'b1_011111001100_110_1_011111001100;
      patterns[48743] = 29'b1_011111001100_111_1_011111001100;
      patterns[48744] = 29'b1_011111001101_000_1_011111001101;
      patterns[48745] = 29'b1_011111001101_001_1_001101011111;
      patterns[48746] = 29'b1_011111001101_010_0_111110011011;
      patterns[48747] = 29'b1_011111001101_011_1_111100110110;
      patterns[48748] = 29'b1_011111001101_100_1_101111100110;
      patterns[48749] = 29'b1_011111001101_101_0_110111110011;
      patterns[48750] = 29'b1_011111001101_110_1_011111001101;
      patterns[48751] = 29'b1_011111001101_111_1_011111001101;
      patterns[48752] = 29'b1_011111001110_000_1_011111001110;
      patterns[48753] = 29'b1_011111001110_001_1_001110011111;
      patterns[48754] = 29'b1_011111001110_010_0_111110011101;
      patterns[48755] = 29'b1_011111001110_011_1_111100111010;
      patterns[48756] = 29'b1_011111001110_100_0_101111100111;
      patterns[48757] = 29'b1_011111001110_101_1_010111110011;
      patterns[48758] = 29'b1_011111001110_110_1_011111001110;
      patterns[48759] = 29'b1_011111001110_111_1_011111001110;
      patterns[48760] = 29'b1_011111001111_000_1_011111001111;
      patterns[48761] = 29'b1_011111001111_001_1_001111011111;
      patterns[48762] = 29'b1_011111001111_010_0_111110011111;
      patterns[48763] = 29'b1_011111001111_011_1_111100111110;
      patterns[48764] = 29'b1_011111001111_100_1_101111100111;
      patterns[48765] = 29'b1_011111001111_101_1_110111110011;
      patterns[48766] = 29'b1_011111001111_110_1_011111001111;
      patterns[48767] = 29'b1_011111001111_111_1_011111001111;
      patterns[48768] = 29'b1_011111010000_000_1_011111010000;
      patterns[48769] = 29'b1_011111010000_001_1_010000011111;
      patterns[48770] = 29'b1_011111010000_010_0_111110100001;
      patterns[48771] = 29'b1_011111010000_011_1_111101000010;
      patterns[48772] = 29'b1_011111010000_100_0_101111101000;
      patterns[48773] = 29'b1_011111010000_101_0_010111110100;
      patterns[48774] = 29'b1_011111010000_110_1_011111010000;
      patterns[48775] = 29'b1_011111010000_111_1_011111010000;
      patterns[48776] = 29'b1_011111010001_000_1_011111010001;
      patterns[48777] = 29'b1_011111010001_001_1_010001011111;
      patterns[48778] = 29'b1_011111010001_010_0_111110100011;
      patterns[48779] = 29'b1_011111010001_011_1_111101000110;
      patterns[48780] = 29'b1_011111010001_100_1_101111101000;
      patterns[48781] = 29'b1_011111010001_101_0_110111110100;
      patterns[48782] = 29'b1_011111010001_110_1_011111010001;
      patterns[48783] = 29'b1_011111010001_111_1_011111010001;
      patterns[48784] = 29'b1_011111010010_000_1_011111010010;
      patterns[48785] = 29'b1_011111010010_001_1_010010011111;
      patterns[48786] = 29'b1_011111010010_010_0_111110100101;
      patterns[48787] = 29'b1_011111010010_011_1_111101001010;
      patterns[48788] = 29'b1_011111010010_100_0_101111101001;
      patterns[48789] = 29'b1_011111010010_101_1_010111110100;
      patterns[48790] = 29'b1_011111010010_110_1_011111010010;
      patterns[48791] = 29'b1_011111010010_111_1_011111010010;
      patterns[48792] = 29'b1_011111010011_000_1_011111010011;
      patterns[48793] = 29'b1_011111010011_001_1_010011011111;
      patterns[48794] = 29'b1_011111010011_010_0_111110100111;
      patterns[48795] = 29'b1_011111010011_011_1_111101001110;
      patterns[48796] = 29'b1_011111010011_100_1_101111101001;
      patterns[48797] = 29'b1_011111010011_101_1_110111110100;
      patterns[48798] = 29'b1_011111010011_110_1_011111010011;
      patterns[48799] = 29'b1_011111010011_111_1_011111010011;
      patterns[48800] = 29'b1_011111010100_000_1_011111010100;
      patterns[48801] = 29'b1_011111010100_001_1_010100011111;
      patterns[48802] = 29'b1_011111010100_010_0_111110101001;
      patterns[48803] = 29'b1_011111010100_011_1_111101010010;
      patterns[48804] = 29'b1_011111010100_100_0_101111101010;
      patterns[48805] = 29'b1_011111010100_101_0_010111110101;
      patterns[48806] = 29'b1_011111010100_110_1_011111010100;
      patterns[48807] = 29'b1_011111010100_111_1_011111010100;
      patterns[48808] = 29'b1_011111010101_000_1_011111010101;
      patterns[48809] = 29'b1_011111010101_001_1_010101011111;
      patterns[48810] = 29'b1_011111010101_010_0_111110101011;
      patterns[48811] = 29'b1_011111010101_011_1_111101010110;
      patterns[48812] = 29'b1_011111010101_100_1_101111101010;
      patterns[48813] = 29'b1_011111010101_101_0_110111110101;
      patterns[48814] = 29'b1_011111010101_110_1_011111010101;
      patterns[48815] = 29'b1_011111010101_111_1_011111010101;
      patterns[48816] = 29'b1_011111010110_000_1_011111010110;
      patterns[48817] = 29'b1_011111010110_001_1_010110011111;
      patterns[48818] = 29'b1_011111010110_010_0_111110101101;
      patterns[48819] = 29'b1_011111010110_011_1_111101011010;
      patterns[48820] = 29'b1_011111010110_100_0_101111101011;
      patterns[48821] = 29'b1_011111010110_101_1_010111110101;
      patterns[48822] = 29'b1_011111010110_110_1_011111010110;
      patterns[48823] = 29'b1_011111010110_111_1_011111010110;
      patterns[48824] = 29'b1_011111010111_000_1_011111010111;
      patterns[48825] = 29'b1_011111010111_001_1_010111011111;
      patterns[48826] = 29'b1_011111010111_010_0_111110101111;
      patterns[48827] = 29'b1_011111010111_011_1_111101011110;
      patterns[48828] = 29'b1_011111010111_100_1_101111101011;
      patterns[48829] = 29'b1_011111010111_101_1_110111110101;
      patterns[48830] = 29'b1_011111010111_110_1_011111010111;
      patterns[48831] = 29'b1_011111010111_111_1_011111010111;
      patterns[48832] = 29'b1_011111011000_000_1_011111011000;
      patterns[48833] = 29'b1_011111011000_001_1_011000011111;
      patterns[48834] = 29'b1_011111011000_010_0_111110110001;
      patterns[48835] = 29'b1_011111011000_011_1_111101100010;
      patterns[48836] = 29'b1_011111011000_100_0_101111101100;
      patterns[48837] = 29'b1_011111011000_101_0_010111110110;
      patterns[48838] = 29'b1_011111011000_110_1_011111011000;
      patterns[48839] = 29'b1_011111011000_111_1_011111011000;
      patterns[48840] = 29'b1_011111011001_000_1_011111011001;
      patterns[48841] = 29'b1_011111011001_001_1_011001011111;
      patterns[48842] = 29'b1_011111011001_010_0_111110110011;
      patterns[48843] = 29'b1_011111011001_011_1_111101100110;
      patterns[48844] = 29'b1_011111011001_100_1_101111101100;
      patterns[48845] = 29'b1_011111011001_101_0_110111110110;
      patterns[48846] = 29'b1_011111011001_110_1_011111011001;
      patterns[48847] = 29'b1_011111011001_111_1_011111011001;
      patterns[48848] = 29'b1_011111011010_000_1_011111011010;
      patterns[48849] = 29'b1_011111011010_001_1_011010011111;
      patterns[48850] = 29'b1_011111011010_010_0_111110110101;
      patterns[48851] = 29'b1_011111011010_011_1_111101101010;
      patterns[48852] = 29'b1_011111011010_100_0_101111101101;
      patterns[48853] = 29'b1_011111011010_101_1_010111110110;
      patterns[48854] = 29'b1_011111011010_110_1_011111011010;
      patterns[48855] = 29'b1_011111011010_111_1_011111011010;
      patterns[48856] = 29'b1_011111011011_000_1_011111011011;
      patterns[48857] = 29'b1_011111011011_001_1_011011011111;
      patterns[48858] = 29'b1_011111011011_010_0_111110110111;
      patterns[48859] = 29'b1_011111011011_011_1_111101101110;
      patterns[48860] = 29'b1_011111011011_100_1_101111101101;
      patterns[48861] = 29'b1_011111011011_101_1_110111110110;
      patterns[48862] = 29'b1_011111011011_110_1_011111011011;
      patterns[48863] = 29'b1_011111011011_111_1_011111011011;
      patterns[48864] = 29'b1_011111011100_000_1_011111011100;
      patterns[48865] = 29'b1_011111011100_001_1_011100011111;
      patterns[48866] = 29'b1_011111011100_010_0_111110111001;
      patterns[48867] = 29'b1_011111011100_011_1_111101110010;
      patterns[48868] = 29'b1_011111011100_100_0_101111101110;
      patterns[48869] = 29'b1_011111011100_101_0_010111110111;
      patterns[48870] = 29'b1_011111011100_110_1_011111011100;
      patterns[48871] = 29'b1_011111011100_111_1_011111011100;
      patterns[48872] = 29'b1_011111011101_000_1_011111011101;
      patterns[48873] = 29'b1_011111011101_001_1_011101011111;
      patterns[48874] = 29'b1_011111011101_010_0_111110111011;
      patterns[48875] = 29'b1_011111011101_011_1_111101110110;
      patterns[48876] = 29'b1_011111011101_100_1_101111101110;
      patterns[48877] = 29'b1_011111011101_101_0_110111110111;
      patterns[48878] = 29'b1_011111011101_110_1_011111011101;
      patterns[48879] = 29'b1_011111011101_111_1_011111011101;
      patterns[48880] = 29'b1_011111011110_000_1_011111011110;
      patterns[48881] = 29'b1_011111011110_001_1_011110011111;
      patterns[48882] = 29'b1_011111011110_010_0_111110111101;
      patterns[48883] = 29'b1_011111011110_011_1_111101111010;
      patterns[48884] = 29'b1_011111011110_100_0_101111101111;
      patterns[48885] = 29'b1_011111011110_101_1_010111110111;
      patterns[48886] = 29'b1_011111011110_110_1_011111011110;
      patterns[48887] = 29'b1_011111011110_111_1_011111011110;
      patterns[48888] = 29'b1_011111011111_000_1_011111011111;
      patterns[48889] = 29'b1_011111011111_001_1_011111011111;
      patterns[48890] = 29'b1_011111011111_010_0_111110111111;
      patterns[48891] = 29'b1_011111011111_011_1_111101111110;
      patterns[48892] = 29'b1_011111011111_100_1_101111101111;
      patterns[48893] = 29'b1_011111011111_101_1_110111110111;
      patterns[48894] = 29'b1_011111011111_110_1_011111011111;
      patterns[48895] = 29'b1_011111011111_111_1_011111011111;
      patterns[48896] = 29'b1_011111100000_000_1_011111100000;
      patterns[48897] = 29'b1_011111100000_001_1_100000011111;
      patterns[48898] = 29'b1_011111100000_010_0_111111000001;
      patterns[48899] = 29'b1_011111100000_011_1_111110000010;
      patterns[48900] = 29'b1_011111100000_100_0_101111110000;
      patterns[48901] = 29'b1_011111100000_101_0_010111111000;
      patterns[48902] = 29'b1_011111100000_110_1_011111100000;
      patterns[48903] = 29'b1_011111100000_111_1_011111100000;
      patterns[48904] = 29'b1_011111100001_000_1_011111100001;
      patterns[48905] = 29'b1_011111100001_001_1_100001011111;
      patterns[48906] = 29'b1_011111100001_010_0_111111000011;
      patterns[48907] = 29'b1_011111100001_011_1_111110000110;
      patterns[48908] = 29'b1_011111100001_100_1_101111110000;
      patterns[48909] = 29'b1_011111100001_101_0_110111111000;
      patterns[48910] = 29'b1_011111100001_110_1_011111100001;
      patterns[48911] = 29'b1_011111100001_111_1_011111100001;
      patterns[48912] = 29'b1_011111100010_000_1_011111100010;
      patterns[48913] = 29'b1_011111100010_001_1_100010011111;
      patterns[48914] = 29'b1_011111100010_010_0_111111000101;
      patterns[48915] = 29'b1_011111100010_011_1_111110001010;
      patterns[48916] = 29'b1_011111100010_100_0_101111110001;
      patterns[48917] = 29'b1_011111100010_101_1_010111111000;
      patterns[48918] = 29'b1_011111100010_110_1_011111100010;
      patterns[48919] = 29'b1_011111100010_111_1_011111100010;
      patterns[48920] = 29'b1_011111100011_000_1_011111100011;
      patterns[48921] = 29'b1_011111100011_001_1_100011011111;
      patterns[48922] = 29'b1_011111100011_010_0_111111000111;
      patterns[48923] = 29'b1_011111100011_011_1_111110001110;
      patterns[48924] = 29'b1_011111100011_100_1_101111110001;
      patterns[48925] = 29'b1_011111100011_101_1_110111111000;
      patterns[48926] = 29'b1_011111100011_110_1_011111100011;
      patterns[48927] = 29'b1_011111100011_111_1_011111100011;
      patterns[48928] = 29'b1_011111100100_000_1_011111100100;
      patterns[48929] = 29'b1_011111100100_001_1_100100011111;
      patterns[48930] = 29'b1_011111100100_010_0_111111001001;
      patterns[48931] = 29'b1_011111100100_011_1_111110010010;
      patterns[48932] = 29'b1_011111100100_100_0_101111110010;
      patterns[48933] = 29'b1_011111100100_101_0_010111111001;
      patterns[48934] = 29'b1_011111100100_110_1_011111100100;
      patterns[48935] = 29'b1_011111100100_111_1_011111100100;
      patterns[48936] = 29'b1_011111100101_000_1_011111100101;
      patterns[48937] = 29'b1_011111100101_001_1_100101011111;
      patterns[48938] = 29'b1_011111100101_010_0_111111001011;
      patterns[48939] = 29'b1_011111100101_011_1_111110010110;
      patterns[48940] = 29'b1_011111100101_100_1_101111110010;
      patterns[48941] = 29'b1_011111100101_101_0_110111111001;
      patterns[48942] = 29'b1_011111100101_110_1_011111100101;
      patterns[48943] = 29'b1_011111100101_111_1_011111100101;
      patterns[48944] = 29'b1_011111100110_000_1_011111100110;
      patterns[48945] = 29'b1_011111100110_001_1_100110011111;
      patterns[48946] = 29'b1_011111100110_010_0_111111001101;
      patterns[48947] = 29'b1_011111100110_011_1_111110011010;
      patterns[48948] = 29'b1_011111100110_100_0_101111110011;
      patterns[48949] = 29'b1_011111100110_101_1_010111111001;
      patterns[48950] = 29'b1_011111100110_110_1_011111100110;
      patterns[48951] = 29'b1_011111100110_111_1_011111100110;
      patterns[48952] = 29'b1_011111100111_000_1_011111100111;
      patterns[48953] = 29'b1_011111100111_001_1_100111011111;
      patterns[48954] = 29'b1_011111100111_010_0_111111001111;
      patterns[48955] = 29'b1_011111100111_011_1_111110011110;
      patterns[48956] = 29'b1_011111100111_100_1_101111110011;
      patterns[48957] = 29'b1_011111100111_101_1_110111111001;
      patterns[48958] = 29'b1_011111100111_110_1_011111100111;
      patterns[48959] = 29'b1_011111100111_111_1_011111100111;
      patterns[48960] = 29'b1_011111101000_000_1_011111101000;
      patterns[48961] = 29'b1_011111101000_001_1_101000011111;
      patterns[48962] = 29'b1_011111101000_010_0_111111010001;
      patterns[48963] = 29'b1_011111101000_011_1_111110100010;
      patterns[48964] = 29'b1_011111101000_100_0_101111110100;
      patterns[48965] = 29'b1_011111101000_101_0_010111111010;
      patterns[48966] = 29'b1_011111101000_110_1_011111101000;
      patterns[48967] = 29'b1_011111101000_111_1_011111101000;
      patterns[48968] = 29'b1_011111101001_000_1_011111101001;
      patterns[48969] = 29'b1_011111101001_001_1_101001011111;
      patterns[48970] = 29'b1_011111101001_010_0_111111010011;
      patterns[48971] = 29'b1_011111101001_011_1_111110100110;
      patterns[48972] = 29'b1_011111101001_100_1_101111110100;
      patterns[48973] = 29'b1_011111101001_101_0_110111111010;
      patterns[48974] = 29'b1_011111101001_110_1_011111101001;
      patterns[48975] = 29'b1_011111101001_111_1_011111101001;
      patterns[48976] = 29'b1_011111101010_000_1_011111101010;
      patterns[48977] = 29'b1_011111101010_001_1_101010011111;
      patterns[48978] = 29'b1_011111101010_010_0_111111010101;
      patterns[48979] = 29'b1_011111101010_011_1_111110101010;
      patterns[48980] = 29'b1_011111101010_100_0_101111110101;
      patterns[48981] = 29'b1_011111101010_101_1_010111111010;
      patterns[48982] = 29'b1_011111101010_110_1_011111101010;
      patterns[48983] = 29'b1_011111101010_111_1_011111101010;
      patterns[48984] = 29'b1_011111101011_000_1_011111101011;
      patterns[48985] = 29'b1_011111101011_001_1_101011011111;
      patterns[48986] = 29'b1_011111101011_010_0_111111010111;
      patterns[48987] = 29'b1_011111101011_011_1_111110101110;
      patterns[48988] = 29'b1_011111101011_100_1_101111110101;
      patterns[48989] = 29'b1_011111101011_101_1_110111111010;
      patterns[48990] = 29'b1_011111101011_110_1_011111101011;
      patterns[48991] = 29'b1_011111101011_111_1_011111101011;
      patterns[48992] = 29'b1_011111101100_000_1_011111101100;
      patterns[48993] = 29'b1_011111101100_001_1_101100011111;
      patterns[48994] = 29'b1_011111101100_010_0_111111011001;
      patterns[48995] = 29'b1_011111101100_011_1_111110110010;
      patterns[48996] = 29'b1_011111101100_100_0_101111110110;
      patterns[48997] = 29'b1_011111101100_101_0_010111111011;
      patterns[48998] = 29'b1_011111101100_110_1_011111101100;
      patterns[48999] = 29'b1_011111101100_111_1_011111101100;
      patterns[49000] = 29'b1_011111101101_000_1_011111101101;
      patterns[49001] = 29'b1_011111101101_001_1_101101011111;
      patterns[49002] = 29'b1_011111101101_010_0_111111011011;
      patterns[49003] = 29'b1_011111101101_011_1_111110110110;
      patterns[49004] = 29'b1_011111101101_100_1_101111110110;
      patterns[49005] = 29'b1_011111101101_101_0_110111111011;
      patterns[49006] = 29'b1_011111101101_110_1_011111101101;
      patterns[49007] = 29'b1_011111101101_111_1_011111101101;
      patterns[49008] = 29'b1_011111101110_000_1_011111101110;
      patterns[49009] = 29'b1_011111101110_001_1_101110011111;
      patterns[49010] = 29'b1_011111101110_010_0_111111011101;
      patterns[49011] = 29'b1_011111101110_011_1_111110111010;
      patterns[49012] = 29'b1_011111101110_100_0_101111110111;
      patterns[49013] = 29'b1_011111101110_101_1_010111111011;
      patterns[49014] = 29'b1_011111101110_110_1_011111101110;
      patterns[49015] = 29'b1_011111101110_111_1_011111101110;
      patterns[49016] = 29'b1_011111101111_000_1_011111101111;
      patterns[49017] = 29'b1_011111101111_001_1_101111011111;
      patterns[49018] = 29'b1_011111101111_010_0_111111011111;
      patterns[49019] = 29'b1_011111101111_011_1_111110111110;
      patterns[49020] = 29'b1_011111101111_100_1_101111110111;
      patterns[49021] = 29'b1_011111101111_101_1_110111111011;
      patterns[49022] = 29'b1_011111101111_110_1_011111101111;
      patterns[49023] = 29'b1_011111101111_111_1_011111101111;
      patterns[49024] = 29'b1_011111110000_000_1_011111110000;
      patterns[49025] = 29'b1_011111110000_001_1_110000011111;
      patterns[49026] = 29'b1_011111110000_010_0_111111100001;
      patterns[49027] = 29'b1_011111110000_011_1_111111000010;
      patterns[49028] = 29'b1_011111110000_100_0_101111111000;
      patterns[49029] = 29'b1_011111110000_101_0_010111111100;
      patterns[49030] = 29'b1_011111110000_110_1_011111110000;
      patterns[49031] = 29'b1_011111110000_111_1_011111110000;
      patterns[49032] = 29'b1_011111110001_000_1_011111110001;
      patterns[49033] = 29'b1_011111110001_001_1_110001011111;
      patterns[49034] = 29'b1_011111110001_010_0_111111100011;
      patterns[49035] = 29'b1_011111110001_011_1_111111000110;
      patterns[49036] = 29'b1_011111110001_100_1_101111111000;
      patterns[49037] = 29'b1_011111110001_101_0_110111111100;
      patterns[49038] = 29'b1_011111110001_110_1_011111110001;
      patterns[49039] = 29'b1_011111110001_111_1_011111110001;
      patterns[49040] = 29'b1_011111110010_000_1_011111110010;
      patterns[49041] = 29'b1_011111110010_001_1_110010011111;
      patterns[49042] = 29'b1_011111110010_010_0_111111100101;
      patterns[49043] = 29'b1_011111110010_011_1_111111001010;
      patterns[49044] = 29'b1_011111110010_100_0_101111111001;
      patterns[49045] = 29'b1_011111110010_101_1_010111111100;
      patterns[49046] = 29'b1_011111110010_110_1_011111110010;
      patterns[49047] = 29'b1_011111110010_111_1_011111110010;
      patterns[49048] = 29'b1_011111110011_000_1_011111110011;
      patterns[49049] = 29'b1_011111110011_001_1_110011011111;
      patterns[49050] = 29'b1_011111110011_010_0_111111100111;
      patterns[49051] = 29'b1_011111110011_011_1_111111001110;
      patterns[49052] = 29'b1_011111110011_100_1_101111111001;
      patterns[49053] = 29'b1_011111110011_101_1_110111111100;
      patterns[49054] = 29'b1_011111110011_110_1_011111110011;
      patterns[49055] = 29'b1_011111110011_111_1_011111110011;
      patterns[49056] = 29'b1_011111110100_000_1_011111110100;
      patterns[49057] = 29'b1_011111110100_001_1_110100011111;
      patterns[49058] = 29'b1_011111110100_010_0_111111101001;
      patterns[49059] = 29'b1_011111110100_011_1_111111010010;
      patterns[49060] = 29'b1_011111110100_100_0_101111111010;
      patterns[49061] = 29'b1_011111110100_101_0_010111111101;
      patterns[49062] = 29'b1_011111110100_110_1_011111110100;
      patterns[49063] = 29'b1_011111110100_111_1_011111110100;
      patterns[49064] = 29'b1_011111110101_000_1_011111110101;
      patterns[49065] = 29'b1_011111110101_001_1_110101011111;
      patterns[49066] = 29'b1_011111110101_010_0_111111101011;
      patterns[49067] = 29'b1_011111110101_011_1_111111010110;
      patterns[49068] = 29'b1_011111110101_100_1_101111111010;
      patterns[49069] = 29'b1_011111110101_101_0_110111111101;
      patterns[49070] = 29'b1_011111110101_110_1_011111110101;
      patterns[49071] = 29'b1_011111110101_111_1_011111110101;
      patterns[49072] = 29'b1_011111110110_000_1_011111110110;
      patterns[49073] = 29'b1_011111110110_001_1_110110011111;
      patterns[49074] = 29'b1_011111110110_010_0_111111101101;
      patterns[49075] = 29'b1_011111110110_011_1_111111011010;
      patterns[49076] = 29'b1_011111110110_100_0_101111111011;
      patterns[49077] = 29'b1_011111110110_101_1_010111111101;
      patterns[49078] = 29'b1_011111110110_110_1_011111110110;
      patterns[49079] = 29'b1_011111110110_111_1_011111110110;
      patterns[49080] = 29'b1_011111110111_000_1_011111110111;
      patterns[49081] = 29'b1_011111110111_001_1_110111011111;
      patterns[49082] = 29'b1_011111110111_010_0_111111101111;
      patterns[49083] = 29'b1_011111110111_011_1_111111011110;
      patterns[49084] = 29'b1_011111110111_100_1_101111111011;
      patterns[49085] = 29'b1_011111110111_101_1_110111111101;
      patterns[49086] = 29'b1_011111110111_110_1_011111110111;
      patterns[49087] = 29'b1_011111110111_111_1_011111110111;
      patterns[49088] = 29'b1_011111111000_000_1_011111111000;
      patterns[49089] = 29'b1_011111111000_001_1_111000011111;
      patterns[49090] = 29'b1_011111111000_010_0_111111110001;
      patterns[49091] = 29'b1_011111111000_011_1_111111100010;
      patterns[49092] = 29'b1_011111111000_100_0_101111111100;
      patterns[49093] = 29'b1_011111111000_101_0_010111111110;
      patterns[49094] = 29'b1_011111111000_110_1_011111111000;
      patterns[49095] = 29'b1_011111111000_111_1_011111111000;
      patterns[49096] = 29'b1_011111111001_000_1_011111111001;
      patterns[49097] = 29'b1_011111111001_001_1_111001011111;
      patterns[49098] = 29'b1_011111111001_010_0_111111110011;
      patterns[49099] = 29'b1_011111111001_011_1_111111100110;
      patterns[49100] = 29'b1_011111111001_100_1_101111111100;
      patterns[49101] = 29'b1_011111111001_101_0_110111111110;
      patterns[49102] = 29'b1_011111111001_110_1_011111111001;
      patterns[49103] = 29'b1_011111111001_111_1_011111111001;
      patterns[49104] = 29'b1_011111111010_000_1_011111111010;
      patterns[49105] = 29'b1_011111111010_001_1_111010011111;
      patterns[49106] = 29'b1_011111111010_010_0_111111110101;
      patterns[49107] = 29'b1_011111111010_011_1_111111101010;
      patterns[49108] = 29'b1_011111111010_100_0_101111111101;
      patterns[49109] = 29'b1_011111111010_101_1_010111111110;
      patterns[49110] = 29'b1_011111111010_110_1_011111111010;
      patterns[49111] = 29'b1_011111111010_111_1_011111111010;
      patterns[49112] = 29'b1_011111111011_000_1_011111111011;
      patterns[49113] = 29'b1_011111111011_001_1_111011011111;
      patterns[49114] = 29'b1_011111111011_010_0_111111110111;
      patterns[49115] = 29'b1_011111111011_011_1_111111101110;
      patterns[49116] = 29'b1_011111111011_100_1_101111111101;
      patterns[49117] = 29'b1_011111111011_101_1_110111111110;
      patterns[49118] = 29'b1_011111111011_110_1_011111111011;
      patterns[49119] = 29'b1_011111111011_111_1_011111111011;
      patterns[49120] = 29'b1_011111111100_000_1_011111111100;
      patterns[49121] = 29'b1_011111111100_001_1_111100011111;
      patterns[49122] = 29'b1_011111111100_010_0_111111111001;
      patterns[49123] = 29'b1_011111111100_011_1_111111110010;
      patterns[49124] = 29'b1_011111111100_100_0_101111111110;
      patterns[49125] = 29'b1_011111111100_101_0_010111111111;
      patterns[49126] = 29'b1_011111111100_110_1_011111111100;
      patterns[49127] = 29'b1_011111111100_111_1_011111111100;
      patterns[49128] = 29'b1_011111111101_000_1_011111111101;
      patterns[49129] = 29'b1_011111111101_001_1_111101011111;
      patterns[49130] = 29'b1_011111111101_010_0_111111111011;
      patterns[49131] = 29'b1_011111111101_011_1_111111110110;
      patterns[49132] = 29'b1_011111111101_100_1_101111111110;
      patterns[49133] = 29'b1_011111111101_101_0_110111111111;
      patterns[49134] = 29'b1_011111111101_110_1_011111111101;
      patterns[49135] = 29'b1_011111111101_111_1_011111111101;
      patterns[49136] = 29'b1_011111111110_000_1_011111111110;
      patterns[49137] = 29'b1_011111111110_001_1_111110011111;
      patterns[49138] = 29'b1_011111111110_010_0_111111111101;
      patterns[49139] = 29'b1_011111111110_011_1_111111111010;
      patterns[49140] = 29'b1_011111111110_100_0_101111111111;
      patterns[49141] = 29'b1_011111111110_101_1_010111111111;
      patterns[49142] = 29'b1_011111111110_110_1_011111111110;
      patterns[49143] = 29'b1_011111111110_111_1_011111111110;
      patterns[49144] = 29'b1_011111111111_000_1_011111111111;
      patterns[49145] = 29'b1_011111111111_001_1_111111011111;
      patterns[49146] = 29'b1_011111111111_010_0_111111111111;
      patterns[49147] = 29'b1_011111111111_011_1_111111111110;
      patterns[49148] = 29'b1_011111111111_100_1_101111111111;
      patterns[49149] = 29'b1_011111111111_101_1_110111111111;
      patterns[49150] = 29'b1_011111111111_110_1_011111111111;
      patterns[49151] = 29'b1_011111111111_111_1_011111111111;
      patterns[49152] = 29'b1_100000000000_000_1_100000000000;
      patterns[49153] = 29'b1_100000000000_001_1_000000100000;
      patterns[49154] = 29'b1_100000000000_010_1_000000000001;
      patterns[49155] = 29'b1_100000000000_011_0_000000000011;
      patterns[49156] = 29'b1_100000000000_100_0_110000000000;
      patterns[49157] = 29'b1_100000000000_101_0_011000000000;
      patterns[49158] = 29'b1_100000000000_110_1_100000000000;
      patterns[49159] = 29'b1_100000000000_111_1_100000000000;
      patterns[49160] = 29'b1_100000000001_000_1_100000000001;
      patterns[49161] = 29'b1_100000000001_001_1_000001100000;
      patterns[49162] = 29'b1_100000000001_010_1_000000000011;
      patterns[49163] = 29'b1_100000000001_011_0_000000000111;
      patterns[49164] = 29'b1_100000000001_100_1_110000000000;
      patterns[49165] = 29'b1_100000000001_101_0_111000000000;
      patterns[49166] = 29'b1_100000000001_110_1_100000000001;
      patterns[49167] = 29'b1_100000000001_111_1_100000000001;
      patterns[49168] = 29'b1_100000000010_000_1_100000000010;
      patterns[49169] = 29'b1_100000000010_001_1_000010100000;
      patterns[49170] = 29'b1_100000000010_010_1_000000000101;
      patterns[49171] = 29'b1_100000000010_011_0_000000001011;
      patterns[49172] = 29'b1_100000000010_100_0_110000000001;
      patterns[49173] = 29'b1_100000000010_101_1_011000000000;
      patterns[49174] = 29'b1_100000000010_110_1_100000000010;
      patterns[49175] = 29'b1_100000000010_111_1_100000000010;
      patterns[49176] = 29'b1_100000000011_000_1_100000000011;
      patterns[49177] = 29'b1_100000000011_001_1_000011100000;
      patterns[49178] = 29'b1_100000000011_010_1_000000000111;
      patterns[49179] = 29'b1_100000000011_011_0_000000001111;
      patterns[49180] = 29'b1_100000000011_100_1_110000000001;
      patterns[49181] = 29'b1_100000000011_101_1_111000000000;
      patterns[49182] = 29'b1_100000000011_110_1_100000000011;
      patterns[49183] = 29'b1_100000000011_111_1_100000000011;
      patterns[49184] = 29'b1_100000000100_000_1_100000000100;
      patterns[49185] = 29'b1_100000000100_001_1_000100100000;
      patterns[49186] = 29'b1_100000000100_010_1_000000001001;
      patterns[49187] = 29'b1_100000000100_011_0_000000010011;
      patterns[49188] = 29'b1_100000000100_100_0_110000000010;
      patterns[49189] = 29'b1_100000000100_101_0_011000000001;
      patterns[49190] = 29'b1_100000000100_110_1_100000000100;
      patterns[49191] = 29'b1_100000000100_111_1_100000000100;
      patterns[49192] = 29'b1_100000000101_000_1_100000000101;
      patterns[49193] = 29'b1_100000000101_001_1_000101100000;
      patterns[49194] = 29'b1_100000000101_010_1_000000001011;
      patterns[49195] = 29'b1_100000000101_011_0_000000010111;
      patterns[49196] = 29'b1_100000000101_100_1_110000000010;
      patterns[49197] = 29'b1_100000000101_101_0_111000000001;
      patterns[49198] = 29'b1_100000000101_110_1_100000000101;
      patterns[49199] = 29'b1_100000000101_111_1_100000000101;
      patterns[49200] = 29'b1_100000000110_000_1_100000000110;
      patterns[49201] = 29'b1_100000000110_001_1_000110100000;
      patterns[49202] = 29'b1_100000000110_010_1_000000001101;
      patterns[49203] = 29'b1_100000000110_011_0_000000011011;
      patterns[49204] = 29'b1_100000000110_100_0_110000000011;
      patterns[49205] = 29'b1_100000000110_101_1_011000000001;
      patterns[49206] = 29'b1_100000000110_110_1_100000000110;
      patterns[49207] = 29'b1_100000000110_111_1_100000000110;
      patterns[49208] = 29'b1_100000000111_000_1_100000000111;
      patterns[49209] = 29'b1_100000000111_001_1_000111100000;
      patterns[49210] = 29'b1_100000000111_010_1_000000001111;
      patterns[49211] = 29'b1_100000000111_011_0_000000011111;
      patterns[49212] = 29'b1_100000000111_100_1_110000000011;
      patterns[49213] = 29'b1_100000000111_101_1_111000000001;
      patterns[49214] = 29'b1_100000000111_110_1_100000000111;
      patterns[49215] = 29'b1_100000000111_111_1_100000000111;
      patterns[49216] = 29'b1_100000001000_000_1_100000001000;
      patterns[49217] = 29'b1_100000001000_001_1_001000100000;
      patterns[49218] = 29'b1_100000001000_010_1_000000010001;
      patterns[49219] = 29'b1_100000001000_011_0_000000100011;
      patterns[49220] = 29'b1_100000001000_100_0_110000000100;
      patterns[49221] = 29'b1_100000001000_101_0_011000000010;
      patterns[49222] = 29'b1_100000001000_110_1_100000001000;
      patterns[49223] = 29'b1_100000001000_111_1_100000001000;
      patterns[49224] = 29'b1_100000001001_000_1_100000001001;
      patterns[49225] = 29'b1_100000001001_001_1_001001100000;
      patterns[49226] = 29'b1_100000001001_010_1_000000010011;
      patterns[49227] = 29'b1_100000001001_011_0_000000100111;
      patterns[49228] = 29'b1_100000001001_100_1_110000000100;
      patterns[49229] = 29'b1_100000001001_101_0_111000000010;
      patterns[49230] = 29'b1_100000001001_110_1_100000001001;
      patterns[49231] = 29'b1_100000001001_111_1_100000001001;
      patterns[49232] = 29'b1_100000001010_000_1_100000001010;
      patterns[49233] = 29'b1_100000001010_001_1_001010100000;
      patterns[49234] = 29'b1_100000001010_010_1_000000010101;
      patterns[49235] = 29'b1_100000001010_011_0_000000101011;
      patterns[49236] = 29'b1_100000001010_100_0_110000000101;
      patterns[49237] = 29'b1_100000001010_101_1_011000000010;
      patterns[49238] = 29'b1_100000001010_110_1_100000001010;
      patterns[49239] = 29'b1_100000001010_111_1_100000001010;
      patterns[49240] = 29'b1_100000001011_000_1_100000001011;
      patterns[49241] = 29'b1_100000001011_001_1_001011100000;
      patterns[49242] = 29'b1_100000001011_010_1_000000010111;
      patterns[49243] = 29'b1_100000001011_011_0_000000101111;
      patterns[49244] = 29'b1_100000001011_100_1_110000000101;
      patterns[49245] = 29'b1_100000001011_101_1_111000000010;
      patterns[49246] = 29'b1_100000001011_110_1_100000001011;
      patterns[49247] = 29'b1_100000001011_111_1_100000001011;
      patterns[49248] = 29'b1_100000001100_000_1_100000001100;
      patterns[49249] = 29'b1_100000001100_001_1_001100100000;
      patterns[49250] = 29'b1_100000001100_010_1_000000011001;
      patterns[49251] = 29'b1_100000001100_011_0_000000110011;
      patterns[49252] = 29'b1_100000001100_100_0_110000000110;
      patterns[49253] = 29'b1_100000001100_101_0_011000000011;
      patterns[49254] = 29'b1_100000001100_110_1_100000001100;
      patterns[49255] = 29'b1_100000001100_111_1_100000001100;
      patterns[49256] = 29'b1_100000001101_000_1_100000001101;
      patterns[49257] = 29'b1_100000001101_001_1_001101100000;
      patterns[49258] = 29'b1_100000001101_010_1_000000011011;
      patterns[49259] = 29'b1_100000001101_011_0_000000110111;
      patterns[49260] = 29'b1_100000001101_100_1_110000000110;
      patterns[49261] = 29'b1_100000001101_101_0_111000000011;
      patterns[49262] = 29'b1_100000001101_110_1_100000001101;
      patterns[49263] = 29'b1_100000001101_111_1_100000001101;
      patterns[49264] = 29'b1_100000001110_000_1_100000001110;
      patterns[49265] = 29'b1_100000001110_001_1_001110100000;
      patterns[49266] = 29'b1_100000001110_010_1_000000011101;
      patterns[49267] = 29'b1_100000001110_011_0_000000111011;
      patterns[49268] = 29'b1_100000001110_100_0_110000000111;
      patterns[49269] = 29'b1_100000001110_101_1_011000000011;
      patterns[49270] = 29'b1_100000001110_110_1_100000001110;
      patterns[49271] = 29'b1_100000001110_111_1_100000001110;
      patterns[49272] = 29'b1_100000001111_000_1_100000001111;
      patterns[49273] = 29'b1_100000001111_001_1_001111100000;
      patterns[49274] = 29'b1_100000001111_010_1_000000011111;
      patterns[49275] = 29'b1_100000001111_011_0_000000111111;
      patterns[49276] = 29'b1_100000001111_100_1_110000000111;
      patterns[49277] = 29'b1_100000001111_101_1_111000000011;
      patterns[49278] = 29'b1_100000001111_110_1_100000001111;
      patterns[49279] = 29'b1_100000001111_111_1_100000001111;
      patterns[49280] = 29'b1_100000010000_000_1_100000010000;
      patterns[49281] = 29'b1_100000010000_001_1_010000100000;
      patterns[49282] = 29'b1_100000010000_010_1_000000100001;
      patterns[49283] = 29'b1_100000010000_011_0_000001000011;
      patterns[49284] = 29'b1_100000010000_100_0_110000001000;
      patterns[49285] = 29'b1_100000010000_101_0_011000000100;
      patterns[49286] = 29'b1_100000010000_110_1_100000010000;
      patterns[49287] = 29'b1_100000010000_111_1_100000010000;
      patterns[49288] = 29'b1_100000010001_000_1_100000010001;
      patterns[49289] = 29'b1_100000010001_001_1_010001100000;
      patterns[49290] = 29'b1_100000010001_010_1_000000100011;
      patterns[49291] = 29'b1_100000010001_011_0_000001000111;
      patterns[49292] = 29'b1_100000010001_100_1_110000001000;
      patterns[49293] = 29'b1_100000010001_101_0_111000000100;
      patterns[49294] = 29'b1_100000010001_110_1_100000010001;
      patterns[49295] = 29'b1_100000010001_111_1_100000010001;
      patterns[49296] = 29'b1_100000010010_000_1_100000010010;
      patterns[49297] = 29'b1_100000010010_001_1_010010100000;
      patterns[49298] = 29'b1_100000010010_010_1_000000100101;
      patterns[49299] = 29'b1_100000010010_011_0_000001001011;
      patterns[49300] = 29'b1_100000010010_100_0_110000001001;
      patterns[49301] = 29'b1_100000010010_101_1_011000000100;
      patterns[49302] = 29'b1_100000010010_110_1_100000010010;
      patterns[49303] = 29'b1_100000010010_111_1_100000010010;
      patterns[49304] = 29'b1_100000010011_000_1_100000010011;
      patterns[49305] = 29'b1_100000010011_001_1_010011100000;
      patterns[49306] = 29'b1_100000010011_010_1_000000100111;
      patterns[49307] = 29'b1_100000010011_011_0_000001001111;
      patterns[49308] = 29'b1_100000010011_100_1_110000001001;
      patterns[49309] = 29'b1_100000010011_101_1_111000000100;
      patterns[49310] = 29'b1_100000010011_110_1_100000010011;
      patterns[49311] = 29'b1_100000010011_111_1_100000010011;
      patterns[49312] = 29'b1_100000010100_000_1_100000010100;
      patterns[49313] = 29'b1_100000010100_001_1_010100100000;
      patterns[49314] = 29'b1_100000010100_010_1_000000101001;
      patterns[49315] = 29'b1_100000010100_011_0_000001010011;
      patterns[49316] = 29'b1_100000010100_100_0_110000001010;
      patterns[49317] = 29'b1_100000010100_101_0_011000000101;
      patterns[49318] = 29'b1_100000010100_110_1_100000010100;
      patterns[49319] = 29'b1_100000010100_111_1_100000010100;
      patterns[49320] = 29'b1_100000010101_000_1_100000010101;
      patterns[49321] = 29'b1_100000010101_001_1_010101100000;
      patterns[49322] = 29'b1_100000010101_010_1_000000101011;
      patterns[49323] = 29'b1_100000010101_011_0_000001010111;
      patterns[49324] = 29'b1_100000010101_100_1_110000001010;
      patterns[49325] = 29'b1_100000010101_101_0_111000000101;
      patterns[49326] = 29'b1_100000010101_110_1_100000010101;
      patterns[49327] = 29'b1_100000010101_111_1_100000010101;
      patterns[49328] = 29'b1_100000010110_000_1_100000010110;
      patterns[49329] = 29'b1_100000010110_001_1_010110100000;
      patterns[49330] = 29'b1_100000010110_010_1_000000101101;
      patterns[49331] = 29'b1_100000010110_011_0_000001011011;
      patterns[49332] = 29'b1_100000010110_100_0_110000001011;
      patterns[49333] = 29'b1_100000010110_101_1_011000000101;
      patterns[49334] = 29'b1_100000010110_110_1_100000010110;
      patterns[49335] = 29'b1_100000010110_111_1_100000010110;
      patterns[49336] = 29'b1_100000010111_000_1_100000010111;
      patterns[49337] = 29'b1_100000010111_001_1_010111100000;
      patterns[49338] = 29'b1_100000010111_010_1_000000101111;
      patterns[49339] = 29'b1_100000010111_011_0_000001011111;
      patterns[49340] = 29'b1_100000010111_100_1_110000001011;
      patterns[49341] = 29'b1_100000010111_101_1_111000000101;
      patterns[49342] = 29'b1_100000010111_110_1_100000010111;
      patterns[49343] = 29'b1_100000010111_111_1_100000010111;
      patterns[49344] = 29'b1_100000011000_000_1_100000011000;
      patterns[49345] = 29'b1_100000011000_001_1_011000100000;
      patterns[49346] = 29'b1_100000011000_010_1_000000110001;
      patterns[49347] = 29'b1_100000011000_011_0_000001100011;
      patterns[49348] = 29'b1_100000011000_100_0_110000001100;
      patterns[49349] = 29'b1_100000011000_101_0_011000000110;
      patterns[49350] = 29'b1_100000011000_110_1_100000011000;
      patterns[49351] = 29'b1_100000011000_111_1_100000011000;
      patterns[49352] = 29'b1_100000011001_000_1_100000011001;
      patterns[49353] = 29'b1_100000011001_001_1_011001100000;
      patterns[49354] = 29'b1_100000011001_010_1_000000110011;
      patterns[49355] = 29'b1_100000011001_011_0_000001100111;
      patterns[49356] = 29'b1_100000011001_100_1_110000001100;
      patterns[49357] = 29'b1_100000011001_101_0_111000000110;
      patterns[49358] = 29'b1_100000011001_110_1_100000011001;
      patterns[49359] = 29'b1_100000011001_111_1_100000011001;
      patterns[49360] = 29'b1_100000011010_000_1_100000011010;
      patterns[49361] = 29'b1_100000011010_001_1_011010100000;
      patterns[49362] = 29'b1_100000011010_010_1_000000110101;
      patterns[49363] = 29'b1_100000011010_011_0_000001101011;
      patterns[49364] = 29'b1_100000011010_100_0_110000001101;
      patterns[49365] = 29'b1_100000011010_101_1_011000000110;
      patterns[49366] = 29'b1_100000011010_110_1_100000011010;
      patterns[49367] = 29'b1_100000011010_111_1_100000011010;
      patterns[49368] = 29'b1_100000011011_000_1_100000011011;
      patterns[49369] = 29'b1_100000011011_001_1_011011100000;
      patterns[49370] = 29'b1_100000011011_010_1_000000110111;
      patterns[49371] = 29'b1_100000011011_011_0_000001101111;
      patterns[49372] = 29'b1_100000011011_100_1_110000001101;
      patterns[49373] = 29'b1_100000011011_101_1_111000000110;
      patterns[49374] = 29'b1_100000011011_110_1_100000011011;
      patterns[49375] = 29'b1_100000011011_111_1_100000011011;
      patterns[49376] = 29'b1_100000011100_000_1_100000011100;
      patterns[49377] = 29'b1_100000011100_001_1_011100100000;
      patterns[49378] = 29'b1_100000011100_010_1_000000111001;
      patterns[49379] = 29'b1_100000011100_011_0_000001110011;
      patterns[49380] = 29'b1_100000011100_100_0_110000001110;
      patterns[49381] = 29'b1_100000011100_101_0_011000000111;
      patterns[49382] = 29'b1_100000011100_110_1_100000011100;
      patterns[49383] = 29'b1_100000011100_111_1_100000011100;
      patterns[49384] = 29'b1_100000011101_000_1_100000011101;
      patterns[49385] = 29'b1_100000011101_001_1_011101100000;
      patterns[49386] = 29'b1_100000011101_010_1_000000111011;
      patterns[49387] = 29'b1_100000011101_011_0_000001110111;
      patterns[49388] = 29'b1_100000011101_100_1_110000001110;
      patterns[49389] = 29'b1_100000011101_101_0_111000000111;
      patterns[49390] = 29'b1_100000011101_110_1_100000011101;
      patterns[49391] = 29'b1_100000011101_111_1_100000011101;
      patterns[49392] = 29'b1_100000011110_000_1_100000011110;
      patterns[49393] = 29'b1_100000011110_001_1_011110100000;
      patterns[49394] = 29'b1_100000011110_010_1_000000111101;
      patterns[49395] = 29'b1_100000011110_011_0_000001111011;
      patterns[49396] = 29'b1_100000011110_100_0_110000001111;
      patterns[49397] = 29'b1_100000011110_101_1_011000000111;
      patterns[49398] = 29'b1_100000011110_110_1_100000011110;
      patterns[49399] = 29'b1_100000011110_111_1_100000011110;
      patterns[49400] = 29'b1_100000011111_000_1_100000011111;
      patterns[49401] = 29'b1_100000011111_001_1_011111100000;
      patterns[49402] = 29'b1_100000011111_010_1_000000111111;
      patterns[49403] = 29'b1_100000011111_011_0_000001111111;
      patterns[49404] = 29'b1_100000011111_100_1_110000001111;
      patterns[49405] = 29'b1_100000011111_101_1_111000000111;
      patterns[49406] = 29'b1_100000011111_110_1_100000011111;
      patterns[49407] = 29'b1_100000011111_111_1_100000011111;
      patterns[49408] = 29'b1_100000100000_000_1_100000100000;
      patterns[49409] = 29'b1_100000100000_001_1_100000100000;
      patterns[49410] = 29'b1_100000100000_010_1_000001000001;
      patterns[49411] = 29'b1_100000100000_011_0_000010000011;
      patterns[49412] = 29'b1_100000100000_100_0_110000010000;
      patterns[49413] = 29'b1_100000100000_101_0_011000001000;
      patterns[49414] = 29'b1_100000100000_110_1_100000100000;
      patterns[49415] = 29'b1_100000100000_111_1_100000100000;
      patterns[49416] = 29'b1_100000100001_000_1_100000100001;
      patterns[49417] = 29'b1_100000100001_001_1_100001100000;
      patterns[49418] = 29'b1_100000100001_010_1_000001000011;
      patterns[49419] = 29'b1_100000100001_011_0_000010000111;
      patterns[49420] = 29'b1_100000100001_100_1_110000010000;
      patterns[49421] = 29'b1_100000100001_101_0_111000001000;
      patterns[49422] = 29'b1_100000100001_110_1_100000100001;
      patterns[49423] = 29'b1_100000100001_111_1_100000100001;
      patterns[49424] = 29'b1_100000100010_000_1_100000100010;
      patterns[49425] = 29'b1_100000100010_001_1_100010100000;
      patterns[49426] = 29'b1_100000100010_010_1_000001000101;
      patterns[49427] = 29'b1_100000100010_011_0_000010001011;
      patterns[49428] = 29'b1_100000100010_100_0_110000010001;
      patterns[49429] = 29'b1_100000100010_101_1_011000001000;
      patterns[49430] = 29'b1_100000100010_110_1_100000100010;
      patterns[49431] = 29'b1_100000100010_111_1_100000100010;
      patterns[49432] = 29'b1_100000100011_000_1_100000100011;
      patterns[49433] = 29'b1_100000100011_001_1_100011100000;
      patterns[49434] = 29'b1_100000100011_010_1_000001000111;
      patterns[49435] = 29'b1_100000100011_011_0_000010001111;
      patterns[49436] = 29'b1_100000100011_100_1_110000010001;
      patterns[49437] = 29'b1_100000100011_101_1_111000001000;
      patterns[49438] = 29'b1_100000100011_110_1_100000100011;
      patterns[49439] = 29'b1_100000100011_111_1_100000100011;
      patterns[49440] = 29'b1_100000100100_000_1_100000100100;
      patterns[49441] = 29'b1_100000100100_001_1_100100100000;
      patterns[49442] = 29'b1_100000100100_010_1_000001001001;
      patterns[49443] = 29'b1_100000100100_011_0_000010010011;
      patterns[49444] = 29'b1_100000100100_100_0_110000010010;
      patterns[49445] = 29'b1_100000100100_101_0_011000001001;
      patterns[49446] = 29'b1_100000100100_110_1_100000100100;
      patterns[49447] = 29'b1_100000100100_111_1_100000100100;
      patterns[49448] = 29'b1_100000100101_000_1_100000100101;
      patterns[49449] = 29'b1_100000100101_001_1_100101100000;
      patterns[49450] = 29'b1_100000100101_010_1_000001001011;
      patterns[49451] = 29'b1_100000100101_011_0_000010010111;
      patterns[49452] = 29'b1_100000100101_100_1_110000010010;
      patterns[49453] = 29'b1_100000100101_101_0_111000001001;
      patterns[49454] = 29'b1_100000100101_110_1_100000100101;
      patterns[49455] = 29'b1_100000100101_111_1_100000100101;
      patterns[49456] = 29'b1_100000100110_000_1_100000100110;
      patterns[49457] = 29'b1_100000100110_001_1_100110100000;
      patterns[49458] = 29'b1_100000100110_010_1_000001001101;
      patterns[49459] = 29'b1_100000100110_011_0_000010011011;
      patterns[49460] = 29'b1_100000100110_100_0_110000010011;
      patterns[49461] = 29'b1_100000100110_101_1_011000001001;
      patterns[49462] = 29'b1_100000100110_110_1_100000100110;
      patterns[49463] = 29'b1_100000100110_111_1_100000100110;
      patterns[49464] = 29'b1_100000100111_000_1_100000100111;
      patterns[49465] = 29'b1_100000100111_001_1_100111100000;
      patterns[49466] = 29'b1_100000100111_010_1_000001001111;
      patterns[49467] = 29'b1_100000100111_011_0_000010011111;
      patterns[49468] = 29'b1_100000100111_100_1_110000010011;
      patterns[49469] = 29'b1_100000100111_101_1_111000001001;
      patterns[49470] = 29'b1_100000100111_110_1_100000100111;
      patterns[49471] = 29'b1_100000100111_111_1_100000100111;
      patterns[49472] = 29'b1_100000101000_000_1_100000101000;
      patterns[49473] = 29'b1_100000101000_001_1_101000100000;
      patterns[49474] = 29'b1_100000101000_010_1_000001010001;
      patterns[49475] = 29'b1_100000101000_011_0_000010100011;
      patterns[49476] = 29'b1_100000101000_100_0_110000010100;
      patterns[49477] = 29'b1_100000101000_101_0_011000001010;
      patterns[49478] = 29'b1_100000101000_110_1_100000101000;
      patterns[49479] = 29'b1_100000101000_111_1_100000101000;
      patterns[49480] = 29'b1_100000101001_000_1_100000101001;
      patterns[49481] = 29'b1_100000101001_001_1_101001100000;
      patterns[49482] = 29'b1_100000101001_010_1_000001010011;
      patterns[49483] = 29'b1_100000101001_011_0_000010100111;
      patterns[49484] = 29'b1_100000101001_100_1_110000010100;
      patterns[49485] = 29'b1_100000101001_101_0_111000001010;
      patterns[49486] = 29'b1_100000101001_110_1_100000101001;
      patterns[49487] = 29'b1_100000101001_111_1_100000101001;
      patterns[49488] = 29'b1_100000101010_000_1_100000101010;
      patterns[49489] = 29'b1_100000101010_001_1_101010100000;
      patterns[49490] = 29'b1_100000101010_010_1_000001010101;
      patterns[49491] = 29'b1_100000101010_011_0_000010101011;
      patterns[49492] = 29'b1_100000101010_100_0_110000010101;
      patterns[49493] = 29'b1_100000101010_101_1_011000001010;
      patterns[49494] = 29'b1_100000101010_110_1_100000101010;
      patterns[49495] = 29'b1_100000101010_111_1_100000101010;
      patterns[49496] = 29'b1_100000101011_000_1_100000101011;
      patterns[49497] = 29'b1_100000101011_001_1_101011100000;
      patterns[49498] = 29'b1_100000101011_010_1_000001010111;
      patterns[49499] = 29'b1_100000101011_011_0_000010101111;
      patterns[49500] = 29'b1_100000101011_100_1_110000010101;
      patterns[49501] = 29'b1_100000101011_101_1_111000001010;
      patterns[49502] = 29'b1_100000101011_110_1_100000101011;
      patterns[49503] = 29'b1_100000101011_111_1_100000101011;
      patterns[49504] = 29'b1_100000101100_000_1_100000101100;
      patterns[49505] = 29'b1_100000101100_001_1_101100100000;
      patterns[49506] = 29'b1_100000101100_010_1_000001011001;
      patterns[49507] = 29'b1_100000101100_011_0_000010110011;
      patterns[49508] = 29'b1_100000101100_100_0_110000010110;
      patterns[49509] = 29'b1_100000101100_101_0_011000001011;
      patterns[49510] = 29'b1_100000101100_110_1_100000101100;
      patterns[49511] = 29'b1_100000101100_111_1_100000101100;
      patterns[49512] = 29'b1_100000101101_000_1_100000101101;
      patterns[49513] = 29'b1_100000101101_001_1_101101100000;
      patterns[49514] = 29'b1_100000101101_010_1_000001011011;
      patterns[49515] = 29'b1_100000101101_011_0_000010110111;
      patterns[49516] = 29'b1_100000101101_100_1_110000010110;
      patterns[49517] = 29'b1_100000101101_101_0_111000001011;
      patterns[49518] = 29'b1_100000101101_110_1_100000101101;
      patterns[49519] = 29'b1_100000101101_111_1_100000101101;
      patterns[49520] = 29'b1_100000101110_000_1_100000101110;
      patterns[49521] = 29'b1_100000101110_001_1_101110100000;
      patterns[49522] = 29'b1_100000101110_010_1_000001011101;
      patterns[49523] = 29'b1_100000101110_011_0_000010111011;
      patterns[49524] = 29'b1_100000101110_100_0_110000010111;
      patterns[49525] = 29'b1_100000101110_101_1_011000001011;
      patterns[49526] = 29'b1_100000101110_110_1_100000101110;
      patterns[49527] = 29'b1_100000101110_111_1_100000101110;
      patterns[49528] = 29'b1_100000101111_000_1_100000101111;
      patterns[49529] = 29'b1_100000101111_001_1_101111100000;
      patterns[49530] = 29'b1_100000101111_010_1_000001011111;
      patterns[49531] = 29'b1_100000101111_011_0_000010111111;
      patterns[49532] = 29'b1_100000101111_100_1_110000010111;
      patterns[49533] = 29'b1_100000101111_101_1_111000001011;
      patterns[49534] = 29'b1_100000101111_110_1_100000101111;
      patterns[49535] = 29'b1_100000101111_111_1_100000101111;
      patterns[49536] = 29'b1_100000110000_000_1_100000110000;
      patterns[49537] = 29'b1_100000110000_001_1_110000100000;
      patterns[49538] = 29'b1_100000110000_010_1_000001100001;
      patterns[49539] = 29'b1_100000110000_011_0_000011000011;
      patterns[49540] = 29'b1_100000110000_100_0_110000011000;
      patterns[49541] = 29'b1_100000110000_101_0_011000001100;
      patterns[49542] = 29'b1_100000110000_110_1_100000110000;
      patterns[49543] = 29'b1_100000110000_111_1_100000110000;
      patterns[49544] = 29'b1_100000110001_000_1_100000110001;
      patterns[49545] = 29'b1_100000110001_001_1_110001100000;
      patterns[49546] = 29'b1_100000110001_010_1_000001100011;
      patterns[49547] = 29'b1_100000110001_011_0_000011000111;
      patterns[49548] = 29'b1_100000110001_100_1_110000011000;
      patterns[49549] = 29'b1_100000110001_101_0_111000001100;
      patterns[49550] = 29'b1_100000110001_110_1_100000110001;
      patterns[49551] = 29'b1_100000110001_111_1_100000110001;
      patterns[49552] = 29'b1_100000110010_000_1_100000110010;
      patterns[49553] = 29'b1_100000110010_001_1_110010100000;
      patterns[49554] = 29'b1_100000110010_010_1_000001100101;
      patterns[49555] = 29'b1_100000110010_011_0_000011001011;
      patterns[49556] = 29'b1_100000110010_100_0_110000011001;
      patterns[49557] = 29'b1_100000110010_101_1_011000001100;
      patterns[49558] = 29'b1_100000110010_110_1_100000110010;
      patterns[49559] = 29'b1_100000110010_111_1_100000110010;
      patterns[49560] = 29'b1_100000110011_000_1_100000110011;
      patterns[49561] = 29'b1_100000110011_001_1_110011100000;
      patterns[49562] = 29'b1_100000110011_010_1_000001100111;
      patterns[49563] = 29'b1_100000110011_011_0_000011001111;
      patterns[49564] = 29'b1_100000110011_100_1_110000011001;
      patterns[49565] = 29'b1_100000110011_101_1_111000001100;
      patterns[49566] = 29'b1_100000110011_110_1_100000110011;
      patterns[49567] = 29'b1_100000110011_111_1_100000110011;
      patterns[49568] = 29'b1_100000110100_000_1_100000110100;
      patterns[49569] = 29'b1_100000110100_001_1_110100100000;
      patterns[49570] = 29'b1_100000110100_010_1_000001101001;
      patterns[49571] = 29'b1_100000110100_011_0_000011010011;
      patterns[49572] = 29'b1_100000110100_100_0_110000011010;
      patterns[49573] = 29'b1_100000110100_101_0_011000001101;
      patterns[49574] = 29'b1_100000110100_110_1_100000110100;
      patterns[49575] = 29'b1_100000110100_111_1_100000110100;
      patterns[49576] = 29'b1_100000110101_000_1_100000110101;
      patterns[49577] = 29'b1_100000110101_001_1_110101100000;
      patterns[49578] = 29'b1_100000110101_010_1_000001101011;
      patterns[49579] = 29'b1_100000110101_011_0_000011010111;
      patterns[49580] = 29'b1_100000110101_100_1_110000011010;
      patterns[49581] = 29'b1_100000110101_101_0_111000001101;
      patterns[49582] = 29'b1_100000110101_110_1_100000110101;
      patterns[49583] = 29'b1_100000110101_111_1_100000110101;
      patterns[49584] = 29'b1_100000110110_000_1_100000110110;
      patterns[49585] = 29'b1_100000110110_001_1_110110100000;
      patterns[49586] = 29'b1_100000110110_010_1_000001101101;
      patterns[49587] = 29'b1_100000110110_011_0_000011011011;
      patterns[49588] = 29'b1_100000110110_100_0_110000011011;
      patterns[49589] = 29'b1_100000110110_101_1_011000001101;
      patterns[49590] = 29'b1_100000110110_110_1_100000110110;
      patterns[49591] = 29'b1_100000110110_111_1_100000110110;
      patterns[49592] = 29'b1_100000110111_000_1_100000110111;
      patterns[49593] = 29'b1_100000110111_001_1_110111100000;
      patterns[49594] = 29'b1_100000110111_010_1_000001101111;
      patterns[49595] = 29'b1_100000110111_011_0_000011011111;
      patterns[49596] = 29'b1_100000110111_100_1_110000011011;
      patterns[49597] = 29'b1_100000110111_101_1_111000001101;
      patterns[49598] = 29'b1_100000110111_110_1_100000110111;
      patterns[49599] = 29'b1_100000110111_111_1_100000110111;
      patterns[49600] = 29'b1_100000111000_000_1_100000111000;
      patterns[49601] = 29'b1_100000111000_001_1_111000100000;
      patterns[49602] = 29'b1_100000111000_010_1_000001110001;
      patterns[49603] = 29'b1_100000111000_011_0_000011100011;
      patterns[49604] = 29'b1_100000111000_100_0_110000011100;
      patterns[49605] = 29'b1_100000111000_101_0_011000001110;
      patterns[49606] = 29'b1_100000111000_110_1_100000111000;
      patterns[49607] = 29'b1_100000111000_111_1_100000111000;
      patterns[49608] = 29'b1_100000111001_000_1_100000111001;
      patterns[49609] = 29'b1_100000111001_001_1_111001100000;
      patterns[49610] = 29'b1_100000111001_010_1_000001110011;
      patterns[49611] = 29'b1_100000111001_011_0_000011100111;
      patterns[49612] = 29'b1_100000111001_100_1_110000011100;
      patterns[49613] = 29'b1_100000111001_101_0_111000001110;
      patterns[49614] = 29'b1_100000111001_110_1_100000111001;
      patterns[49615] = 29'b1_100000111001_111_1_100000111001;
      patterns[49616] = 29'b1_100000111010_000_1_100000111010;
      patterns[49617] = 29'b1_100000111010_001_1_111010100000;
      patterns[49618] = 29'b1_100000111010_010_1_000001110101;
      patterns[49619] = 29'b1_100000111010_011_0_000011101011;
      patterns[49620] = 29'b1_100000111010_100_0_110000011101;
      patterns[49621] = 29'b1_100000111010_101_1_011000001110;
      patterns[49622] = 29'b1_100000111010_110_1_100000111010;
      patterns[49623] = 29'b1_100000111010_111_1_100000111010;
      patterns[49624] = 29'b1_100000111011_000_1_100000111011;
      patterns[49625] = 29'b1_100000111011_001_1_111011100000;
      patterns[49626] = 29'b1_100000111011_010_1_000001110111;
      patterns[49627] = 29'b1_100000111011_011_0_000011101111;
      patterns[49628] = 29'b1_100000111011_100_1_110000011101;
      patterns[49629] = 29'b1_100000111011_101_1_111000001110;
      patterns[49630] = 29'b1_100000111011_110_1_100000111011;
      patterns[49631] = 29'b1_100000111011_111_1_100000111011;
      patterns[49632] = 29'b1_100000111100_000_1_100000111100;
      patterns[49633] = 29'b1_100000111100_001_1_111100100000;
      patterns[49634] = 29'b1_100000111100_010_1_000001111001;
      patterns[49635] = 29'b1_100000111100_011_0_000011110011;
      patterns[49636] = 29'b1_100000111100_100_0_110000011110;
      patterns[49637] = 29'b1_100000111100_101_0_011000001111;
      patterns[49638] = 29'b1_100000111100_110_1_100000111100;
      patterns[49639] = 29'b1_100000111100_111_1_100000111100;
      patterns[49640] = 29'b1_100000111101_000_1_100000111101;
      patterns[49641] = 29'b1_100000111101_001_1_111101100000;
      patterns[49642] = 29'b1_100000111101_010_1_000001111011;
      patterns[49643] = 29'b1_100000111101_011_0_000011110111;
      patterns[49644] = 29'b1_100000111101_100_1_110000011110;
      patterns[49645] = 29'b1_100000111101_101_0_111000001111;
      patterns[49646] = 29'b1_100000111101_110_1_100000111101;
      patterns[49647] = 29'b1_100000111101_111_1_100000111101;
      patterns[49648] = 29'b1_100000111110_000_1_100000111110;
      patterns[49649] = 29'b1_100000111110_001_1_111110100000;
      patterns[49650] = 29'b1_100000111110_010_1_000001111101;
      patterns[49651] = 29'b1_100000111110_011_0_000011111011;
      patterns[49652] = 29'b1_100000111110_100_0_110000011111;
      patterns[49653] = 29'b1_100000111110_101_1_011000001111;
      patterns[49654] = 29'b1_100000111110_110_1_100000111110;
      patterns[49655] = 29'b1_100000111110_111_1_100000111110;
      patterns[49656] = 29'b1_100000111111_000_1_100000111111;
      patterns[49657] = 29'b1_100000111111_001_1_111111100000;
      patterns[49658] = 29'b1_100000111111_010_1_000001111111;
      patterns[49659] = 29'b1_100000111111_011_0_000011111111;
      patterns[49660] = 29'b1_100000111111_100_1_110000011111;
      patterns[49661] = 29'b1_100000111111_101_1_111000001111;
      patterns[49662] = 29'b1_100000111111_110_1_100000111111;
      patterns[49663] = 29'b1_100000111111_111_1_100000111111;
      patterns[49664] = 29'b1_100001000000_000_1_100001000000;
      patterns[49665] = 29'b1_100001000000_001_1_000000100001;
      patterns[49666] = 29'b1_100001000000_010_1_000010000001;
      patterns[49667] = 29'b1_100001000000_011_0_000100000011;
      patterns[49668] = 29'b1_100001000000_100_0_110000100000;
      patterns[49669] = 29'b1_100001000000_101_0_011000010000;
      patterns[49670] = 29'b1_100001000000_110_1_100001000000;
      patterns[49671] = 29'b1_100001000000_111_1_100001000000;
      patterns[49672] = 29'b1_100001000001_000_1_100001000001;
      patterns[49673] = 29'b1_100001000001_001_1_000001100001;
      patterns[49674] = 29'b1_100001000001_010_1_000010000011;
      patterns[49675] = 29'b1_100001000001_011_0_000100000111;
      patterns[49676] = 29'b1_100001000001_100_1_110000100000;
      patterns[49677] = 29'b1_100001000001_101_0_111000010000;
      patterns[49678] = 29'b1_100001000001_110_1_100001000001;
      patterns[49679] = 29'b1_100001000001_111_1_100001000001;
      patterns[49680] = 29'b1_100001000010_000_1_100001000010;
      patterns[49681] = 29'b1_100001000010_001_1_000010100001;
      patterns[49682] = 29'b1_100001000010_010_1_000010000101;
      patterns[49683] = 29'b1_100001000010_011_0_000100001011;
      patterns[49684] = 29'b1_100001000010_100_0_110000100001;
      patterns[49685] = 29'b1_100001000010_101_1_011000010000;
      patterns[49686] = 29'b1_100001000010_110_1_100001000010;
      patterns[49687] = 29'b1_100001000010_111_1_100001000010;
      patterns[49688] = 29'b1_100001000011_000_1_100001000011;
      patterns[49689] = 29'b1_100001000011_001_1_000011100001;
      patterns[49690] = 29'b1_100001000011_010_1_000010000111;
      patterns[49691] = 29'b1_100001000011_011_0_000100001111;
      patterns[49692] = 29'b1_100001000011_100_1_110000100001;
      patterns[49693] = 29'b1_100001000011_101_1_111000010000;
      patterns[49694] = 29'b1_100001000011_110_1_100001000011;
      patterns[49695] = 29'b1_100001000011_111_1_100001000011;
      patterns[49696] = 29'b1_100001000100_000_1_100001000100;
      patterns[49697] = 29'b1_100001000100_001_1_000100100001;
      patterns[49698] = 29'b1_100001000100_010_1_000010001001;
      patterns[49699] = 29'b1_100001000100_011_0_000100010011;
      patterns[49700] = 29'b1_100001000100_100_0_110000100010;
      patterns[49701] = 29'b1_100001000100_101_0_011000010001;
      patterns[49702] = 29'b1_100001000100_110_1_100001000100;
      patterns[49703] = 29'b1_100001000100_111_1_100001000100;
      patterns[49704] = 29'b1_100001000101_000_1_100001000101;
      patterns[49705] = 29'b1_100001000101_001_1_000101100001;
      patterns[49706] = 29'b1_100001000101_010_1_000010001011;
      patterns[49707] = 29'b1_100001000101_011_0_000100010111;
      patterns[49708] = 29'b1_100001000101_100_1_110000100010;
      patterns[49709] = 29'b1_100001000101_101_0_111000010001;
      patterns[49710] = 29'b1_100001000101_110_1_100001000101;
      patterns[49711] = 29'b1_100001000101_111_1_100001000101;
      patterns[49712] = 29'b1_100001000110_000_1_100001000110;
      patterns[49713] = 29'b1_100001000110_001_1_000110100001;
      patterns[49714] = 29'b1_100001000110_010_1_000010001101;
      patterns[49715] = 29'b1_100001000110_011_0_000100011011;
      patterns[49716] = 29'b1_100001000110_100_0_110000100011;
      patterns[49717] = 29'b1_100001000110_101_1_011000010001;
      patterns[49718] = 29'b1_100001000110_110_1_100001000110;
      patterns[49719] = 29'b1_100001000110_111_1_100001000110;
      patterns[49720] = 29'b1_100001000111_000_1_100001000111;
      patterns[49721] = 29'b1_100001000111_001_1_000111100001;
      patterns[49722] = 29'b1_100001000111_010_1_000010001111;
      patterns[49723] = 29'b1_100001000111_011_0_000100011111;
      patterns[49724] = 29'b1_100001000111_100_1_110000100011;
      patterns[49725] = 29'b1_100001000111_101_1_111000010001;
      patterns[49726] = 29'b1_100001000111_110_1_100001000111;
      patterns[49727] = 29'b1_100001000111_111_1_100001000111;
      patterns[49728] = 29'b1_100001001000_000_1_100001001000;
      patterns[49729] = 29'b1_100001001000_001_1_001000100001;
      patterns[49730] = 29'b1_100001001000_010_1_000010010001;
      patterns[49731] = 29'b1_100001001000_011_0_000100100011;
      patterns[49732] = 29'b1_100001001000_100_0_110000100100;
      patterns[49733] = 29'b1_100001001000_101_0_011000010010;
      patterns[49734] = 29'b1_100001001000_110_1_100001001000;
      patterns[49735] = 29'b1_100001001000_111_1_100001001000;
      patterns[49736] = 29'b1_100001001001_000_1_100001001001;
      patterns[49737] = 29'b1_100001001001_001_1_001001100001;
      patterns[49738] = 29'b1_100001001001_010_1_000010010011;
      patterns[49739] = 29'b1_100001001001_011_0_000100100111;
      patterns[49740] = 29'b1_100001001001_100_1_110000100100;
      patterns[49741] = 29'b1_100001001001_101_0_111000010010;
      patterns[49742] = 29'b1_100001001001_110_1_100001001001;
      patterns[49743] = 29'b1_100001001001_111_1_100001001001;
      patterns[49744] = 29'b1_100001001010_000_1_100001001010;
      patterns[49745] = 29'b1_100001001010_001_1_001010100001;
      patterns[49746] = 29'b1_100001001010_010_1_000010010101;
      patterns[49747] = 29'b1_100001001010_011_0_000100101011;
      patterns[49748] = 29'b1_100001001010_100_0_110000100101;
      patterns[49749] = 29'b1_100001001010_101_1_011000010010;
      patterns[49750] = 29'b1_100001001010_110_1_100001001010;
      patterns[49751] = 29'b1_100001001010_111_1_100001001010;
      patterns[49752] = 29'b1_100001001011_000_1_100001001011;
      patterns[49753] = 29'b1_100001001011_001_1_001011100001;
      patterns[49754] = 29'b1_100001001011_010_1_000010010111;
      patterns[49755] = 29'b1_100001001011_011_0_000100101111;
      patterns[49756] = 29'b1_100001001011_100_1_110000100101;
      patterns[49757] = 29'b1_100001001011_101_1_111000010010;
      patterns[49758] = 29'b1_100001001011_110_1_100001001011;
      patterns[49759] = 29'b1_100001001011_111_1_100001001011;
      patterns[49760] = 29'b1_100001001100_000_1_100001001100;
      patterns[49761] = 29'b1_100001001100_001_1_001100100001;
      patterns[49762] = 29'b1_100001001100_010_1_000010011001;
      patterns[49763] = 29'b1_100001001100_011_0_000100110011;
      patterns[49764] = 29'b1_100001001100_100_0_110000100110;
      patterns[49765] = 29'b1_100001001100_101_0_011000010011;
      patterns[49766] = 29'b1_100001001100_110_1_100001001100;
      patterns[49767] = 29'b1_100001001100_111_1_100001001100;
      patterns[49768] = 29'b1_100001001101_000_1_100001001101;
      patterns[49769] = 29'b1_100001001101_001_1_001101100001;
      patterns[49770] = 29'b1_100001001101_010_1_000010011011;
      patterns[49771] = 29'b1_100001001101_011_0_000100110111;
      patterns[49772] = 29'b1_100001001101_100_1_110000100110;
      patterns[49773] = 29'b1_100001001101_101_0_111000010011;
      patterns[49774] = 29'b1_100001001101_110_1_100001001101;
      patterns[49775] = 29'b1_100001001101_111_1_100001001101;
      patterns[49776] = 29'b1_100001001110_000_1_100001001110;
      patterns[49777] = 29'b1_100001001110_001_1_001110100001;
      patterns[49778] = 29'b1_100001001110_010_1_000010011101;
      patterns[49779] = 29'b1_100001001110_011_0_000100111011;
      patterns[49780] = 29'b1_100001001110_100_0_110000100111;
      patterns[49781] = 29'b1_100001001110_101_1_011000010011;
      patterns[49782] = 29'b1_100001001110_110_1_100001001110;
      patterns[49783] = 29'b1_100001001110_111_1_100001001110;
      patterns[49784] = 29'b1_100001001111_000_1_100001001111;
      patterns[49785] = 29'b1_100001001111_001_1_001111100001;
      patterns[49786] = 29'b1_100001001111_010_1_000010011111;
      patterns[49787] = 29'b1_100001001111_011_0_000100111111;
      patterns[49788] = 29'b1_100001001111_100_1_110000100111;
      patterns[49789] = 29'b1_100001001111_101_1_111000010011;
      patterns[49790] = 29'b1_100001001111_110_1_100001001111;
      patterns[49791] = 29'b1_100001001111_111_1_100001001111;
      patterns[49792] = 29'b1_100001010000_000_1_100001010000;
      patterns[49793] = 29'b1_100001010000_001_1_010000100001;
      patterns[49794] = 29'b1_100001010000_010_1_000010100001;
      patterns[49795] = 29'b1_100001010000_011_0_000101000011;
      patterns[49796] = 29'b1_100001010000_100_0_110000101000;
      patterns[49797] = 29'b1_100001010000_101_0_011000010100;
      patterns[49798] = 29'b1_100001010000_110_1_100001010000;
      patterns[49799] = 29'b1_100001010000_111_1_100001010000;
      patterns[49800] = 29'b1_100001010001_000_1_100001010001;
      patterns[49801] = 29'b1_100001010001_001_1_010001100001;
      patterns[49802] = 29'b1_100001010001_010_1_000010100011;
      patterns[49803] = 29'b1_100001010001_011_0_000101000111;
      patterns[49804] = 29'b1_100001010001_100_1_110000101000;
      patterns[49805] = 29'b1_100001010001_101_0_111000010100;
      patterns[49806] = 29'b1_100001010001_110_1_100001010001;
      patterns[49807] = 29'b1_100001010001_111_1_100001010001;
      patterns[49808] = 29'b1_100001010010_000_1_100001010010;
      patterns[49809] = 29'b1_100001010010_001_1_010010100001;
      patterns[49810] = 29'b1_100001010010_010_1_000010100101;
      patterns[49811] = 29'b1_100001010010_011_0_000101001011;
      patterns[49812] = 29'b1_100001010010_100_0_110000101001;
      patterns[49813] = 29'b1_100001010010_101_1_011000010100;
      patterns[49814] = 29'b1_100001010010_110_1_100001010010;
      patterns[49815] = 29'b1_100001010010_111_1_100001010010;
      patterns[49816] = 29'b1_100001010011_000_1_100001010011;
      patterns[49817] = 29'b1_100001010011_001_1_010011100001;
      patterns[49818] = 29'b1_100001010011_010_1_000010100111;
      patterns[49819] = 29'b1_100001010011_011_0_000101001111;
      patterns[49820] = 29'b1_100001010011_100_1_110000101001;
      patterns[49821] = 29'b1_100001010011_101_1_111000010100;
      patterns[49822] = 29'b1_100001010011_110_1_100001010011;
      patterns[49823] = 29'b1_100001010011_111_1_100001010011;
      patterns[49824] = 29'b1_100001010100_000_1_100001010100;
      patterns[49825] = 29'b1_100001010100_001_1_010100100001;
      patterns[49826] = 29'b1_100001010100_010_1_000010101001;
      patterns[49827] = 29'b1_100001010100_011_0_000101010011;
      patterns[49828] = 29'b1_100001010100_100_0_110000101010;
      patterns[49829] = 29'b1_100001010100_101_0_011000010101;
      patterns[49830] = 29'b1_100001010100_110_1_100001010100;
      patterns[49831] = 29'b1_100001010100_111_1_100001010100;
      patterns[49832] = 29'b1_100001010101_000_1_100001010101;
      patterns[49833] = 29'b1_100001010101_001_1_010101100001;
      patterns[49834] = 29'b1_100001010101_010_1_000010101011;
      patterns[49835] = 29'b1_100001010101_011_0_000101010111;
      patterns[49836] = 29'b1_100001010101_100_1_110000101010;
      patterns[49837] = 29'b1_100001010101_101_0_111000010101;
      patterns[49838] = 29'b1_100001010101_110_1_100001010101;
      patterns[49839] = 29'b1_100001010101_111_1_100001010101;
      patterns[49840] = 29'b1_100001010110_000_1_100001010110;
      patterns[49841] = 29'b1_100001010110_001_1_010110100001;
      patterns[49842] = 29'b1_100001010110_010_1_000010101101;
      patterns[49843] = 29'b1_100001010110_011_0_000101011011;
      patterns[49844] = 29'b1_100001010110_100_0_110000101011;
      patterns[49845] = 29'b1_100001010110_101_1_011000010101;
      patterns[49846] = 29'b1_100001010110_110_1_100001010110;
      patterns[49847] = 29'b1_100001010110_111_1_100001010110;
      patterns[49848] = 29'b1_100001010111_000_1_100001010111;
      patterns[49849] = 29'b1_100001010111_001_1_010111100001;
      patterns[49850] = 29'b1_100001010111_010_1_000010101111;
      patterns[49851] = 29'b1_100001010111_011_0_000101011111;
      patterns[49852] = 29'b1_100001010111_100_1_110000101011;
      patterns[49853] = 29'b1_100001010111_101_1_111000010101;
      patterns[49854] = 29'b1_100001010111_110_1_100001010111;
      patterns[49855] = 29'b1_100001010111_111_1_100001010111;
      patterns[49856] = 29'b1_100001011000_000_1_100001011000;
      patterns[49857] = 29'b1_100001011000_001_1_011000100001;
      patterns[49858] = 29'b1_100001011000_010_1_000010110001;
      patterns[49859] = 29'b1_100001011000_011_0_000101100011;
      patterns[49860] = 29'b1_100001011000_100_0_110000101100;
      patterns[49861] = 29'b1_100001011000_101_0_011000010110;
      patterns[49862] = 29'b1_100001011000_110_1_100001011000;
      patterns[49863] = 29'b1_100001011000_111_1_100001011000;
      patterns[49864] = 29'b1_100001011001_000_1_100001011001;
      patterns[49865] = 29'b1_100001011001_001_1_011001100001;
      patterns[49866] = 29'b1_100001011001_010_1_000010110011;
      patterns[49867] = 29'b1_100001011001_011_0_000101100111;
      patterns[49868] = 29'b1_100001011001_100_1_110000101100;
      patterns[49869] = 29'b1_100001011001_101_0_111000010110;
      patterns[49870] = 29'b1_100001011001_110_1_100001011001;
      patterns[49871] = 29'b1_100001011001_111_1_100001011001;
      patterns[49872] = 29'b1_100001011010_000_1_100001011010;
      patterns[49873] = 29'b1_100001011010_001_1_011010100001;
      patterns[49874] = 29'b1_100001011010_010_1_000010110101;
      patterns[49875] = 29'b1_100001011010_011_0_000101101011;
      patterns[49876] = 29'b1_100001011010_100_0_110000101101;
      patterns[49877] = 29'b1_100001011010_101_1_011000010110;
      patterns[49878] = 29'b1_100001011010_110_1_100001011010;
      patterns[49879] = 29'b1_100001011010_111_1_100001011010;
      patterns[49880] = 29'b1_100001011011_000_1_100001011011;
      patterns[49881] = 29'b1_100001011011_001_1_011011100001;
      patterns[49882] = 29'b1_100001011011_010_1_000010110111;
      patterns[49883] = 29'b1_100001011011_011_0_000101101111;
      patterns[49884] = 29'b1_100001011011_100_1_110000101101;
      patterns[49885] = 29'b1_100001011011_101_1_111000010110;
      patterns[49886] = 29'b1_100001011011_110_1_100001011011;
      patterns[49887] = 29'b1_100001011011_111_1_100001011011;
      patterns[49888] = 29'b1_100001011100_000_1_100001011100;
      patterns[49889] = 29'b1_100001011100_001_1_011100100001;
      patterns[49890] = 29'b1_100001011100_010_1_000010111001;
      patterns[49891] = 29'b1_100001011100_011_0_000101110011;
      patterns[49892] = 29'b1_100001011100_100_0_110000101110;
      patterns[49893] = 29'b1_100001011100_101_0_011000010111;
      patterns[49894] = 29'b1_100001011100_110_1_100001011100;
      patterns[49895] = 29'b1_100001011100_111_1_100001011100;
      patterns[49896] = 29'b1_100001011101_000_1_100001011101;
      patterns[49897] = 29'b1_100001011101_001_1_011101100001;
      patterns[49898] = 29'b1_100001011101_010_1_000010111011;
      patterns[49899] = 29'b1_100001011101_011_0_000101110111;
      patterns[49900] = 29'b1_100001011101_100_1_110000101110;
      patterns[49901] = 29'b1_100001011101_101_0_111000010111;
      patterns[49902] = 29'b1_100001011101_110_1_100001011101;
      patterns[49903] = 29'b1_100001011101_111_1_100001011101;
      patterns[49904] = 29'b1_100001011110_000_1_100001011110;
      patterns[49905] = 29'b1_100001011110_001_1_011110100001;
      patterns[49906] = 29'b1_100001011110_010_1_000010111101;
      patterns[49907] = 29'b1_100001011110_011_0_000101111011;
      patterns[49908] = 29'b1_100001011110_100_0_110000101111;
      patterns[49909] = 29'b1_100001011110_101_1_011000010111;
      patterns[49910] = 29'b1_100001011110_110_1_100001011110;
      patterns[49911] = 29'b1_100001011110_111_1_100001011110;
      patterns[49912] = 29'b1_100001011111_000_1_100001011111;
      patterns[49913] = 29'b1_100001011111_001_1_011111100001;
      patterns[49914] = 29'b1_100001011111_010_1_000010111111;
      patterns[49915] = 29'b1_100001011111_011_0_000101111111;
      patterns[49916] = 29'b1_100001011111_100_1_110000101111;
      patterns[49917] = 29'b1_100001011111_101_1_111000010111;
      patterns[49918] = 29'b1_100001011111_110_1_100001011111;
      patterns[49919] = 29'b1_100001011111_111_1_100001011111;
      patterns[49920] = 29'b1_100001100000_000_1_100001100000;
      patterns[49921] = 29'b1_100001100000_001_1_100000100001;
      patterns[49922] = 29'b1_100001100000_010_1_000011000001;
      patterns[49923] = 29'b1_100001100000_011_0_000110000011;
      patterns[49924] = 29'b1_100001100000_100_0_110000110000;
      patterns[49925] = 29'b1_100001100000_101_0_011000011000;
      patterns[49926] = 29'b1_100001100000_110_1_100001100000;
      patterns[49927] = 29'b1_100001100000_111_1_100001100000;
      patterns[49928] = 29'b1_100001100001_000_1_100001100001;
      patterns[49929] = 29'b1_100001100001_001_1_100001100001;
      patterns[49930] = 29'b1_100001100001_010_1_000011000011;
      patterns[49931] = 29'b1_100001100001_011_0_000110000111;
      patterns[49932] = 29'b1_100001100001_100_1_110000110000;
      patterns[49933] = 29'b1_100001100001_101_0_111000011000;
      patterns[49934] = 29'b1_100001100001_110_1_100001100001;
      patterns[49935] = 29'b1_100001100001_111_1_100001100001;
      patterns[49936] = 29'b1_100001100010_000_1_100001100010;
      patterns[49937] = 29'b1_100001100010_001_1_100010100001;
      patterns[49938] = 29'b1_100001100010_010_1_000011000101;
      patterns[49939] = 29'b1_100001100010_011_0_000110001011;
      patterns[49940] = 29'b1_100001100010_100_0_110000110001;
      patterns[49941] = 29'b1_100001100010_101_1_011000011000;
      patterns[49942] = 29'b1_100001100010_110_1_100001100010;
      patterns[49943] = 29'b1_100001100010_111_1_100001100010;
      patterns[49944] = 29'b1_100001100011_000_1_100001100011;
      patterns[49945] = 29'b1_100001100011_001_1_100011100001;
      patterns[49946] = 29'b1_100001100011_010_1_000011000111;
      patterns[49947] = 29'b1_100001100011_011_0_000110001111;
      patterns[49948] = 29'b1_100001100011_100_1_110000110001;
      patterns[49949] = 29'b1_100001100011_101_1_111000011000;
      patterns[49950] = 29'b1_100001100011_110_1_100001100011;
      patterns[49951] = 29'b1_100001100011_111_1_100001100011;
      patterns[49952] = 29'b1_100001100100_000_1_100001100100;
      patterns[49953] = 29'b1_100001100100_001_1_100100100001;
      patterns[49954] = 29'b1_100001100100_010_1_000011001001;
      patterns[49955] = 29'b1_100001100100_011_0_000110010011;
      patterns[49956] = 29'b1_100001100100_100_0_110000110010;
      patterns[49957] = 29'b1_100001100100_101_0_011000011001;
      patterns[49958] = 29'b1_100001100100_110_1_100001100100;
      patterns[49959] = 29'b1_100001100100_111_1_100001100100;
      patterns[49960] = 29'b1_100001100101_000_1_100001100101;
      patterns[49961] = 29'b1_100001100101_001_1_100101100001;
      patterns[49962] = 29'b1_100001100101_010_1_000011001011;
      patterns[49963] = 29'b1_100001100101_011_0_000110010111;
      patterns[49964] = 29'b1_100001100101_100_1_110000110010;
      patterns[49965] = 29'b1_100001100101_101_0_111000011001;
      patterns[49966] = 29'b1_100001100101_110_1_100001100101;
      patterns[49967] = 29'b1_100001100101_111_1_100001100101;
      patterns[49968] = 29'b1_100001100110_000_1_100001100110;
      patterns[49969] = 29'b1_100001100110_001_1_100110100001;
      patterns[49970] = 29'b1_100001100110_010_1_000011001101;
      patterns[49971] = 29'b1_100001100110_011_0_000110011011;
      patterns[49972] = 29'b1_100001100110_100_0_110000110011;
      patterns[49973] = 29'b1_100001100110_101_1_011000011001;
      patterns[49974] = 29'b1_100001100110_110_1_100001100110;
      patterns[49975] = 29'b1_100001100110_111_1_100001100110;
      patterns[49976] = 29'b1_100001100111_000_1_100001100111;
      patterns[49977] = 29'b1_100001100111_001_1_100111100001;
      patterns[49978] = 29'b1_100001100111_010_1_000011001111;
      patterns[49979] = 29'b1_100001100111_011_0_000110011111;
      patterns[49980] = 29'b1_100001100111_100_1_110000110011;
      patterns[49981] = 29'b1_100001100111_101_1_111000011001;
      patterns[49982] = 29'b1_100001100111_110_1_100001100111;
      patterns[49983] = 29'b1_100001100111_111_1_100001100111;
      patterns[49984] = 29'b1_100001101000_000_1_100001101000;
      patterns[49985] = 29'b1_100001101000_001_1_101000100001;
      patterns[49986] = 29'b1_100001101000_010_1_000011010001;
      patterns[49987] = 29'b1_100001101000_011_0_000110100011;
      patterns[49988] = 29'b1_100001101000_100_0_110000110100;
      patterns[49989] = 29'b1_100001101000_101_0_011000011010;
      patterns[49990] = 29'b1_100001101000_110_1_100001101000;
      patterns[49991] = 29'b1_100001101000_111_1_100001101000;
      patterns[49992] = 29'b1_100001101001_000_1_100001101001;
      patterns[49993] = 29'b1_100001101001_001_1_101001100001;
      patterns[49994] = 29'b1_100001101001_010_1_000011010011;
      patterns[49995] = 29'b1_100001101001_011_0_000110100111;
      patterns[49996] = 29'b1_100001101001_100_1_110000110100;
      patterns[49997] = 29'b1_100001101001_101_0_111000011010;
      patterns[49998] = 29'b1_100001101001_110_1_100001101001;
      patterns[49999] = 29'b1_100001101001_111_1_100001101001;
      patterns[50000] = 29'b1_100001101010_000_1_100001101010;
      patterns[50001] = 29'b1_100001101010_001_1_101010100001;
      patterns[50002] = 29'b1_100001101010_010_1_000011010101;
      patterns[50003] = 29'b1_100001101010_011_0_000110101011;
      patterns[50004] = 29'b1_100001101010_100_0_110000110101;
      patterns[50005] = 29'b1_100001101010_101_1_011000011010;
      patterns[50006] = 29'b1_100001101010_110_1_100001101010;
      patterns[50007] = 29'b1_100001101010_111_1_100001101010;
      patterns[50008] = 29'b1_100001101011_000_1_100001101011;
      patterns[50009] = 29'b1_100001101011_001_1_101011100001;
      patterns[50010] = 29'b1_100001101011_010_1_000011010111;
      patterns[50011] = 29'b1_100001101011_011_0_000110101111;
      patterns[50012] = 29'b1_100001101011_100_1_110000110101;
      patterns[50013] = 29'b1_100001101011_101_1_111000011010;
      patterns[50014] = 29'b1_100001101011_110_1_100001101011;
      patterns[50015] = 29'b1_100001101011_111_1_100001101011;
      patterns[50016] = 29'b1_100001101100_000_1_100001101100;
      patterns[50017] = 29'b1_100001101100_001_1_101100100001;
      patterns[50018] = 29'b1_100001101100_010_1_000011011001;
      patterns[50019] = 29'b1_100001101100_011_0_000110110011;
      patterns[50020] = 29'b1_100001101100_100_0_110000110110;
      patterns[50021] = 29'b1_100001101100_101_0_011000011011;
      patterns[50022] = 29'b1_100001101100_110_1_100001101100;
      patterns[50023] = 29'b1_100001101100_111_1_100001101100;
      patterns[50024] = 29'b1_100001101101_000_1_100001101101;
      patterns[50025] = 29'b1_100001101101_001_1_101101100001;
      patterns[50026] = 29'b1_100001101101_010_1_000011011011;
      patterns[50027] = 29'b1_100001101101_011_0_000110110111;
      patterns[50028] = 29'b1_100001101101_100_1_110000110110;
      patterns[50029] = 29'b1_100001101101_101_0_111000011011;
      patterns[50030] = 29'b1_100001101101_110_1_100001101101;
      patterns[50031] = 29'b1_100001101101_111_1_100001101101;
      patterns[50032] = 29'b1_100001101110_000_1_100001101110;
      patterns[50033] = 29'b1_100001101110_001_1_101110100001;
      patterns[50034] = 29'b1_100001101110_010_1_000011011101;
      patterns[50035] = 29'b1_100001101110_011_0_000110111011;
      patterns[50036] = 29'b1_100001101110_100_0_110000110111;
      patterns[50037] = 29'b1_100001101110_101_1_011000011011;
      patterns[50038] = 29'b1_100001101110_110_1_100001101110;
      patterns[50039] = 29'b1_100001101110_111_1_100001101110;
      patterns[50040] = 29'b1_100001101111_000_1_100001101111;
      patterns[50041] = 29'b1_100001101111_001_1_101111100001;
      patterns[50042] = 29'b1_100001101111_010_1_000011011111;
      patterns[50043] = 29'b1_100001101111_011_0_000110111111;
      patterns[50044] = 29'b1_100001101111_100_1_110000110111;
      patterns[50045] = 29'b1_100001101111_101_1_111000011011;
      patterns[50046] = 29'b1_100001101111_110_1_100001101111;
      patterns[50047] = 29'b1_100001101111_111_1_100001101111;
      patterns[50048] = 29'b1_100001110000_000_1_100001110000;
      patterns[50049] = 29'b1_100001110000_001_1_110000100001;
      patterns[50050] = 29'b1_100001110000_010_1_000011100001;
      patterns[50051] = 29'b1_100001110000_011_0_000111000011;
      patterns[50052] = 29'b1_100001110000_100_0_110000111000;
      patterns[50053] = 29'b1_100001110000_101_0_011000011100;
      patterns[50054] = 29'b1_100001110000_110_1_100001110000;
      patterns[50055] = 29'b1_100001110000_111_1_100001110000;
      patterns[50056] = 29'b1_100001110001_000_1_100001110001;
      patterns[50057] = 29'b1_100001110001_001_1_110001100001;
      patterns[50058] = 29'b1_100001110001_010_1_000011100011;
      patterns[50059] = 29'b1_100001110001_011_0_000111000111;
      patterns[50060] = 29'b1_100001110001_100_1_110000111000;
      patterns[50061] = 29'b1_100001110001_101_0_111000011100;
      patterns[50062] = 29'b1_100001110001_110_1_100001110001;
      patterns[50063] = 29'b1_100001110001_111_1_100001110001;
      patterns[50064] = 29'b1_100001110010_000_1_100001110010;
      patterns[50065] = 29'b1_100001110010_001_1_110010100001;
      patterns[50066] = 29'b1_100001110010_010_1_000011100101;
      patterns[50067] = 29'b1_100001110010_011_0_000111001011;
      patterns[50068] = 29'b1_100001110010_100_0_110000111001;
      patterns[50069] = 29'b1_100001110010_101_1_011000011100;
      patterns[50070] = 29'b1_100001110010_110_1_100001110010;
      patterns[50071] = 29'b1_100001110010_111_1_100001110010;
      patterns[50072] = 29'b1_100001110011_000_1_100001110011;
      patterns[50073] = 29'b1_100001110011_001_1_110011100001;
      patterns[50074] = 29'b1_100001110011_010_1_000011100111;
      patterns[50075] = 29'b1_100001110011_011_0_000111001111;
      patterns[50076] = 29'b1_100001110011_100_1_110000111001;
      patterns[50077] = 29'b1_100001110011_101_1_111000011100;
      patterns[50078] = 29'b1_100001110011_110_1_100001110011;
      patterns[50079] = 29'b1_100001110011_111_1_100001110011;
      patterns[50080] = 29'b1_100001110100_000_1_100001110100;
      patterns[50081] = 29'b1_100001110100_001_1_110100100001;
      patterns[50082] = 29'b1_100001110100_010_1_000011101001;
      patterns[50083] = 29'b1_100001110100_011_0_000111010011;
      patterns[50084] = 29'b1_100001110100_100_0_110000111010;
      patterns[50085] = 29'b1_100001110100_101_0_011000011101;
      patterns[50086] = 29'b1_100001110100_110_1_100001110100;
      patterns[50087] = 29'b1_100001110100_111_1_100001110100;
      patterns[50088] = 29'b1_100001110101_000_1_100001110101;
      patterns[50089] = 29'b1_100001110101_001_1_110101100001;
      patterns[50090] = 29'b1_100001110101_010_1_000011101011;
      patterns[50091] = 29'b1_100001110101_011_0_000111010111;
      patterns[50092] = 29'b1_100001110101_100_1_110000111010;
      patterns[50093] = 29'b1_100001110101_101_0_111000011101;
      patterns[50094] = 29'b1_100001110101_110_1_100001110101;
      patterns[50095] = 29'b1_100001110101_111_1_100001110101;
      patterns[50096] = 29'b1_100001110110_000_1_100001110110;
      patterns[50097] = 29'b1_100001110110_001_1_110110100001;
      patterns[50098] = 29'b1_100001110110_010_1_000011101101;
      patterns[50099] = 29'b1_100001110110_011_0_000111011011;
      patterns[50100] = 29'b1_100001110110_100_0_110000111011;
      patterns[50101] = 29'b1_100001110110_101_1_011000011101;
      patterns[50102] = 29'b1_100001110110_110_1_100001110110;
      patterns[50103] = 29'b1_100001110110_111_1_100001110110;
      patterns[50104] = 29'b1_100001110111_000_1_100001110111;
      patterns[50105] = 29'b1_100001110111_001_1_110111100001;
      patterns[50106] = 29'b1_100001110111_010_1_000011101111;
      patterns[50107] = 29'b1_100001110111_011_0_000111011111;
      patterns[50108] = 29'b1_100001110111_100_1_110000111011;
      patterns[50109] = 29'b1_100001110111_101_1_111000011101;
      patterns[50110] = 29'b1_100001110111_110_1_100001110111;
      patterns[50111] = 29'b1_100001110111_111_1_100001110111;
      patterns[50112] = 29'b1_100001111000_000_1_100001111000;
      patterns[50113] = 29'b1_100001111000_001_1_111000100001;
      patterns[50114] = 29'b1_100001111000_010_1_000011110001;
      patterns[50115] = 29'b1_100001111000_011_0_000111100011;
      patterns[50116] = 29'b1_100001111000_100_0_110000111100;
      patterns[50117] = 29'b1_100001111000_101_0_011000011110;
      patterns[50118] = 29'b1_100001111000_110_1_100001111000;
      patterns[50119] = 29'b1_100001111000_111_1_100001111000;
      patterns[50120] = 29'b1_100001111001_000_1_100001111001;
      patterns[50121] = 29'b1_100001111001_001_1_111001100001;
      patterns[50122] = 29'b1_100001111001_010_1_000011110011;
      patterns[50123] = 29'b1_100001111001_011_0_000111100111;
      patterns[50124] = 29'b1_100001111001_100_1_110000111100;
      patterns[50125] = 29'b1_100001111001_101_0_111000011110;
      patterns[50126] = 29'b1_100001111001_110_1_100001111001;
      patterns[50127] = 29'b1_100001111001_111_1_100001111001;
      patterns[50128] = 29'b1_100001111010_000_1_100001111010;
      patterns[50129] = 29'b1_100001111010_001_1_111010100001;
      patterns[50130] = 29'b1_100001111010_010_1_000011110101;
      patterns[50131] = 29'b1_100001111010_011_0_000111101011;
      patterns[50132] = 29'b1_100001111010_100_0_110000111101;
      patterns[50133] = 29'b1_100001111010_101_1_011000011110;
      patterns[50134] = 29'b1_100001111010_110_1_100001111010;
      patterns[50135] = 29'b1_100001111010_111_1_100001111010;
      patterns[50136] = 29'b1_100001111011_000_1_100001111011;
      patterns[50137] = 29'b1_100001111011_001_1_111011100001;
      patterns[50138] = 29'b1_100001111011_010_1_000011110111;
      patterns[50139] = 29'b1_100001111011_011_0_000111101111;
      patterns[50140] = 29'b1_100001111011_100_1_110000111101;
      patterns[50141] = 29'b1_100001111011_101_1_111000011110;
      patterns[50142] = 29'b1_100001111011_110_1_100001111011;
      patterns[50143] = 29'b1_100001111011_111_1_100001111011;
      patterns[50144] = 29'b1_100001111100_000_1_100001111100;
      patterns[50145] = 29'b1_100001111100_001_1_111100100001;
      patterns[50146] = 29'b1_100001111100_010_1_000011111001;
      patterns[50147] = 29'b1_100001111100_011_0_000111110011;
      patterns[50148] = 29'b1_100001111100_100_0_110000111110;
      patterns[50149] = 29'b1_100001111100_101_0_011000011111;
      patterns[50150] = 29'b1_100001111100_110_1_100001111100;
      patterns[50151] = 29'b1_100001111100_111_1_100001111100;
      patterns[50152] = 29'b1_100001111101_000_1_100001111101;
      patterns[50153] = 29'b1_100001111101_001_1_111101100001;
      patterns[50154] = 29'b1_100001111101_010_1_000011111011;
      patterns[50155] = 29'b1_100001111101_011_0_000111110111;
      patterns[50156] = 29'b1_100001111101_100_1_110000111110;
      patterns[50157] = 29'b1_100001111101_101_0_111000011111;
      patterns[50158] = 29'b1_100001111101_110_1_100001111101;
      patterns[50159] = 29'b1_100001111101_111_1_100001111101;
      patterns[50160] = 29'b1_100001111110_000_1_100001111110;
      patterns[50161] = 29'b1_100001111110_001_1_111110100001;
      patterns[50162] = 29'b1_100001111110_010_1_000011111101;
      patterns[50163] = 29'b1_100001111110_011_0_000111111011;
      patterns[50164] = 29'b1_100001111110_100_0_110000111111;
      patterns[50165] = 29'b1_100001111110_101_1_011000011111;
      patterns[50166] = 29'b1_100001111110_110_1_100001111110;
      patterns[50167] = 29'b1_100001111110_111_1_100001111110;
      patterns[50168] = 29'b1_100001111111_000_1_100001111111;
      patterns[50169] = 29'b1_100001111111_001_1_111111100001;
      patterns[50170] = 29'b1_100001111111_010_1_000011111111;
      patterns[50171] = 29'b1_100001111111_011_0_000111111111;
      patterns[50172] = 29'b1_100001111111_100_1_110000111111;
      patterns[50173] = 29'b1_100001111111_101_1_111000011111;
      patterns[50174] = 29'b1_100001111111_110_1_100001111111;
      patterns[50175] = 29'b1_100001111111_111_1_100001111111;
      patterns[50176] = 29'b1_100010000000_000_1_100010000000;
      patterns[50177] = 29'b1_100010000000_001_1_000000100010;
      patterns[50178] = 29'b1_100010000000_010_1_000100000001;
      patterns[50179] = 29'b1_100010000000_011_0_001000000011;
      patterns[50180] = 29'b1_100010000000_100_0_110001000000;
      patterns[50181] = 29'b1_100010000000_101_0_011000100000;
      patterns[50182] = 29'b1_100010000000_110_1_100010000000;
      patterns[50183] = 29'b1_100010000000_111_1_100010000000;
      patterns[50184] = 29'b1_100010000001_000_1_100010000001;
      patterns[50185] = 29'b1_100010000001_001_1_000001100010;
      patterns[50186] = 29'b1_100010000001_010_1_000100000011;
      patterns[50187] = 29'b1_100010000001_011_0_001000000111;
      patterns[50188] = 29'b1_100010000001_100_1_110001000000;
      patterns[50189] = 29'b1_100010000001_101_0_111000100000;
      patterns[50190] = 29'b1_100010000001_110_1_100010000001;
      patterns[50191] = 29'b1_100010000001_111_1_100010000001;
      patterns[50192] = 29'b1_100010000010_000_1_100010000010;
      patterns[50193] = 29'b1_100010000010_001_1_000010100010;
      patterns[50194] = 29'b1_100010000010_010_1_000100000101;
      patterns[50195] = 29'b1_100010000010_011_0_001000001011;
      patterns[50196] = 29'b1_100010000010_100_0_110001000001;
      patterns[50197] = 29'b1_100010000010_101_1_011000100000;
      patterns[50198] = 29'b1_100010000010_110_1_100010000010;
      patterns[50199] = 29'b1_100010000010_111_1_100010000010;
      patterns[50200] = 29'b1_100010000011_000_1_100010000011;
      patterns[50201] = 29'b1_100010000011_001_1_000011100010;
      patterns[50202] = 29'b1_100010000011_010_1_000100000111;
      patterns[50203] = 29'b1_100010000011_011_0_001000001111;
      patterns[50204] = 29'b1_100010000011_100_1_110001000001;
      patterns[50205] = 29'b1_100010000011_101_1_111000100000;
      patterns[50206] = 29'b1_100010000011_110_1_100010000011;
      patterns[50207] = 29'b1_100010000011_111_1_100010000011;
      patterns[50208] = 29'b1_100010000100_000_1_100010000100;
      patterns[50209] = 29'b1_100010000100_001_1_000100100010;
      patterns[50210] = 29'b1_100010000100_010_1_000100001001;
      patterns[50211] = 29'b1_100010000100_011_0_001000010011;
      patterns[50212] = 29'b1_100010000100_100_0_110001000010;
      patterns[50213] = 29'b1_100010000100_101_0_011000100001;
      patterns[50214] = 29'b1_100010000100_110_1_100010000100;
      patterns[50215] = 29'b1_100010000100_111_1_100010000100;
      patterns[50216] = 29'b1_100010000101_000_1_100010000101;
      patterns[50217] = 29'b1_100010000101_001_1_000101100010;
      patterns[50218] = 29'b1_100010000101_010_1_000100001011;
      patterns[50219] = 29'b1_100010000101_011_0_001000010111;
      patterns[50220] = 29'b1_100010000101_100_1_110001000010;
      patterns[50221] = 29'b1_100010000101_101_0_111000100001;
      patterns[50222] = 29'b1_100010000101_110_1_100010000101;
      patterns[50223] = 29'b1_100010000101_111_1_100010000101;
      patterns[50224] = 29'b1_100010000110_000_1_100010000110;
      patterns[50225] = 29'b1_100010000110_001_1_000110100010;
      patterns[50226] = 29'b1_100010000110_010_1_000100001101;
      patterns[50227] = 29'b1_100010000110_011_0_001000011011;
      patterns[50228] = 29'b1_100010000110_100_0_110001000011;
      patterns[50229] = 29'b1_100010000110_101_1_011000100001;
      patterns[50230] = 29'b1_100010000110_110_1_100010000110;
      patterns[50231] = 29'b1_100010000110_111_1_100010000110;
      patterns[50232] = 29'b1_100010000111_000_1_100010000111;
      patterns[50233] = 29'b1_100010000111_001_1_000111100010;
      patterns[50234] = 29'b1_100010000111_010_1_000100001111;
      patterns[50235] = 29'b1_100010000111_011_0_001000011111;
      patterns[50236] = 29'b1_100010000111_100_1_110001000011;
      patterns[50237] = 29'b1_100010000111_101_1_111000100001;
      patterns[50238] = 29'b1_100010000111_110_1_100010000111;
      patterns[50239] = 29'b1_100010000111_111_1_100010000111;
      patterns[50240] = 29'b1_100010001000_000_1_100010001000;
      patterns[50241] = 29'b1_100010001000_001_1_001000100010;
      patterns[50242] = 29'b1_100010001000_010_1_000100010001;
      patterns[50243] = 29'b1_100010001000_011_0_001000100011;
      patterns[50244] = 29'b1_100010001000_100_0_110001000100;
      patterns[50245] = 29'b1_100010001000_101_0_011000100010;
      patterns[50246] = 29'b1_100010001000_110_1_100010001000;
      patterns[50247] = 29'b1_100010001000_111_1_100010001000;
      patterns[50248] = 29'b1_100010001001_000_1_100010001001;
      patterns[50249] = 29'b1_100010001001_001_1_001001100010;
      patterns[50250] = 29'b1_100010001001_010_1_000100010011;
      patterns[50251] = 29'b1_100010001001_011_0_001000100111;
      patterns[50252] = 29'b1_100010001001_100_1_110001000100;
      patterns[50253] = 29'b1_100010001001_101_0_111000100010;
      patterns[50254] = 29'b1_100010001001_110_1_100010001001;
      patterns[50255] = 29'b1_100010001001_111_1_100010001001;
      patterns[50256] = 29'b1_100010001010_000_1_100010001010;
      patterns[50257] = 29'b1_100010001010_001_1_001010100010;
      patterns[50258] = 29'b1_100010001010_010_1_000100010101;
      patterns[50259] = 29'b1_100010001010_011_0_001000101011;
      patterns[50260] = 29'b1_100010001010_100_0_110001000101;
      patterns[50261] = 29'b1_100010001010_101_1_011000100010;
      patterns[50262] = 29'b1_100010001010_110_1_100010001010;
      patterns[50263] = 29'b1_100010001010_111_1_100010001010;
      patterns[50264] = 29'b1_100010001011_000_1_100010001011;
      patterns[50265] = 29'b1_100010001011_001_1_001011100010;
      patterns[50266] = 29'b1_100010001011_010_1_000100010111;
      patterns[50267] = 29'b1_100010001011_011_0_001000101111;
      patterns[50268] = 29'b1_100010001011_100_1_110001000101;
      patterns[50269] = 29'b1_100010001011_101_1_111000100010;
      patterns[50270] = 29'b1_100010001011_110_1_100010001011;
      patterns[50271] = 29'b1_100010001011_111_1_100010001011;
      patterns[50272] = 29'b1_100010001100_000_1_100010001100;
      patterns[50273] = 29'b1_100010001100_001_1_001100100010;
      patterns[50274] = 29'b1_100010001100_010_1_000100011001;
      patterns[50275] = 29'b1_100010001100_011_0_001000110011;
      patterns[50276] = 29'b1_100010001100_100_0_110001000110;
      patterns[50277] = 29'b1_100010001100_101_0_011000100011;
      patterns[50278] = 29'b1_100010001100_110_1_100010001100;
      patterns[50279] = 29'b1_100010001100_111_1_100010001100;
      patterns[50280] = 29'b1_100010001101_000_1_100010001101;
      patterns[50281] = 29'b1_100010001101_001_1_001101100010;
      patterns[50282] = 29'b1_100010001101_010_1_000100011011;
      patterns[50283] = 29'b1_100010001101_011_0_001000110111;
      patterns[50284] = 29'b1_100010001101_100_1_110001000110;
      patterns[50285] = 29'b1_100010001101_101_0_111000100011;
      patterns[50286] = 29'b1_100010001101_110_1_100010001101;
      patterns[50287] = 29'b1_100010001101_111_1_100010001101;
      patterns[50288] = 29'b1_100010001110_000_1_100010001110;
      patterns[50289] = 29'b1_100010001110_001_1_001110100010;
      patterns[50290] = 29'b1_100010001110_010_1_000100011101;
      patterns[50291] = 29'b1_100010001110_011_0_001000111011;
      patterns[50292] = 29'b1_100010001110_100_0_110001000111;
      patterns[50293] = 29'b1_100010001110_101_1_011000100011;
      patterns[50294] = 29'b1_100010001110_110_1_100010001110;
      patterns[50295] = 29'b1_100010001110_111_1_100010001110;
      patterns[50296] = 29'b1_100010001111_000_1_100010001111;
      patterns[50297] = 29'b1_100010001111_001_1_001111100010;
      patterns[50298] = 29'b1_100010001111_010_1_000100011111;
      patterns[50299] = 29'b1_100010001111_011_0_001000111111;
      patterns[50300] = 29'b1_100010001111_100_1_110001000111;
      patterns[50301] = 29'b1_100010001111_101_1_111000100011;
      patterns[50302] = 29'b1_100010001111_110_1_100010001111;
      patterns[50303] = 29'b1_100010001111_111_1_100010001111;
      patterns[50304] = 29'b1_100010010000_000_1_100010010000;
      patterns[50305] = 29'b1_100010010000_001_1_010000100010;
      patterns[50306] = 29'b1_100010010000_010_1_000100100001;
      patterns[50307] = 29'b1_100010010000_011_0_001001000011;
      patterns[50308] = 29'b1_100010010000_100_0_110001001000;
      patterns[50309] = 29'b1_100010010000_101_0_011000100100;
      patterns[50310] = 29'b1_100010010000_110_1_100010010000;
      patterns[50311] = 29'b1_100010010000_111_1_100010010000;
      patterns[50312] = 29'b1_100010010001_000_1_100010010001;
      patterns[50313] = 29'b1_100010010001_001_1_010001100010;
      patterns[50314] = 29'b1_100010010001_010_1_000100100011;
      patterns[50315] = 29'b1_100010010001_011_0_001001000111;
      patterns[50316] = 29'b1_100010010001_100_1_110001001000;
      patterns[50317] = 29'b1_100010010001_101_0_111000100100;
      patterns[50318] = 29'b1_100010010001_110_1_100010010001;
      patterns[50319] = 29'b1_100010010001_111_1_100010010001;
      patterns[50320] = 29'b1_100010010010_000_1_100010010010;
      patterns[50321] = 29'b1_100010010010_001_1_010010100010;
      patterns[50322] = 29'b1_100010010010_010_1_000100100101;
      patterns[50323] = 29'b1_100010010010_011_0_001001001011;
      patterns[50324] = 29'b1_100010010010_100_0_110001001001;
      patterns[50325] = 29'b1_100010010010_101_1_011000100100;
      patterns[50326] = 29'b1_100010010010_110_1_100010010010;
      patterns[50327] = 29'b1_100010010010_111_1_100010010010;
      patterns[50328] = 29'b1_100010010011_000_1_100010010011;
      patterns[50329] = 29'b1_100010010011_001_1_010011100010;
      patterns[50330] = 29'b1_100010010011_010_1_000100100111;
      patterns[50331] = 29'b1_100010010011_011_0_001001001111;
      patterns[50332] = 29'b1_100010010011_100_1_110001001001;
      patterns[50333] = 29'b1_100010010011_101_1_111000100100;
      patterns[50334] = 29'b1_100010010011_110_1_100010010011;
      patterns[50335] = 29'b1_100010010011_111_1_100010010011;
      patterns[50336] = 29'b1_100010010100_000_1_100010010100;
      patterns[50337] = 29'b1_100010010100_001_1_010100100010;
      patterns[50338] = 29'b1_100010010100_010_1_000100101001;
      patterns[50339] = 29'b1_100010010100_011_0_001001010011;
      patterns[50340] = 29'b1_100010010100_100_0_110001001010;
      patterns[50341] = 29'b1_100010010100_101_0_011000100101;
      patterns[50342] = 29'b1_100010010100_110_1_100010010100;
      patterns[50343] = 29'b1_100010010100_111_1_100010010100;
      patterns[50344] = 29'b1_100010010101_000_1_100010010101;
      patterns[50345] = 29'b1_100010010101_001_1_010101100010;
      patterns[50346] = 29'b1_100010010101_010_1_000100101011;
      patterns[50347] = 29'b1_100010010101_011_0_001001010111;
      patterns[50348] = 29'b1_100010010101_100_1_110001001010;
      patterns[50349] = 29'b1_100010010101_101_0_111000100101;
      patterns[50350] = 29'b1_100010010101_110_1_100010010101;
      patterns[50351] = 29'b1_100010010101_111_1_100010010101;
      patterns[50352] = 29'b1_100010010110_000_1_100010010110;
      patterns[50353] = 29'b1_100010010110_001_1_010110100010;
      patterns[50354] = 29'b1_100010010110_010_1_000100101101;
      patterns[50355] = 29'b1_100010010110_011_0_001001011011;
      patterns[50356] = 29'b1_100010010110_100_0_110001001011;
      patterns[50357] = 29'b1_100010010110_101_1_011000100101;
      patterns[50358] = 29'b1_100010010110_110_1_100010010110;
      patterns[50359] = 29'b1_100010010110_111_1_100010010110;
      patterns[50360] = 29'b1_100010010111_000_1_100010010111;
      patterns[50361] = 29'b1_100010010111_001_1_010111100010;
      patterns[50362] = 29'b1_100010010111_010_1_000100101111;
      patterns[50363] = 29'b1_100010010111_011_0_001001011111;
      patterns[50364] = 29'b1_100010010111_100_1_110001001011;
      patterns[50365] = 29'b1_100010010111_101_1_111000100101;
      patterns[50366] = 29'b1_100010010111_110_1_100010010111;
      patterns[50367] = 29'b1_100010010111_111_1_100010010111;
      patterns[50368] = 29'b1_100010011000_000_1_100010011000;
      patterns[50369] = 29'b1_100010011000_001_1_011000100010;
      patterns[50370] = 29'b1_100010011000_010_1_000100110001;
      patterns[50371] = 29'b1_100010011000_011_0_001001100011;
      patterns[50372] = 29'b1_100010011000_100_0_110001001100;
      patterns[50373] = 29'b1_100010011000_101_0_011000100110;
      patterns[50374] = 29'b1_100010011000_110_1_100010011000;
      patterns[50375] = 29'b1_100010011000_111_1_100010011000;
      patterns[50376] = 29'b1_100010011001_000_1_100010011001;
      patterns[50377] = 29'b1_100010011001_001_1_011001100010;
      patterns[50378] = 29'b1_100010011001_010_1_000100110011;
      patterns[50379] = 29'b1_100010011001_011_0_001001100111;
      patterns[50380] = 29'b1_100010011001_100_1_110001001100;
      patterns[50381] = 29'b1_100010011001_101_0_111000100110;
      patterns[50382] = 29'b1_100010011001_110_1_100010011001;
      patterns[50383] = 29'b1_100010011001_111_1_100010011001;
      patterns[50384] = 29'b1_100010011010_000_1_100010011010;
      patterns[50385] = 29'b1_100010011010_001_1_011010100010;
      patterns[50386] = 29'b1_100010011010_010_1_000100110101;
      patterns[50387] = 29'b1_100010011010_011_0_001001101011;
      patterns[50388] = 29'b1_100010011010_100_0_110001001101;
      patterns[50389] = 29'b1_100010011010_101_1_011000100110;
      patterns[50390] = 29'b1_100010011010_110_1_100010011010;
      patterns[50391] = 29'b1_100010011010_111_1_100010011010;
      patterns[50392] = 29'b1_100010011011_000_1_100010011011;
      patterns[50393] = 29'b1_100010011011_001_1_011011100010;
      patterns[50394] = 29'b1_100010011011_010_1_000100110111;
      patterns[50395] = 29'b1_100010011011_011_0_001001101111;
      patterns[50396] = 29'b1_100010011011_100_1_110001001101;
      patterns[50397] = 29'b1_100010011011_101_1_111000100110;
      patterns[50398] = 29'b1_100010011011_110_1_100010011011;
      patterns[50399] = 29'b1_100010011011_111_1_100010011011;
      patterns[50400] = 29'b1_100010011100_000_1_100010011100;
      patterns[50401] = 29'b1_100010011100_001_1_011100100010;
      patterns[50402] = 29'b1_100010011100_010_1_000100111001;
      patterns[50403] = 29'b1_100010011100_011_0_001001110011;
      patterns[50404] = 29'b1_100010011100_100_0_110001001110;
      patterns[50405] = 29'b1_100010011100_101_0_011000100111;
      patterns[50406] = 29'b1_100010011100_110_1_100010011100;
      patterns[50407] = 29'b1_100010011100_111_1_100010011100;
      patterns[50408] = 29'b1_100010011101_000_1_100010011101;
      patterns[50409] = 29'b1_100010011101_001_1_011101100010;
      patterns[50410] = 29'b1_100010011101_010_1_000100111011;
      patterns[50411] = 29'b1_100010011101_011_0_001001110111;
      patterns[50412] = 29'b1_100010011101_100_1_110001001110;
      patterns[50413] = 29'b1_100010011101_101_0_111000100111;
      patterns[50414] = 29'b1_100010011101_110_1_100010011101;
      patterns[50415] = 29'b1_100010011101_111_1_100010011101;
      patterns[50416] = 29'b1_100010011110_000_1_100010011110;
      patterns[50417] = 29'b1_100010011110_001_1_011110100010;
      patterns[50418] = 29'b1_100010011110_010_1_000100111101;
      patterns[50419] = 29'b1_100010011110_011_0_001001111011;
      patterns[50420] = 29'b1_100010011110_100_0_110001001111;
      patterns[50421] = 29'b1_100010011110_101_1_011000100111;
      patterns[50422] = 29'b1_100010011110_110_1_100010011110;
      patterns[50423] = 29'b1_100010011110_111_1_100010011110;
      patterns[50424] = 29'b1_100010011111_000_1_100010011111;
      patterns[50425] = 29'b1_100010011111_001_1_011111100010;
      patterns[50426] = 29'b1_100010011111_010_1_000100111111;
      patterns[50427] = 29'b1_100010011111_011_0_001001111111;
      patterns[50428] = 29'b1_100010011111_100_1_110001001111;
      patterns[50429] = 29'b1_100010011111_101_1_111000100111;
      patterns[50430] = 29'b1_100010011111_110_1_100010011111;
      patterns[50431] = 29'b1_100010011111_111_1_100010011111;
      patterns[50432] = 29'b1_100010100000_000_1_100010100000;
      patterns[50433] = 29'b1_100010100000_001_1_100000100010;
      patterns[50434] = 29'b1_100010100000_010_1_000101000001;
      patterns[50435] = 29'b1_100010100000_011_0_001010000011;
      patterns[50436] = 29'b1_100010100000_100_0_110001010000;
      patterns[50437] = 29'b1_100010100000_101_0_011000101000;
      patterns[50438] = 29'b1_100010100000_110_1_100010100000;
      patterns[50439] = 29'b1_100010100000_111_1_100010100000;
      patterns[50440] = 29'b1_100010100001_000_1_100010100001;
      patterns[50441] = 29'b1_100010100001_001_1_100001100010;
      patterns[50442] = 29'b1_100010100001_010_1_000101000011;
      patterns[50443] = 29'b1_100010100001_011_0_001010000111;
      patterns[50444] = 29'b1_100010100001_100_1_110001010000;
      patterns[50445] = 29'b1_100010100001_101_0_111000101000;
      patterns[50446] = 29'b1_100010100001_110_1_100010100001;
      patterns[50447] = 29'b1_100010100001_111_1_100010100001;
      patterns[50448] = 29'b1_100010100010_000_1_100010100010;
      patterns[50449] = 29'b1_100010100010_001_1_100010100010;
      patterns[50450] = 29'b1_100010100010_010_1_000101000101;
      patterns[50451] = 29'b1_100010100010_011_0_001010001011;
      patterns[50452] = 29'b1_100010100010_100_0_110001010001;
      patterns[50453] = 29'b1_100010100010_101_1_011000101000;
      patterns[50454] = 29'b1_100010100010_110_1_100010100010;
      patterns[50455] = 29'b1_100010100010_111_1_100010100010;
      patterns[50456] = 29'b1_100010100011_000_1_100010100011;
      patterns[50457] = 29'b1_100010100011_001_1_100011100010;
      patterns[50458] = 29'b1_100010100011_010_1_000101000111;
      patterns[50459] = 29'b1_100010100011_011_0_001010001111;
      patterns[50460] = 29'b1_100010100011_100_1_110001010001;
      patterns[50461] = 29'b1_100010100011_101_1_111000101000;
      patterns[50462] = 29'b1_100010100011_110_1_100010100011;
      patterns[50463] = 29'b1_100010100011_111_1_100010100011;
      patterns[50464] = 29'b1_100010100100_000_1_100010100100;
      patterns[50465] = 29'b1_100010100100_001_1_100100100010;
      patterns[50466] = 29'b1_100010100100_010_1_000101001001;
      patterns[50467] = 29'b1_100010100100_011_0_001010010011;
      patterns[50468] = 29'b1_100010100100_100_0_110001010010;
      patterns[50469] = 29'b1_100010100100_101_0_011000101001;
      patterns[50470] = 29'b1_100010100100_110_1_100010100100;
      patterns[50471] = 29'b1_100010100100_111_1_100010100100;
      patterns[50472] = 29'b1_100010100101_000_1_100010100101;
      patterns[50473] = 29'b1_100010100101_001_1_100101100010;
      patterns[50474] = 29'b1_100010100101_010_1_000101001011;
      patterns[50475] = 29'b1_100010100101_011_0_001010010111;
      patterns[50476] = 29'b1_100010100101_100_1_110001010010;
      patterns[50477] = 29'b1_100010100101_101_0_111000101001;
      patterns[50478] = 29'b1_100010100101_110_1_100010100101;
      patterns[50479] = 29'b1_100010100101_111_1_100010100101;
      patterns[50480] = 29'b1_100010100110_000_1_100010100110;
      patterns[50481] = 29'b1_100010100110_001_1_100110100010;
      patterns[50482] = 29'b1_100010100110_010_1_000101001101;
      patterns[50483] = 29'b1_100010100110_011_0_001010011011;
      patterns[50484] = 29'b1_100010100110_100_0_110001010011;
      patterns[50485] = 29'b1_100010100110_101_1_011000101001;
      patterns[50486] = 29'b1_100010100110_110_1_100010100110;
      patterns[50487] = 29'b1_100010100110_111_1_100010100110;
      patterns[50488] = 29'b1_100010100111_000_1_100010100111;
      patterns[50489] = 29'b1_100010100111_001_1_100111100010;
      patterns[50490] = 29'b1_100010100111_010_1_000101001111;
      patterns[50491] = 29'b1_100010100111_011_0_001010011111;
      patterns[50492] = 29'b1_100010100111_100_1_110001010011;
      patterns[50493] = 29'b1_100010100111_101_1_111000101001;
      patterns[50494] = 29'b1_100010100111_110_1_100010100111;
      patterns[50495] = 29'b1_100010100111_111_1_100010100111;
      patterns[50496] = 29'b1_100010101000_000_1_100010101000;
      patterns[50497] = 29'b1_100010101000_001_1_101000100010;
      patterns[50498] = 29'b1_100010101000_010_1_000101010001;
      patterns[50499] = 29'b1_100010101000_011_0_001010100011;
      patterns[50500] = 29'b1_100010101000_100_0_110001010100;
      patterns[50501] = 29'b1_100010101000_101_0_011000101010;
      patterns[50502] = 29'b1_100010101000_110_1_100010101000;
      patterns[50503] = 29'b1_100010101000_111_1_100010101000;
      patterns[50504] = 29'b1_100010101001_000_1_100010101001;
      patterns[50505] = 29'b1_100010101001_001_1_101001100010;
      patterns[50506] = 29'b1_100010101001_010_1_000101010011;
      patterns[50507] = 29'b1_100010101001_011_0_001010100111;
      patterns[50508] = 29'b1_100010101001_100_1_110001010100;
      patterns[50509] = 29'b1_100010101001_101_0_111000101010;
      patterns[50510] = 29'b1_100010101001_110_1_100010101001;
      patterns[50511] = 29'b1_100010101001_111_1_100010101001;
      patterns[50512] = 29'b1_100010101010_000_1_100010101010;
      patterns[50513] = 29'b1_100010101010_001_1_101010100010;
      patterns[50514] = 29'b1_100010101010_010_1_000101010101;
      patterns[50515] = 29'b1_100010101010_011_0_001010101011;
      patterns[50516] = 29'b1_100010101010_100_0_110001010101;
      patterns[50517] = 29'b1_100010101010_101_1_011000101010;
      patterns[50518] = 29'b1_100010101010_110_1_100010101010;
      patterns[50519] = 29'b1_100010101010_111_1_100010101010;
      patterns[50520] = 29'b1_100010101011_000_1_100010101011;
      patterns[50521] = 29'b1_100010101011_001_1_101011100010;
      patterns[50522] = 29'b1_100010101011_010_1_000101010111;
      patterns[50523] = 29'b1_100010101011_011_0_001010101111;
      patterns[50524] = 29'b1_100010101011_100_1_110001010101;
      patterns[50525] = 29'b1_100010101011_101_1_111000101010;
      patterns[50526] = 29'b1_100010101011_110_1_100010101011;
      patterns[50527] = 29'b1_100010101011_111_1_100010101011;
      patterns[50528] = 29'b1_100010101100_000_1_100010101100;
      patterns[50529] = 29'b1_100010101100_001_1_101100100010;
      patterns[50530] = 29'b1_100010101100_010_1_000101011001;
      patterns[50531] = 29'b1_100010101100_011_0_001010110011;
      patterns[50532] = 29'b1_100010101100_100_0_110001010110;
      patterns[50533] = 29'b1_100010101100_101_0_011000101011;
      patterns[50534] = 29'b1_100010101100_110_1_100010101100;
      patterns[50535] = 29'b1_100010101100_111_1_100010101100;
      patterns[50536] = 29'b1_100010101101_000_1_100010101101;
      patterns[50537] = 29'b1_100010101101_001_1_101101100010;
      patterns[50538] = 29'b1_100010101101_010_1_000101011011;
      patterns[50539] = 29'b1_100010101101_011_0_001010110111;
      patterns[50540] = 29'b1_100010101101_100_1_110001010110;
      patterns[50541] = 29'b1_100010101101_101_0_111000101011;
      patterns[50542] = 29'b1_100010101101_110_1_100010101101;
      patterns[50543] = 29'b1_100010101101_111_1_100010101101;
      patterns[50544] = 29'b1_100010101110_000_1_100010101110;
      patterns[50545] = 29'b1_100010101110_001_1_101110100010;
      patterns[50546] = 29'b1_100010101110_010_1_000101011101;
      patterns[50547] = 29'b1_100010101110_011_0_001010111011;
      patterns[50548] = 29'b1_100010101110_100_0_110001010111;
      patterns[50549] = 29'b1_100010101110_101_1_011000101011;
      patterns[50550] = 29'b1_100010101110_110_1_100010101110;
      patterns[50551] = 29'b1_100010101110_111_1_100010101110;
      patterns[50552] = 29'b1_100010101111_000_1_100010101111;
      patterns[50553] = 29'b1_100010101111_001_1_101111100010;
      patterns[50554] = 29'b1_100010101111_010_1_000101011111;
      patterns[50555] = 29'b1_100010101111_011_0_001010111111;
      patterns[50556] = 29'b1_100010101111_100_1_110001010111;
      patterns[50557] = 29'b1_100010101111_101_1_111000101011;
      patterns[50558] = 29'b1_100010101111_110_1_100010101111;
      patterns[50559] = 29'b1_100010101111_111_1_100010101111;
      patterns[50560] = 29'b1_100010110000_000_1_100010110000;
      patterns[50561] = 29'b1_100010110000_001_1_110000100010;
      patterns[50562] = 29'b1_100010110000_010_1_000101100001;
      patterns[50563] = 29'b1_100010110000_011_0_001011000011;
      patterns[50564] = 29'b1_100010110000_100_0_110001011000;
      patterns[50565] = 29'b1_100010110000_101_0_011000101100;
      patterns[50566] = 29'b1_100010110000_110_1_100010110000;
      patterns[50567] = 29'b1_100010110000_111_1_100010110000;
      patterns[50568] = 29'b1_100010110001_000_1_100010110001;
      patterns[50569] = 29'b1_100010110001_001_1_110001100010;
      patterns[50570] = 29'b1_100010110001_010_1_000101100011;
      patterns[50571] = 29'b1_100010110001_011_0_001011000111;
      patterns[50572] = 29'b1_100010110001_100_1_110001011000;
      patterns[50573] = 29'b1_100010110001_101_0_111000101100;
      patterns[50574] = 29'b1_100010110001_110_1_100010110001;
      patterns[50575] = 29'b1_100010110001_111_1_100010110001;
      patterns[50576] = 29'b1_100010110010_000_1_100010110010;
      patterns[50577] = 29'b1_100010110010_001_1_110010100010;
      patterns[50578] = 29'b1_100010110010_010_1_000101100101;
      patterns[50579] = 29'b1_100010110010_011_0_001011001011;
      patterns[50580] = 29'b1_100010110010_100_0_110001011001;
      patterns[50581] = 29'b1_100010110010_101_1_011000101100;
      patterns[50582] = 29'b1_100010110010_110_1_100010110010;
      patterns[50583] = 29'b1_100010110010_111_1_100010110010;
      patterns[50584] = 29'b1_100010110011_000_1_100010110011;
      patterns[50585] = 29'b1_100010110011_001_1_110011100010;
      patterns[50586] = 29'b1_100010110011_010_1_000101100111;
      patterns[50587] = 29'b1_100010110011_011_0_001011001111;
      patterns[50588] = 29'b1_100010110011_100_1_110001011001;
      patterns[50589] = 29'b1_100010110011_101_1_111000101100;
      patterns[50590] = 29'b1_100010110011_110_1_100010110011;
      patterns[50591] = 29'b1_100010110011_111_1_100010110011;
      patterns[50592] = 29'b1_100010110100_000_1_100010110100;
      patterns[50593] = 29'b1_100010110100_001_1_110100100010;
      patterns[50594] = 29'b1_100010110100_010_1_000101101001;
      patterns[50595] = 29'b1_100010110100_011_0_001011010011;
      patterns[50596] = 29'b1_100010110100_100_0_110001011010;
      patterns[50597] = 29'b1_100010110100_101_0_011000101101;
      patterns[50598] = 29'b1_100010110100_110_1_100010110100;
      patterns[50599] = 29'b1_100010110100_111_1_100010110100;
      patterns[50600] = 29'b1_100010110101_000_1_100010110101;
      patterns[50601] = 29'b1_100010110101_001_1_110101100010;
      patterns[50602] = 29'b1_100010110101_010_1_000101101011;
      patterns[50603] = 29'b1_100010110101_011_0_001011010111;
      patterns[50604] = 29'b1_100010110101_100_1_110001011010;
      patterns[50605] = 29'b1_100010110101_101_0_111000101101;
      patterns[50606] = 29'b1_100010110101_110_1_100010110101;
      patterns[50607] = 29'b1_100010110101_111_1_100010110101;
      patterns[50608] = 29'b1_100010110110_000_1_100010110110;
      patterns[50609] = 29'b1_100010110110_001_1_110110100010;
      patterns[50610] = 29'b1_100010110110_010_1_000101101101;
      patterns[50611] = 29'b1_100010110110_011_0_001011011011;
      patterns[50612] = 29'b1_100010110110_100_0_110001011011;
      patterns[50613] = 29'b1_100010110110_101_1_011000101101;
      patterns[50614] = 29'b1_100010110110_110_1_100010110110;
      patterns[50615] = 29'b1_100010110110_111_1_100010110110;
      patterns[50616] = 29'b1_100010110111_000_1_100010110111;
      patterns[50617] = 29'b1_100010110111_001_1_110111100010;
      patterns[50618] = 29'b1_100010110111_010_1_000101101111;
      patterns[50619] = 29'b1_100010110111_011_0_001011011111;
      patterns[50620] = 29'b1_100010110111_100_1_110001011011;
      patterns[50621] = 29'b1_100010110111_101_1_111000101101;
      patterns[50622] = 29'b1_100010110111_110_1_100010110111;
      patterns[50623] = 29'b1_100010110111_111_1_100010110111;
      patterns[50624] = 29'b1_100010111000_000_1_100010111000;
      patterns[50625] = 29'b1_100010111000_001_1_111000100010;
      patterns[50626] = 29'b1_100010111000_010_1_000101110001;
      patterns[50627] = 29'b1_100010111000_011_0_001011100011;
      patterns[50628] = 29'b1_100010111000_100_0_110001011100;
      patterns[50629] = 29'b1_100010111000_101_0_011000101110;
      patterns[50630] = 29'b1_100010111000_110_1_100010111000;
      patterns[50631] = 29'b1_100010111000_111_1_100010111000;
      patterns[50632] = 29'b1_100010111001_000_1_100010111001;
      patterns[50633] = 29'b1_100010111001_001_1_111001100010;
      patterns[50634] = 29'b1_100010111001_010_1_000101110011;
      patterns[50635] = 29'b1_100010111001_011_0_001011100111;
      patterns[50636] = 29'b1_100010111001_100_1_110001011100;
      patterns[50637] = 29'b1_100010111001_101_0_111000101110;
      patterns[50638] = 29'b1_100010111001_110_1_100010111001;
      patterns[50639] = 29'b1_100010111001_111_1_100010111001;
      patterns[50640] = 29'b1_100010111010_000_1_100010111010;
      patterns[50641] = 29'b1_100010111010_001_1_111010100010;
      patterns[50642] = 29'b1_100010111010_010_1_000101110101;
      patterns[50643] = 29'b1_100010111010_011_0_001011101011;
      patterns[50644] = 29'b1_100010111010_100_0_110001011101;
      patterns[50645] = 29'b1_100010111010_101_1_011000101110;
      patterns[50646] = 29'b1_100010111010_110_1_100010111010;
      patterns[50647] = 29'b1_100010111010_111_1_100010111010;
      patterns[50648] = 29'b1_100010111011_000_1_100010111011;
      patterns[50649] = 29'b1_100010111011_001_1_111011100010;
      patterns[50650] = 29'b1_100010111011_010_1_000101110111;
      patterns[50651] = 29'b1_100010111011_011_0_001011101111;
      patterns[50652] = 29'b1_100010111011_100_1_110001011101;
      patterns[50653] = 29'b1_100010111011_101_1_111000101110;
      patterns[50654] = 29'b1_100010111011_110_1_100010111011;
      patterns[50655] = 29'b1_100010111011_111_1_100010111011;
      patterns[50656] = 29'b1_100010111100_000_1_100010111100;
      patterns[50657] = 29'b1_100010111100_001_1_111100100010;
      patterns[50658] = 29'b1_100010111100_010_1_000101111001;
      patterns[50659] = 29'b1_100010111100_011_0_001011110011;
      patterns[50660] = 29'b1_100010111100_100_0_110001011110;
      patterns[50661] = 29'b1_100010111100_101_0_011000101111;
      patterns[50662] = 29'b1_100010111100_110_1_100010111100;
      patterns[50663] = 29'b1_100010111100_111_1_100010111100;
      patterns[50664] = 29'b1_100010111101_000_1_100010111101;
      patterns[50665] = 29'b1_100010111101_001_1_111101100010;
      patterns[50666] = 29'b1_100010111101_010_1_000101111011;
      patterns[50667] = 29'b1_100010111101_011_0_001011110111;
      patterns[50668] = 29'b1_100010111101_100_1_110001011110;
      patterns[50669] = 29'b1_100010111101_101_0_111000101111;
      patterns[50670] = 29'b1_100010111101_110_1_100010111101;
      patterns[50671] = 29'b1_100010111101_111_1_100010111101;
      patterns[50672] = 29'b1_100010111110_000_1_100010111110;
      patterns[50673] = 29'b1_100010111110_001_1_111110100010;
      patterns[50674] = 29'b1_100010111110_010_1_000101111101;
      patterns[50675] = 29'b1_100010111110_011_0_001011111011;
      patterns[50676] = 29'b1_100010111110_100_0_110001011111;
      patterns[50677] = 29'b1_100010111110_101_1_011000101111;
      patterns[50678] = 29'b1_100010111110_110_1_100010111110;
      patterns[50679] = 29'b1_100010111110_111_1_100010111110;
      patterns[50680] = 29'b1_100010111111_000_1_100010111111;
      patterns[50681] = 29'b1_100010111111_001_1_111111100010;
      patterns[50682] = 29'b1_100010111111_010_1_000101111111;
      patterns[50683] = 29'b1_100010111111_011_0_001011111111;
      patterns[50684] = 29'b1_100010111111_100_1_110001011111;
      patterns[50685] = 29'b1_100010111111_101_1_111000101111;
      patterns[50686] = 29'b1_100010111111_110_1_100010111111;
      patterns[50687] = 29'b1_100010111111_111_1_100010111111;
      patterns[50688] = 29'b1_100011000000_000_1_100011000000;
      patterns[50689] = 29'b1_100011000000_001_1_000000100011;
      patterns[50690] = 29'b1_100011000000_010_1_000110000001;
      patterns[50691] = 29'b1_100011000000_011_0_001100000011;
      patterns[50692] = 29'b1_100011000000_100_0_110001100000;
      patterns[50693] = 29'b1_100011000000_101_0_011000110000;
      patterns[50694] = 29'b1_100011000000_110_1_100011000000;
      patterns[50695] = 29'b1_100011000000_111_1_100011000000;
      patterns[50696] = 29'b1_100011000001_000_1_100011000001;
      patterns[50697] = 29'b1_100011000001_001_1_000001100011;
      patterns[50698] = 29'b1_100011000001_010_1_000110000011;
      patterns[50699] = 29'b1_100011000001_011_0_001100000111;
      patterns[50700] = 29'b1_100011000001_100_1_110001100000;
      patterns[50701] = 29'b1_100011000001_101_0_111000110000;
      patterns[50702] = 29'b1_100011000001_110_1_100011000001;
      patterns[50703] = 29'b1_100011000001_111_1_100011000001;
      patterns[50704] = 29'b1_100011000010_000_1_100011000010;
      patterns[50705] = 29'b1_100011000010_001_1_000010100011;
      patterns[50706] = 29'b1_100011000010_010_1_000110000101;
      patterns[50707] = 29'b1_100011000010_011_0_001100001011;
      patterns[50708] = 29'b1_100011000010_100_0_110001100001;
      patterns[50709] = 29'b1_100011000010_101_1_011000110000;
      patterns[50710] = 29'b1_100011000010_110_1_100011000010;
      patterns[50711] = 29'b1_100011000010_111_1_100011000010;
      patterns[50712] = 29'b1_100011000011_000_1_100011000011;
      patterns[50713] = 29'b1_100011000011_001_1_000011100011;
      patterns[50714] = 29'b1_100011000011_010_1_000110000111;
      patterns[50715] = 29'b1_100011000011_011_0_001100001111;
      patterns[50716] = 29'b1_100011000011_100_1_110001100001;
      patterns[50717] = 29'b1_100011000011_101_1_111000110000;
      patterns[50718] = 29'b1_100011000011_110_1_100011000011;
      patterns[50719] = 29'b1_100011000011_111_1_100011000011;
      patterns[50720] = 29'b1_100011000100_000_1_100011000100;
      patterns[50721] = 29'b1_100011000100_001_1_000100100011;
      patterns[50722] = 29'b1_100011000100_010_1_000110001001;
      patterns[50723] = 29'b1_100011000100_011_0_001100010011;
      patterns[50724] = 29'b1_100011000100_100_0_110001100010;
      patterns[50725] = 29'b1_100011000100_101_0_011000110001;
      patterns[50726] = 29'b1_100011000100_110_1_100011000100;
      patterns[50727] = 29'b1_100011000100_111_1_100011000100;
      patterns[50728] = 29'b1_100011000101_000_1_100011000101;
      patterns[50729] = 29'b1_100011000101_001_1_000101100011;
      patterns[50730] = 29'b1_100011000101_010_1_000110001011;
      patterns[50731] = 29'b1_100011000101_011_0_001100010111;
      patterns[50732] = 29'b1_100011000101_100_1_110001100010;
      patterns[50733] = 29'b1_100011000101_101_0_111000110001;
      patterns[50734] = 29'b1_100011000101_110_1_100011000101;
      patterns[50735] = 29'b1_100011000101_111_1_100011000101;
      patterns[50736] = 29'b1_100011000110_000_1_100011000110;
      patterns[50737] = 29'b1_100011000110_001_1_000110100011;
      patterns[50738] = 29'b1_100011000110_010_1_000110001101;
      patterns[50739] = 29'b1_100011000110_011_0_001100011011;
      patterns[50740] = 29'b1_100011000110_100_0_110001100011;
      patterns[50741] = 29'b1_100011000110_101_1_011000110001;
      patterns[50742] = 29'b1_100011000110_110_1_100011000110;
      patterns[50743] = 29'b1_100011000110_111_1_100011000110;
      patterns[50744] = 29'b1_100011000111_000_1_100011000111;
      patterns[50745] = 29'b1_100011000111_001_1_000111100011;
      patterns[50746] = 29'b1_100011000111_010_1_000110001111;
      patterns[50747] = 29'b1_100011000111_011_0_001100011111;
      patterns[50748] = 29'b1_100011000111_100_1_110001100011;
      patterns[50749] = 29'b1_100011000111_101_1_111000110001;
      patterns[50750] = 29'b1_100011000111_110_1_100011000111;
      patterns[50751] = 29'b1_100011000111_111_1_100011000111;
      patterns[50752] = 29'b1_100011001000_000_1_100011001000;
      patterns[50753] = 29'b1_100011001000_001_1_001000100011;
      patterns[50754] = 29'b1_100011001000_010_1_000110010001;
      patterns[50755] = 29'b1_100011001000_011_0_001100100011;
      patterns[50756] = 29'b1_100011001000_100_0_110001100100;
      patterns[50757] = 29'b1_100011001000_101_0_011000110010;
      patterns[50758] = 29'b1_100011001000_110_1_100011001000;
      patterns[50759] = 29'b1_100011001000_111_1_100011001000;
      patterns[50760] = 29'b1_100011001001_000_1_100011001001;
      patterns[50761] = 29'b1_100011001001_001_1_001001100011;
      patterns[50762] = 29'b1_100011001001_010_1_000110010011;
      patterns[50763] = 29'b1_100011001001_011_0_001100100111;
      patterns[50764] = 29'b1_100011001001_100_1_110001100100;
      patterns[50765] = 29'b1_100011001001_101_0_111000110010;
      patterns[50766] = 29'b1_100011001001_110_1_100011001001;
      patterns[50767] = 29'b1_100011001001_111_1_100011001001;
      patterns[50768] = 29'b1_100011001010_000_1_100011001010;
      patterns[50769] = 29'b1_100011001010_001_1_001010100011;
      patterns[50770] = 29'b1_100011001010_010_1_000110010101;
      patterns[50771] = 29'b1_100011001010_011_0_001100101011;
      patterns[50772] = 29'b1_100011001010_100_0_110001100101;
      patterns[50773] = 29'b1_100011001010_101_1_011000110010;
      patterns[50774] = 29'b1_100011001010_110_1_100011001010;
      patterns[50775] = 29'b1_100011001010_111_1_100011001010;
      patterns[50776] = 29'b1_100011001011_000_1_100011001011;
      patterns[50777] = 29'b1_100011001011_001_1_001011100011;
      patterns[50778] = 29'b1_100011001011_010_1_000110010111;
      patterns[50779] = 29'b1_100011001011_011_0_001100101111;
      patterns[50780] = 29'b1_100011001011_100_1_110001100101;
      patterns[50781] = 29'b1_100011001011_101_1_111000110010;
      patterns[50782] = 29'b1_100011001011_110_1_100011001011;
      patterns[50783] = 29'b1_100011001011_111_1_100011001011;
      patterns[50784] = 29'b1_100011001100_000_1_100011001100;
      patterns[50785] = 29'b1_100011001100_001_1_001100100011;
      patterns[50786] = 29'b1_100011001100_010_1_000110011001;
      patterns[50787] = 29'b1_100011001100_011_0_001100110011;
      patterns[50788] = 29'b1_100011001100_100_0_110001100110;
      patterns[50789] = 29'b1_100011001100_101_0_011000110011;
      patterns[50790] = 29'b1_100011001100_110_1_100011001100;
      patterns[50791] = 29'b1_100011001100_111_1_100011001100;
      patterns[50792] = 29'b1_100011001101_000_1_100011001101;
      patterns[50793] = 29'b1_100011001101_001_1_001101100011;
      patterns[50794] = 29'b1_100011001101_010_1_000110011011;
      patterns[50795] = 29'b1_100011001101_011_0_001100110111;
      patterns[50796] = 29'b1_100011001101_100_1_110001100110;
      patterns[50797] = 29'b1_100011001101_101_0_111000110011;
      patterns[50798] = 29'b1_100011001101_110_1_100011001101;
      patterns[50799] = 29'b1_100011001101_111_1_100011001101;
      patterns[50800] = 29'b1_100011001110_000_1_100011001110;
      patterns[50801] = 29'b1_100011001110_001_1_001110100011;
      patterns[50802] = 29'b1_100011001110_010_1_000110011101;
      patterns[50803] = 29'b1_100011001110_011_0_001100111011;
      patterns[50804] = 29'b1_100011001110_100_0_110001100111;
      patterns[50805] = 29'b1_100011001110_101_1_011000110011;
      patterns[50806] = 29'b1_100011001110_110_1_100011001110;
      patterns[50807] = 29'b1_100011001110_111_1_100011001110;
      patterns[50808] = 29'b1_100011001111_000_1_100011001111;
      patterns[50809] = 29'b1_100011001111_001_1_001111100011;
      patterns[50810] = 29'b1_100011001111_010_1_000110011111;
      patterns[50811] = 29'b1_100011001111_011_0_001100111111;
      patterns[50812] = 29'b1_100011001111_100_1_110001100111;
      patterns[50813] = 29'b1_100011001111_101_1_111000110011;
      patterns[50814] = 29'b1_100011001111_110_1_100011001111;
      patterns[50815] = 29'b1_100011001111_111_1_100011001111;
      patterns[50816] = 29'b1_100011010000_000_1_100011010000;
      patterns[50817] = 29'b1_100011010000_001_1_010000100011;
      patterns[50818] = 29'b1_100011010000_010_1_000110100001;
      patterns[50819] = 29'b1_100011010000_011_0_001101000011;
      patterns[50820] = 29'b1_100011010000_100_0_110001101000;
      patterns[50821] = 29'b1_100011010000_101_0_011000110100;
      patterns[50822] = 29'b1_100011010000_110_1_100011010000;
      patterns[50823] = 29'b1_100011010000_111_1_100011010000;
      patterns[50824] = 29'b1_100011010001_000_1_100011010001;
      patterns[50825] = 29'b1_100011010001_001_1_010001100011;
      patterns[50826] = 29'b1_100011010001_010_1_000110100011;
      patterns[50827] = 29'b1_100011010001_011_0_001101000111;
      patterns[50828] = 29'b1_100011010001_100_1_110001101000;
      patterns[50829] = 29'b1_100011010001_101_0_111000110100;
      patterns[50830] = 29'b1_100011010001_110_1_100011010001;
      patterns[50831] = 29'b1_100011010001_111_1_100011010001;
      patterns[50832] = 29'b1_100011010010_000_1_100011010010;
      patterns[50833] = 29'b1_100011010010_001_1_010010100011;
      patterns[50834] = 29'b1_100011010010_010_1_000110100101;
      patterns[50835] = 29'b1_100011010010_011_0_001101001011;
      patterns[50836] = 29'b1_100011010010_100_0_110001101001;
      patterns[50837] = 29'b1_100011010010_101_1_011000110100;
      patterns[50838] = 29'b1_100011010010_110_1_100011010010;
      patterns[50839] = 29'b1_100011010010_111_1_100011010010;
      patterns[50840] = 29'b1_100011010011_000_1_100011010011;
      patterns[50841] = 29'b1_100011010011_001_1_010011100011;
      patterns[50842] = 29'b1_100011010011_010_1_000110100111;
      patterns[50843] = 29'b1_100011010011_011_0_001101001111;
      patterns[50844] = 29'b1_100011010011_100_1_110001101001;
      patterns[50845] = 29'b1_100011010011_101_1_111000110100;
      patterns[50846] = 29'b1_100011010011_110_1_100011010011;
      patterns[50847] = 29'b1_100011010011_111_1_100011010011;
      patterns[50848] = 29'b1_100011010100_000_1_100011010100;
      patterns[50849] = 29'b1_100011010100_001_1_010100100011;
      patterns[50850] = 29'b1_100011010100_010_1_000110101001;
      patterns[50851] = 29'b1_100011010100_011_0_001101010011;
      patterns[50852] = 29'b1_100011010100_100_0_110001101010;
      patterns[50853] = 29'b1_100011010100_101_0_011000110101;
      patterns[50854] = 29'b1_100011010100_110_1_100011010100;
      patterns[50855] = 29'b1_100011010100_111_1_100011010100;
      patterns[50856] = 29'b1_100011010101_000_1_100011010101;
      patterns[50857] = 29'b1_100011010101_001_1_010101100011;
      patterns[50858] = 29'b1_100011010101_010_1_000110101011;
      patterns[50859] = 29'b1_100011010101_011_0_001101010111;
      patterns[50860] = 29'b1_100011010101_100_1_110001101010;
      patterns[50861] = 29'b1_100011010101_101_0_111000110101;
      patterns[50862] = 29'b1_100011010101_110_1_100011010101;
      patterns[50863] = 29'b1_100011010101_111_1_100011010101;
      patterns[50864] = 29'b1_100011010110_000_1_100011010110;
      patterns[50865] = 29'b1_100011010110_001_1_010110100011;
      patterns[50866] = 29'b1_100011010110_010_1_000110101101;
      patterns[50867] = 29'b1_100011010110_011_0_001101011011;
      patterns[50868] = 29'b1_100011010110_100_0_110001101011;
      patterns[50869] = 29'b1_100011010110_101_1_011000110101;
      patterns[50870] = 29'b1_100011010110_110_1_100011010110;
      patterns[50871] = 29'b1_100011010110_111_1_100011010110;
      patterns[50872] = 29'b1_100011010111_000_1_100011010111;
      patterns[50873] = 29'b1_100011010111_001_1_010111100011;
      patterns[50874] = 29'b1_100011010111_010_1_000110101111;
      patterns[50875] = 29'b1_100011010111_011_0_001101011111;
      patterns[50876] = 29'b1_100011010111_100_1_110001101011;
      patterns[50877] = 29'b1_100011010111_101_1_111000110101;
      patterns[50878] = 29'b1_100011010111_110_1_100011010111;
      patterns[50879] = 29'b1_100011010111_111_1_100011010111;
      patterns[50880] = 29'b1_100011011000_000_1_100011011000;
      patterns[50881] = 29'b1_100011011000_001_1_011000100011;
      patterns[50882] = 29'b1_100011011000_010_1_000110110001;
      patterns[50883] = 29'b1_100011011000_011_0_001101100011;
      patterns[50884] = 29'b1_100011011000_100_0_110001101100;
      patterns[50885] = 29'b1_100011011000_101_0_011000110110;
      patterns[50886] = 29'b1_100011011000_110_1_100011011000;
      patterns[50887] = 29'b1_100011011000_111_1_100011011000;
      patterns[50888] = 29'b1_100011011001_000_1_100011011001;
      patterns[50889] = 29'b1_100011011001_001_1_011001100011;
      patterns[50890] = 29'b1_100011011001_010_1_000110110011;
      patterns[50891] = 29'b1_100011011001_011_0_001101100111;
      patterns[50892] = 29'b1_100011011001_100_1_110001101100;
      patterns[50893] = 29'b1_100011011001_101_0_111000110110;
      patterns[50894] = 29'b1_100011011001_110_1_100011011001;
      patterns[50895] = 29'b1_100011011001_111_1_100011011001;
      patterns[50896] = 29'b1_100011011010_000_1_100011011010;
      patterns[50897] = 29'b1_100011011010_001_1_011010100011;
      patterns[50898] = 29'b1_100011011010_010_1_000110110101;
      patterns[50899] = 29'b1_100011011010_011_0_001101101011;
      patterns[50900] = 29'b1_100011011010_100_0_110001101101;
      patterns[50901] = 29'b1_100011011010_101_1_011000110110;
      patterns[50902] = 29'b1_100011011010_110_1_100011011010;
      patterns[50903] = 29'b1_100011011010_111_1_100011011010;
      patterns[50904] = 29'b1_100011011011_000_1_100011011011;
      patterns[50905] = 29'b1_100011011011_001_1_011011100011;
      patterns[50906] = 29'b1_100011011011_010_1_000110110111;
      patterns[50907] = 29'b1_100011011011_011_0_001101101111;
      patterns[50908] = 29'b1_100011011011_100_1_110001101101;
      patterns[50909] = 29'b1_100011011011_101_1_111000110110;
      patterns[50910] = 29'b1_100011011011_110_1_100011011011;
      patterns[50911] = 29'b1_100011011011_111_1_100011011011;
      patterns[50912] = 29'b1_100011011100_000_1_100011011100;
      patterns[50913] = 29'b1_100011011100_001_1_011100100011;
      patterns[50914] = 29'b1_100011011100_010_1_000110111001;
      patterns[50915] = 29'b1_100011011100_011_0_001101110011;
      patterns[50916] = 29'b1_100011011100_100_0_110001101110;
      patterns[50917] = 29'b1_100011011100_101_0_011000110111;
      patterns[50918] = 29'b1_100011011100_110_1_100011011100;
      patterns[50919] = 29'b1_100011011100_111_1_100011011100;
      patterns[50920] = 29'b1_100011011101_000_1_100011011101;
      patterns[50921] = 29'b1_100011011101_001_1_011101100011;
      patterns[50922] = 29'b1_100011011101_010_1_000110111011;
      patterns[50923] = 29'b1_100011011101_011_0_001101110111;
      patterns[50924] = 29'b1_100011011101_100_1_110001101110;
      patterns[50925] = 29'b1_100011011101_101_0_111000110111;
      patterns[50926] = 29'b1_100011011101_110_1_100011011101;
      patterns[50927] = 29'b1_100011011101_111_1_100011011101;
      patterns[50928] = 29'b1_100011011110_000_1_100011011110;
      patterns[50929] = 29'b1_100011011110_001_1_011110100011;
      patterns[50930] = 29'b1_100011011110_010_1_000110111101;
      patterns[50931] = 29'b1_100011011110_011_0_001101111011;
      patterns[50932] = 29'b1_100011011110_100_0_110001101111;
      patterns[50933] = 29'b1_100011011110_101_1_011000110111;
      patterns[50934] = 29'b1_100011011110_110_1_100011011110;
      patterns[50935] = 29'b1_100011011110_111_1_100011011110;
      patterns[50936] = 29'b1_100011011111_000_1_100011011111;
      patterns[50937] = 29'b1_100011011111_001_1_011111100011;
      patterns[50938] = 29'b1_100011011111_010_1_000110111111;
      patterns[50939] = 29'b1_100011011111_011_0_001101111111;
      patterns[50940] = 29'b1_100011011111_100_1_110001101111;
      patterns[50941] = 29'b1_100011011111_101_1_111000110111;
      patterns[50942] = 29'b1_100011011111_110_1_100011011111;
      patterns[50943] = 29'b1_100011011111_111_1_100011011111;
      patterns[50944] = 29'b1_100011100000_000_1_100011100000;
      patterns[50945] = 29'b1_100011100000_001_1_100000100011;
      patterns[50946] = 29'b1_100011100000_010_1_000111000001;
      patterns[50947] = 29'b1_100011100000_011_0_001110000011;
      patterns[50948] = 29'b1_100011100000_100_0_110001110000;
      patterns[50949] = 29'b1_100011100000_101_0_011000111000;
      patterns[50950] = 29'b1_100011100000_110_1_100011100000;
      patterns[50951] = 29'b1_100011100000_111_1_100011100000;
      patterns[50952] = 29'b1_100011100001_000_1_100011100001;
      patterns[50953] = 29'b1_100011100001_001_1_100001100011;
      patterns[50954] = 29'b1_100011100001_010_1_000111000011;
      patterns[50955] = 29'b1_100011100001_011_0_001110000111;
      patterns[50956] = 29'b1_100011100001_100_1_110001110000;
      patterns[50957] = 29'b1_100011100001_101_0_111000111000;
      patterns[50958] = 29'b1_100011100001_110_1_100011100001;
      patterns[50959] = 29'b1_100011100001_111_1_100011100001;
      patterns[50960] = 29'b1_100011100010_000_1_100011100010;
      patterns[50961] = 29'b1_100011100010_001_1_100010100011;
      patterns[50962] = 29'b1_100011100010_010_1_000111000101;
      patterns[50963] = 29'b1_100011100010_011_0_001110001011;
      patterns[50964] = 29'b1_100011100010_100_0_110001110001;
      patterns[50965] = 29'b1_100011100010_101_1_011000111000;
      patterns[50966] = 29'b1_100011100010_110_1_100011100010;
      patterns[50967] = 29'b1_100011100010_111_1_100011100010;
      patterns[50968] = 29'b1_100011100011_000_1_100011100011;
      patterns[50969] = 29'b1_100011100011_001_1_100011100011;
      patterns[50970] = 29'b1_100011100011_010_1_000111000111;
      patterns[50971] = 29'b1_100011100011_011_0_001110001111;
      patterns[50972] = 29'b1_100011100011_100_1_110001110001;
      patterns[50973] = 29'b1_100011100011_101_1_111000111000;
      patterns[50974] = 29'b1_100011100011_110_1_100011100011;
      patterns[50975] = 29'b1_100011100011_111_1_100011100011;
      patterns[50976] = 29'b1_100011100100_000_1_100011100100;
      patterns[50977] = 29'b1_100011100100_001_1_100100100011;
      patterns[50978] = 29'b1_100011100100_010_1_000111001001;
      patterns[50979] = 29'b1_100011100100_011_0_001110010011;
      patterns[50980] = 29'b1_100011100100_100_0_110001110010;
      patterns[50981] = 29'b1_100011100100_101_0_011000111001;
      patterns[50982] = 29'b1_100011100100_110_1_100011100100;
      patterns[50983] = 29'b1_100011100100_111_1_100011100100;
      patterns[50984] = 29'b1_100011100101_000_1_100011100101;
      patterns[50985] = 29'b1_100011100101_001_1_100101100011;
      patterns[50986] = 29'b1_100011100101_010_1_000111001011;
      patterns[50987] = 29'b1_100011100101_011_0_001110010111;
      patterns[50988] = 29'b1_100011100101_100_1_110001110010;
      patterns[50989] = 29'b1_100011100101_101_0_111000111001;
      patterns[50990] = 29'b1_100011100101_110_1_100011100101;
      patterns[50991] = 29'b1_100011100101_111_1_100011100101;
      patterns[50992] = 29'b1_100011100110_000_1_100011100110;
      patterns[50993] = 29'b1_100011100110_001_1_100110100011;
      patterns[50994] = 29'b1_100011100110_010_1_000111001101;
      patterns[50995] = 29'b1_100011100110_011_0_001110011011;
      patterns[50996] = 29'b1_100011100110_100_0_110001110011;
      patterns[50997] = 29'b1_100011100110_101_1_011000111001;
      patterns[50998] = 29'b1_100011100110_110_1_100011100110;
      patterns[50999] = 29'b1_100011100110_111_1_100011100110;
      patterns[51000] = 29'b1_100011100111_000_1_100011100111;
      patterns[51001] = 29'b1_100011100111_001_1_100111100011;
      patterns[51002] = 29'b1_100011100111_010_1_000111001111;
      patterns[51003] = 29'b1_100011100111_011_0_001110011111;
      patterns[51004] = 29'b1_100011100111_100_1_110001110011;
      patterns[51005] = 29'b1_100011100111_101_1_111000111001;
      patterns[51006] = 29'b1_100011100111_110_1_100011100111;
      patterns[51007] = 29'b1_100011100111_111_1_100011100111;
      patterns[51008] = 29'b1_100011101000_000_1_100011101000;
      patterns[51009] = 29'b1_100011101000_001_1_101000100011;
      patterns[51010] = 29'b1_100011101000_010_1_000111010001;
      patterns[51011] = 29'b1_100011101000_011_0_001110100011;
      patterns[51012] = 29'b1_100011101000_100_0_110001110100;
      patterns[51013] = 29'b1_100011101000_101_0_011000111010;
      patterns[51014] = 29'b1_100011101000_110_1_100011101000;
      patterns[51015] = 29'b1_100011101000_111_1_100011101000;
      patterns[51016] = 29'b1_100011101001_000_1_100011101001;
      patterns[51017] = 29'b1_100011101001_001_1_101001100011;
      patterns[51018] = 29'b1_100011101001_010_1_000111010011;
      patterns[51019] = 29'b1_100011101001_011_0_001110100111;
      patterns[51020] = 29'b1_100011101001_100_1_110001110100;
      patterns[51021] = 29'b1_100011101001_101_0_111000111010;
      patterns[51022] = 29'b1_100011101001_110_1_100011101001;
      patterns[51023] = 29'b1_100011101001_111_1_100011101001;
      patterns[51024] = 29'b1_100011101010_000_1_100011101010;
      patterns[51025] = 29'b1_100011101010_001_1_101010100011;
      patterns[51026] = 29'b1_100011101010_010_1_000111010101;
      patterns[51027] = 29'b1_100011101010_011_0_001110101011;
      patterns[51028] = 29'b1_100011101010_100_0_110001110101;
      patterns[51029] = 29'b1_100011101010_101_1_011000111010;
      patterns[51030] = 29'b1_100011101010_110_1_100011101010;
      patterns[51031] = 29'b1_100011101010_111_1_100011101010;
      patterns[51032] = 29'b1_100011101011_000_1_100011101011;
      patterns[51033] = 29'b1_100011101011_001_1_101011100011;
      patterns[51034] = 29'b1_100011101011_010_1_000111010111;
      patterns[51035] = 29'b1_100011101011_011_0_001110101111;
      patterns[51036] = 29'b1_100011101011_100_1_110001110101;
      patterns[51037] = 29'b1_100011101011_101_1_111000111010;
      patterns[51038] = 29'b1_100011101011_110_1_100011101011;
      patterns[51039] = 29'b1_100011101011_111_1_100011101011;
      patterns[51040] = 29'b1_100011101100_000_1_100011101100;
      patterns[51041] = 29'b1_100011101100_001_1_101100100011;
      patterns[51042] = 29'b1_100011101100_010_1_000111011001;
      patterns[51043] = 29'b1_100011101100_011_0_001110110011;
      patterns[51044] = 29'b1_100011101100_100_0_110001110110;
      patterns[51045] = 29'b1_100011101100_101_0_011000111011;
      patterns[51046] = 29'b1_100011101100_110_1_100011101100;
      patterns[51047] = 29'b1_100011101100_111_1_100011101100;
      patterns[51048] = 29'b1_100011101101_000_1_100011101101;
      patterns[51049] = 29'b1_100011101101_001_1_101101100011;
      patterns[51050] = 29'b1_100011101101_010_1_000111011011;
      patterns[51051] = 29'b1_100011101101_011_0_001110110111;
      patterns[51052] = 29'b1_100011101101_100_1_110001110110;
      patterns[51053] = 29'b1_100011101101_101_0_111000111011;
      patterns[51054] = 29'b1_100011101101_110_1_100011101101;
      patterns[51055] = 29'b1_100011101101_111_1_100011101101;
      patterns[51056] = 29'b1_100011101110_000_1_100011101110;
      patterns[51057] = 29'b1_100011101110_001_1_101110100011;
      patterns[51058] = 29'b1_100011101110_010_1_000111011101;
      patterns[51059] = 29'b1_100011101110_011_0_001110111011;
      patterns[51060] = 29'b1_100011101110_100_0_110001110111;
      patterns[51061] = 29'b1_100011101110_101_1_011000111011;
      patterns[51062] = 29'b1_100011101110_110_1_100011101110;
      patterns[51063] = 29'b1_100011101110_111_1_100011101110;
      patterns[51064] = 29'b1_100011101111_000_1_100011101111;
      patterns[51065] = 29'b1_100011101111_001_1_101111100011;
      patterns[51066] = 29'b1_100011101111_010_1_000111011111;
      patterns[51067] = 29'b1_100011101111_011_0_001110111111;
      patterns[51068] = 29'b1_100011101111_100_1_110001110111;
      patterns[51069] = 29'b1_100011101111_101_1_111000111011;
      patterns[51070] = 29'b1_100011101111_110_1_100011101111;
      patterns[51071] = 29'b1_100011101111_111_1_100011101111;
      patterns[51072] = 29'b1_100011110000_000_1_100011110000;
      patterns[51073] = 29'b1_100011110000_001_1_110000100011;
      patterns[51074] = 29'b1_100011110000_010_1_000111100001;
      patterns[51075] = 29'b1_100011110000_011_0_001111000011;
      patterns[51076] = 29'b1_100011110000_100_0_110001111000;
      patterns[51077] = 29'b1_100011110000_101_0_011000111100;
      patterns[51078] = 29'b1_100011110000_110_1_100011110000;
      patterns[51079] = 29'b1_100011110000_111_1_100011110000;
      patterns[51080] = 29'b1_100011110001_000_1_100011110001;
      patterns[51081] = 29'b1_100011110001_001_1_110001100011;
      patterns[51082] = 29'b1_100011110001_010_1_000111100011;
      patterns[51083] = 29'b1_100011110001_011_0_001111000111;
      patterns[51084] = 29'b1_100011110001_100_1_110001111000;
      patterns[51085] = 29'b1_100011110001_101_0_111000111100;
      patterns[51086] = 29'b1_100011110001_110_1_100011110001;
      patterns[51087] = 29'b1_100011110001_111_1_100011110001;
      patterns[51088] = 29'b1_100011110010_000_1_100011110010;
      patterns[51089] = 29'b1_100011110010_001_1_110010100011;
      patterns[51090] = 29'b1_100011110010_010_1_000111100101;
      patterns[51091] = 29'b1_100011110010_011_0_001111001011;
      patterns[51092] = 29'b1_100011110010_100_0_110001111001;
      patterns[51093] = 29'b1_100011110010_101_1_011000111100;
      patterns[51094] = 29'b1_100011110010_110_1_100011110010;
      patterns[51095] = 29'b1_100011110010_111_1_100011110010;
      patterns[51096] = 29'b1_100011110011_000_1_100011110011;
      patterns[51097] = 29'b1_100011110011_001_1_110011100011;
      patterns[51098] = 29'b1_100011110011_010_1_000111100111;
      patterns[51099] = 29'b1_100011110011_011_0_001111001111;
      patterns[51100] = 29'b1_100011110011_100_1_110001111001;
      patterns[51101] = 29'b1_100011110011_101_1_111000111100;
      patterns[51102] = 29'b1_100011110011_110_1_100011110011;
      patterns[51103] = 29'b1_100011110011_111_1_100011110011;
      patterns[51104] = 29'b1_100011110100_000_1_100011110100;
      patterns[51105] = 29'b1_100011110100_001_1_110100100011;
      patterns[51106] = 29'b1_100011110100_010_1_000111101001;
      patterns[51107] = 29'b1_100011110100_011_0_001111010011;
      patterns[51108] = 29'b1_100011110100_100_0_110001111010;
      patterns[51109] = 29'b1_100011110100_101_0_011000111101;
      patterns[51110] = 29'b1_100011110100_110_1_100011110100;
      patterns[51111] = 29'b1_100011110100_111_1_100011110100;
      patterns[51112] = 29'b1_100011110101_000_1_100011110101;
      patterns[51113] = 29'b1_100011110101_001_1_110101100011;
      patterns[51114] = 29'b1_100011110101_010_1_000111101011;
      patterns[51115] = 29'b1_100011110101_011_0_001111010111;
      patterns[51116] = 29'b1_100011110101_100_1_110001111010;
      patterns[51117] = 29'b1_100011110101_101_0_111000111101;
      patterns[51118] = 29'b1_100011110101_110_1_100011110101;
      patterns[51119] = 29'b1_100011110101_111_1_100011110101;
      patterns[51120] = 29'b1_100011110110_000_1_100011110110;
      patterns[51121] = 29'b1_100011110110_001_1_110110100011;
      patterns[51122] = 29'b1_100011110110_010_1_000111101101;
      patterns[51123] = 29'b1_100011110110_011_0_001111011011;
      patterns[51124] = 29'b1_100011110110_100_0_110001111011;
      patterns[51125] = 29'b1_100011110110_101_1_011000111101;
      patterns[51126] = 29'b1_100011110110_110_1_100011110110;
      patterns[51127] = 29'b1_100011110110_111_1_100011110110;
      patterns[51128] = 29'b1_100011110111_000_1_100011110111;
      patterns[51129] = 29'b1_100011110111_001_1_110111100011;
      patterns[51130] = 29'b1_100011110111_010_1_000111101111;
      patterns[51131] = 29'b1_100011110111_011_0_001111011111;
      patterns[51132] = 29'b1_100011110111_100_1_110001111011;
      patterns[51133] = 29'b1_100011110111_101_1_111000111101;
      patterns[51134] = 29'b1_100011110111_110_1_100011110111;
      patterns[51135] = 29'b1_100011110111_111_1_100011110111;
      patterns[51136] = 29'b1_100011111000_000_1_100011111000;
      patterns[51137] = 29'b1_100011111000_001_1_111000100011;
      patterns[51138] = 29'b1_100011111000_010_1_000111110001;
      patterns[51139] = 29'b1_100011111000_011_0_001111100011;
      patterns[51140] = 29'b1_100011111000_100_0_110001111100;
      patterns[51141] = 29'b1_100011111000_101_0_011000111110;
      patterns[51142] = 29'b1_100011111000_110_1_100011111000;
      patterns[51143] = 29'b1_100011111000_111_1_100011111000;
      patterns[51144] = 29'b1_100011111001_000_1_100011111001;
      patterns[51145] = 29'b1_100011111001_001_1_111001100011;
      patterns[51146] = 29'b1_100011111001_010_1_000111110011;
      patterns[51147] = 29'b1_100011111001_011_0_001111100111;
      patterns[51148] = 29'b1_100011111001_100_1_110001111100;
      patterns[51149] = 29'b1_100011111001_101_0_111000111110;
      patterns[51150] = 29'b1_100011111001_110_1_100011111001;
      patterns[51151] = 29'b1_100011111001_111_1_100011111001;
      patterns[51152] = 29'b1_100011111010_000_1_100011111010;
      patterns[51153] = 29'b1_100011111010_001_1_111010100011;
      patterns[51154] = 29'b1_100011111010_010_1_000111110101;
      patterns[51155] = 29'b1_100011111010_011_0_001111101011;
      patterns[51156] = 29'b1_100011111010_100_0_110001111101;
      patterns[51157] = 29'b1_100011111010_101_1_011000111110;
      patterns[51158] = 29'b1_100011111010_110_1_100011111010;
      patterns[51159] = 29'b1_100011111010_111_1_100011111010;
      patterns[51160] = 29'b1_100011111011_000_1_100011111011;
      patterns[51161] = 29'b1_100011111011_001_1_111011100011;
      patterns[51162] = 29'b1_100011111011_010_1_000111110111;
      patterns[51163] = 29'b1_100011111011_011_0_001111101111;
      patterns[51164] = 29'b1_100011111011_100_1_110001111101;
      patterns[51165] = 29'b1_100011111011_101_1_111000111110;
      patterns[51166] = 29'b1_100011111011_110_1_100011111011;
      patterns[51167] = 29'b1_100011111011_111_1_100011111011;
      patterns[51168] = 29'b1_100011111100_000_1_100011111100;
      patterns[51169] = 29'b1_100011111100_001_1_111100100011;
      patterns[51170] = 29'b1_100011111100_010_1_000111111001;
      patterns[51171] = 29'b1_100011111100_011_0_001111110011;
      patterns[51172] = 29'b1_100011111100_100_0_110001111110;
      patterns[51173] = 29'b1_100011111100_101_0_011000111111;
      patterns[51174] = 29'b1_100011111100_110_1_100011111100;
      patterns[51175] = 29'b1_100011111100_111_1_100011111100;
      patterns[51176] = 29'b1_100011111101_000_1_100011111101;
      patterns[51177] = 29'b1_100011111101_001_1_111101100011;
      patterns[51178] = 29'b1_100011111101_010_1_000111111011;
      patterns[51179] = 29'b1_100011111101_011_0_001111110111;
      patterns[51180] = 29'b1_100011111101_100_1_110001111110;
      patterns[51181] = 29'b1_100011111101_101_0_111000111111;
      patterns[51182] = 29'b1_100011111101_110_1_100011111101;
      patterns[51183] = 29'b1_100011111101_111_1_100011111101;
      patterns[51184] = 29'b1_100011111110_000_1_100011111110;
      patterns[51185] = 29'b1_100011111110_001_1_111110100011;
      patterns[51186] = 29'b1_100011111110_010_1_000111111101;
      patterns[51187] = 29'b1_100011111110_011_0_001111111011;
      patterns[51188] = 29'b1_100011111110_100_0_110001111111;
      patterns[51189] = 29'b1_100011111110_101_1_011000111111;
      patterns[51190] = 29'b1_100011111110_110_1_100011111110;
      patterns[51191] = 29'b1_100011111110_111_1_100011111110;
      patterns[51192] = 29'b1_100011111111_000_1_100011111111;
      patterns[51193] = 29'b1_100011111111_001_1_111111100011;
      patterns[51194] = 29'b1_100011111111_010_1_000111111111;
      patterns[51195] = 29'b1_100011111111_011_0_001111111111;
      patterns[51196] = 29'b1_100011111111_100_1_110001111111;
      patterns[51197] = 29'b1_100011111111_101_1_111000111111;
      patterns[51198] = 29'b1_100011111111_110_1_100011111111;
      patterns[51199] = 29'b1_100011111111_111_1_100011111111;
      patterns[51200] = 29'b1_100100000000_000_1_100100000000;
      patterns[51201] = 29'b1_100100000000_001_1_000000100100;
      patterns[51202] = 29'b1_100100000000_010_1_001000000001;
      patterns[51203] = 29'b1_100100000000_011_0_010000000011;
      patterns[51204] = 29'b1_100100000000_100_0_110010000000;
      patterns[51205] = 29'b1_100100000000_101_0_011001000000;
      patterns[51206] = 29'b1_100100000000_110_1_100100000000;
      patterns[51207] = 29'b1_100100000000_111_1_100100000000;
      patterns[51208] = 29'b1_100100000001_000_1_100100000001;
      patterns[51209] = 29'b1_100100000001_001_1_000001100100;
      patterns[51210] = 29'b1_100100000001_010_1_001000000011;
      patterns[51211] = 29'b1_100100000001_011_0_010000000111;
      patterns[51212] = 29'b1_100100000001_100_1_110010000000;
      patterns[51213] = 29'b1_100100000001_101_0_111001000000;
      patterns[51214] = 29'b1_100100000001_110_1_100100000001;
      patterns[51215] = 29'b1_100100000001_111_1_100100000001;
      patterns[51216] = 29'b1_100100000010_000_1_100100000010;
      patterns[51217] = 29'b1_100100000010_001_1_000010100100;
      patterns[51218] = 29'b1_100100000010_010_1_001000000101;
      patterns[51219] = 29'b1_100100000010_011_0_010000001011;
      patterns[51220] = 29'b1_100100000010_100_0_110010000001;
      patterns[51221] = 29'b1_100100000010_101_1_011001000000;
      patterns[51222] = 29'b1_100100000010_110_1_100100000010;
      patterns[51223] = 29'b1_100100000010_111_1_100100000010;
      patterns[51224] = 29'b1_100100000011_000_1_100100000011;
      patterns[51225] = 29'b1_100100000011_001_1_000011100100;
      patterns[51226] = 29'b1_100100000011_010_1_001000000111;
      patterns[51227] = 29'b1_100100000011_011_0_010000001111;
      patterns[51228] = 29'b1_100100000011_100_1_110010000001;
      patterns[51229] = 29'b1_100100000011_101_1_111001000000;
      patterns[51230] = 29'b1_100100000011_110_1_100100000011;
      patterns[51231] = 29'b1_100100000011_111_1_100100000011;
      patterns[51232] = 29'b1_100100000100_000_1_100100000100;
      patterns[51233] = 29'b1_100100000100_001_1_000100100100;
      patterns[51234] = 29'b1_100100000100_010_1_001000001001;
      patterns[51235] = 29'b1_100100000100_011_0_010000010011;
      patterns[51236] = 29'b1_100100000100_100_0_110010000010;
      patterns[51237] = 29'b1_100100000100_101_0_011001000001;
      patterns[51238] = 29'b1_100100000100_110_1_100100000100;
      patterns[51239] = 29'b1_100100000100_111_1_100100000100;
      patterns[51240] = 29'b1_100100000101_000_1_100100000101;
      patterns[51241] = 29'b1_100100000101_001_1_000101100100;
      patterns[51242] = 29'b1_100100000101_010_1_001000001011;
      patterns[51243] = 29'b1_100100000101_011_0_010000010111;
      patterns[51244] = 29'b1_100100000101_100_1_110010000010;
      patterns[51245] = 29'b1_100100000101_101_0_111001000001;
      patterns[51246] = 29'b1_100100000101_110_1_100100000101;
      patterns[51247] = 29'b1_100100000101_111_1_100100000101;
      patterns[51248] = 29'b1_100100000110_000_1_100100000110;
      patterns[51249] = 29'b1_100100000110_001_1_000110100100;
      patterns[51250] = 29'b1_100100000110_010_1_001000001101;
      patterns[51251] = 29'b1_100100000110_011_0_010000011011;
      patterns[51252] = 29'b1_100100000110_100_0_110010000011;
      patterns[51253] = 29'b1_100100000110_101_1_011001000001;
      patterns[51254] = 29'b1_100100000110_110_1_100100000110;
      patterns[51255] = 29'b1_100100000110_111_1_100100000110;
      patterns[51256] = 29'b1_100100000111_000_1_100100000111;
      patterns[51257] = 29'b1_100100000111_001_1_000111100100;
      patterns[51258] = 29'b1_100100000111_010_1_001000001111;
      patterns[51259] = 29'b1_100100000111_011_0_010000011111;
      patterns[51260] = 29'b1_100100000111_100_1_110010000011;
      patterns[51261] = 29'b1_100100000111_101_1_111001000001;
      patterns[51262] = 29'b1_100100000111_110_1_100100000111;
      patterns[51263] = 29'b1_100100000111_111_1_100100000111;
      patterns[51264] = 29'b1_100100001000_000_1_100100001000;
      patterns[51265] = 29'b1_100100001000_001_1_001000100100;
      patterns[51266] = 29'b1_100100001000_010_1_001000010001;
      patterns[51267] = 29'b1_100100001000_011_0_010000100011;
      patterns[51268] = 29'b1_100100001000_100_0_110010000100;
      patterns[51269] = 29'b1_100100001000_101_0_011001000010;
      patterns[51270] = 29'b1_100100001000_110_1_100100001000;
      patterns[51271] = 29'b1_100100001000_111_1_100100001000;
      patterns[51272] = 29'b1_100100001001_000_1_100100001001;
      patterns[51273] = 29'b1_100100001001_001_1_001001100100;
      patterns[51274] = 29'b1_100100001001_010_1_001000010011;
      patterns[51275] = 29'b1_100100001001_011_0_010000100111;
      patterns[51276] = 29'b1_100100001001_100_1_110010000100;
      patterns[51277] = 29'b1_100100001001_101_0_111001000010;
      patterns[51278] = 29'b1_100100001001_110_1_100100001001;
      patterns[51279] = 29'b1_100100001001_111_1_100100001001;
      patterns[51280] = 29'b1_100100001010_000_1_100100001010;
      patterns[51281] = 29'b1_100100001010_001_1_001010100100;
      patterns[51282] = 29'b1_100100001010_010_1_001000010101;
      patterns[51283] = 29'b1_100100001010_011_0_010000101011;
      patterns[51284] = 29'b1_100100001010_100_0_110010000101;
      patterns[51285] = 29'b1_100100001010_101_1_011001000010;
      patterns[51286] = 29'b1_100100001010_110_1_100100001010;
      patterns[51287] = 29'b1_100100001010_111_1_100100001010;
      patterns[51288] = 29'b1_100100001011_000_1_100100001011;
      patterns[51289] = 29'b1_100100001011_001_1_001011100100;
      patterns[51290] = 29'b1_100100001011_010_1_001000010111;
      patterns[51291] = 29'b1_100100001011_011_0_010000101111;
      patterns[51292] = 29'b1_100100001011_100_1_110010000101;
      patterns[51293] = 29'b1_100100001011_101_1_111001000010;
      patterns[51294] = 29'b1_100100001011_110_1_100100001011;
      patterns[51295] = 29'b1_100100001011_111_1_100100001011;
      patterns[51296] = 29'b1_100100001100_000_1_100100001100;
      patterns[51297] = 29'b1_100100001100_001_1_001100100100;
      patterns[51298] = 29'b1_100100001100_010_1_001000011001;
      patterns[51299] = 29'b1_100100001100_011_0_010000110011;
      patterns[51300] = 29'b1_100100001100_100_0_110010000110;
      patterns[51301] = 29'b1_100100001100_101_0_011001000011;
      patterns[51302] = 29'b1_100100001100_110_1_100100001100;
      patterns[51303] = 29'b1_100100001100_111_1_100100001100;
      patterns[51304] = 29'b1_100100001101_000_1_100100001101;
      patterns[51305] = 29'b1_100100001101_001_1_001101100100;
      patterns[51306] = 29'b1_100100001101_010_1_001000011011;
      patterns[51307] = 29'b1_100100001101_011_0_010000110111;
      patterns[51308] = 29'b1_100100001101_100_1_110010000110;
      patterns[51309] = 29'b1_100100001101_101_0_111001000011;
      patterns[51310] = 29'b1_100100001101_110_1_100100001101;
      patterns[51311] = 29'b1_100100001101_111_1_100100001101;
      patterns[51312] = 29'b1_100100001110_000_1_100100001110;
      patterns[51313] = 29'b1_100100001110_001_1_001110100100;
      patterns[51314] = 29'b1_100100001110_010_1_001000011101;
      patterns[51315] = 29'b1_100100001110_011_0_010000111011;
      patterns[51316] = 29'b1_100100001110_100_0_110010000111;
      patterns[51317] = 29'b1_100100001110_101_1_011001000011;
      patterns[51318] = 29'b1_100100001110_110_1_100100001110;
      patterns[51319] = 29'b1_100100001110_111_1_100100001110;
      patterns[51320] = 29'b1_100100001111_000_1_100100001111;
      patterns[51321] = 29'b1_100100001111_001_1_001111100100;
      patterns[51322] = 29'b1_100100001111_010_1_001000011111;
      patterns[51323] = 29'b1_100100001111_011_0_010000111111;
      patterns[51324] = 29'b1_100100001111_100_1_110010000111;
      patterns[51325] = 29'b1_100100001111_101_1_111001000011;
      patterns[51326] = 29'b1_100100001111_110_1_100100001111;
      patterns[51327] = 29'b1_100100001111_111_1_100100001111;
      patterns[51328] = 29'b1_100100010000_000_1_100100010000;
      patterns[51329] = 29'b1_100100010000_001_1_010000100100;
      patterns[51330] = 29'b1_100100010000_010_1_001000100001;
      patterns[51331] = 29'b1_100100010000_011_0_010001000011;
      patterns[51332] = 29'b1_100100010000_100_0_110010001000;
      patterns[51333] = 29'b1_100100010000_101_0_011001000100;
      patterns[51334] = 29'b1_100100010000_110_1_100100010000;
      patterns[51335] = 29'b1_100100010000_111_1_100100010000;
      patterns[51336] = 29'b1_100100010001_000_1_100100010001;
      patterns[51337] = 29'b1_100100010001_001_1_010001100100;
      patterns[51338] = 29'b1_100100010001_010_1_001000100011;
      patterns[51339] = 29'b1_100100010001_011_0_010001000111;
      patterns[51340] = 29'b1_100100010001_100_1_110010001000;
      patterns[51341] = 29'b1_100100010001_101_0_111001000100;
      patterns[51342] = 29'b1_100100010001_110_1_100100010001;
      patterns[51343] = 29'b1_100100010001_111_1_100100010001;
      patterns[51344] = 29'b1_100100010010_000_1_100100010010;
      patterns[51345] = 29'b1_100100010010_001_1_010010100100;
      patterns[51346] = 29'b1_100100010010_010_1_001000100101;
      patterns[51347] = 29'b1_100100010010_011_0_010001001011;
      patterns[51348] = 29'b1_100100010010_100_0_110010001001;
      patterns[51349] = 29'b1_100100010010_101_1_011001000100;
      patterns[51350] = 29'b1_100100010010_110_1_100100010010;
      patterns[51351] = 29'b1_100100010010_111_1_100100010010;
      patterns[51352] = 29'b1_100100010011_000_1_100100010011;
      patterns[51353] = 29'b1_100100010011_001_1_010011100100;
      patterns[51354] = 29'b1_100100010011_010_1_001000100111;
      patterns[51355] = 29'b1_100100010011_011_0_010001001111;
      patterns[51356] = 29'b1_100100010011_100_1_110010001001;
      patterns[51357] = 29'b1_100100010011_101_1_111001000100;
      patterns[51358] = 29'b1_100100010011_110_1_100100010011;
      patterns[51359] = 29'b1_100100010011_111_1_100100010011;
      patterns[51360] = 29'b1_100100010100_000_1_100100010100;
      patterns[51361] = 29'b1_100100010100_001_1_010100100100;
      patterns[51362] = 29'b1_100100010100_010_1_001000101001;
      patterns[51363] = 29'b1_100100010100_011_0_010001010011;
      patterns[51364] = 29'b1_100100010100_100_0_110010001010;
      patterns[51365] = 29'b1_100100010100_101_0_011001000101;
      patterns[51366] = 29'b1_100100010100_110_1_100100010100;
      patterns[51367] = 29'b1_100100010100_111_1_100100010100;
      patterns[51368] = 29'b1_100100010101_000_1_100100010101;
      patterns[51369] = 29'b1_100100010101_001_1_010101100100;
      patterns[51370] = 29'b1_100100010101_010_1_001000101011;
      patterns[51371] = 29'b1_100100010101_011_0_010001010111;
      patterns[51372] = 29'b1_100100010101_100_1_110010001010;
      patterns[51373] = 29'b1_100100010101_101_0_111001000101;
      patterns[51374] = 29'b1_100100010101_110_1_100100010101;
      patterns[51375] = 29'b1_100100010101_111_1_100100010101;
      patterns[51376] = 29'b1_100100010110_000_1_100100010110;
      patterns[51377] = 29'b1_100100010110_001_1_010110100100;
      patterns[51378] = 29'b1_100100010110_010_1_001000101101;
      patterns[51379] = 29'b1_100100010110_011_0_010001011011;
      patterns[51380] = 29'b1_100100010110_100_0_110010001011;
      patterns[51381] = 29'b1_100100010110_101_1_011001000101;
      patterns[51382] = 29'b1_100100010110_110_1_100100010110;
      patterns[51383] = 29'b1_100100010110_111_1_100100010110;
      patterns[51384] = 29'b1_100100010111_000_1_100100010111;
      patterns[51385] = 29'b1_100100010111_001_1_010111100100;
      patterns[51386] = 29'b1_100100010111_010_1_001000101111;
      patterns[51387] = 29'b1_100100010111_011_0_010001011111;
      patterns[51388] = 29'b1_100100010111_100_1_110010001011;
      patterns[51389] = 29'b1_100100010111_101_1_111001000101;
      patterns[51390] = 29'b1_100100010111_110_1_100100010111;
      patterns[51391] = 29'b1_100100010111_111_1_100100010111;
      patterns[51392] = 29'b1_100100011000_000_1_100100011000;
      patterns[51393] = 29'b1_100100011000_001_1_011000100100;
      patterns[51394] = 29'b1_100100011000_010_1_001000110001;
      patterns[51395] = 29'b1_100100011000_011_0_010001100011;
      patterns[51396] = 29'b1_100100011000_100_0_110010001100;
      patterns[51397] = 29'b1_100100011000_101_0_011001000110;
      patterns[51398] = 29'b1_100100011000_110_1_100100011000;
      patterns[51399] = 29'b1_100100011000_111_1_100100011000;
      patterns[51400] = 29'b1_100100011001_000_1_100100011001;
      patterns[51401] = 29'b1_100100011001_001_1_011001100100;
      patterns[51402] = 29'b1_100100011001_010_1_001000110011;
      patterns[51403] = 29'b1_100100011001_011_0_010001100111;
      patterns[51404] = 29'b1_100100011001_100_1_110010001100;
      patterns[51405] = 29'b1_100100011001_101_0_111001000110;
      patterns[51406] = 29'b1_100100011001_110_1_100100011001;
      patterns[51407] = 29'b1_100100011001_111_1_100100011001;
      patterns[51408] = 29'b1_100100011010_000_1_100100011010;
      patterns[51409] = 29'b1_100100011010_001_1_011010100100;
      patterns[51410] = 29'b1_100100011010_010_1_001000110101;
      patterns[51411] = 29'b1_100100011010_011_0_010001101011;
      patterns[51412] = 29'b1_100100011010_100_0_110010001101;
      patterns[51413] = 29'b1_100100011010_101_1_011001000110;
      patterns[51414] = 29'b1_100100011010_110_1_100100011010;
      patterns[51415] = 29'b1_100100011010_111_1_100100011010;
      patterns[51416] = 29'b1_100100011011_000_1_100100011011;
      patterns[51417] = 29'b1_100100011011_001_1_011011100100;
      patterns[51418] = 29'b1_100100011011_010_1_001000110111;
      patterns[51419] = 29'b1_100100011011_011_0_010001101111;
      patterns[51420] = 29'b1_100100011011_100_1_110010001101;
      patterns[51421] = 29'b1_100100011011_101_1_111001000110;
      patterns[51422] = 29'b1_100100011011_110_1_100100011011;
      patterns[51423] = 29'b1_100100011011_111_1_100100011011;
      patterns[51424] = 29'b1_100100011100_000_1_100100011100;
      patterns[51425] = 29'b1_100100011100_001_1_011100100100;
      patterns[51426] = 29'b1_100100011100_010_1_001000111001;
      patterns[51427] = 29'b1_100100011100_011_0_010001110011;
      patterns[51428] = 29'b1_100100011100_100_0_110010001110;
      patterns[51429] = 29'b1_100100011100_101_0_011001000111;
      patterns[51430] = 29'b1_100100011100_110_1_100100011100;
      patterns[51431] = 29'b1_100100011100_111_1_100100011100;
      patterns[51432] = 29'b1_100100011101_000_1_100100011101;
      patterns[51433] = 29'b1_100100011101_001_1_011101100100;
      patterns[51434] = 29'b1_100100011101_010_1_001000111011;
      patterns[51435] = 29'b1_100100011101_011_0_010001110111;
      patterns[51436] = 29'b1_100100011101_100_1_110010001110;
      patterns[51437] = 29'b1_100100011101_101_0_111001000111;
      patterns[51438] = 29'b1_100100011101_110_1_100100011101;
      patterns[51439] = 29'b1_100100011101_111_1_100100011101;
      patterns[51440] = 29'b1_100100011110_000_1_100100011110;
      patterns[51441] = 29'b1_100100011110_001_1_011110100100;
      patterns[51442] = 29'b1_100100011110_010_1_001000111101;
      patterns[51443] = 29'b1_100100011110_011_0_010001111011;
      patterns[51444] = 29'b1_100100011110_100_0_110010001111;
      patterns[51445] = 29'b1_100100011110_101_1_011001000111;
      patterns[51446] = 29'b1_100100011110_110_1_100100011110;
      patterns[51447] = 29'b1_100100011110_111_1_100100011110;
      patterns[51448] = 29'b1_100100011111_000_1_100100011111;
      patterns[51449] = 29'b1_100100011111_001_1_011111100100;
      patterns[51450] = 29'b1_100100011111_010_1_001000111111;
      patterns[51451] = 29'b1_100100011111_011_0_010001111111;
      patterns[51452] = 29'b1_100100011111_100_1_110010001111;
      patterns[51453] = 29'b1_100100011111_101_1_111001000111;
      patterns[51454] = 29'b1_100100011111_110_1_100100011111;
      patterns[51455] = 29'b1_100100011111_111_1_100100011111;
      patterns[51456] = 29'b1_100100100000_000_1_100100100000;
      patterns[51457] = 29'b1_100100100000_001_1_100000100100;
      patterns[51458] = 29'b1_100100100000_010_1_001001000001;
      patterns[51459] = 29'b1_100100100000_011_0_010010000011;
      patterns[51460] = 29'b1_100100100000_100_0_110010010000;
      patterns[51461] = 29'b1_100100100000_101_0_011001001000;
      patterns[51462] = 29'b1_100100100000_110_1_100100100000;
      patterns[51463] = 29'b1_100100100000_111_1_100100100000;
      patterns[51464] = 29'b1_100100100001_000_1_100100100001;
      patterns[51465] = 29'b1_100100100001_001_1_100001100100;
      patterns[51466] = 29'b1_100100100001_010_1_001001000011;
      patterns[51467] = 29'b1_100100100001_011_0_010010000111;
      patterns[51468] = 29'b1_100100100001_100_1_110010010000;
      patterns[51469] = 29'b1_100100100001_101_0_111001001000;
      patterns[51470] = 29'b1_100100100001_110_1_100100100001;
      patterns[51471] = 29'b1_100100100001_111_1_100100100001;
      patterns[51472] = 29'b1_100100100010_000_1_100100100010;
      patterns[51473] = 29'b1_100100100010_001_1_100010100100;
      patterns[51474] = 29'b1_100100100010_010_1_001001000101;
      patterns[51475] = 29'b1_100100100010_011_0_010010001011;
      patterns[51476] = 29'b1_100100100010_100_0_110010010001;
      patterns[51477] = 29'b1_100100100010_101_1_011001001000;
      patterns[51478] = 29'b1_100100100010_110_1_100100100010;
      patterns[51479] = 29'b1_100100100010_111_1_100100100010;
      patterns[51480] = 29'b1_100100100011_000_1_100100100011;
      patterns[51481] = 29'b1_100100100011_001_1_100011100100;
      patterns[51482] = 29'b1_100100100011_010_1_001001000111;
      patterns[51483] = 29'b1_100100100011_011_0_010010001111;
      patterns[51484] = 29'b1_100100100011_100_1_110010010001;
      patterns[51485] = 29'b1_100100100011_101_1_111001001000;
      patterns[51486] = 29'b1_100100100011_110_1_100100100011;
      patterns[51487] = 29'b1_100100100011_111_1_100100100011;
      patterns[51488] = 29'b1_100100100100_000_1_100100100100;
      patterns[51489] = 29'b1_100100100100_001_1_100100100100;
      patterns[51490] = 29'b1_100100100100_010_1_001001001001;
      patterns[51491] = 29'b1_100100100100_011_0_010010010011;
      patterns[51492] = 29'b1_100100100100_100_0_110010010010;
      patterns[51493] = 29'b1_100100100100_101_0_011001001001;
      patterns[51494] = 29'b1_100100100100_110_1_100100100100;
      patterns[51495] = 29'b1_100100100100_111_1_100100100100;
      patterns[51496] = 29'b1_100100100101_000_1_100100100101;
      patterns[51497] = 29'b1_100100100101_001_1_100101100100;
      patterns[51498] = 29'b1_100100100101_010_1_001001001011;
      patterns[51499] = 29'b1_100100100101_011_0_010010010111;
      patterns[51500] = 29'b1_100100100101_100_1_110010010010;
      patterns[51501] = 29'b1_100100100101_101_0_111001001001;
      patterns[51502] = 29'b1_100100100101_110_1_100100100101;
      patterns[51503] = 29'b1_100100100101_111_1_100100100101;
      patterns[51504] = 29'b1_100100100110_000_1_100100100110;
      patterns[51505] = 29'b1_100100100110_001_1_100110100100;
      patterns[51506] = 29'b1_100100100110_010_1_001001001101;
      patterns[51507] = 29'b1_100100100110_011_0_010010011011;
      patterns[51508] = 29'b1_100100100110_100_0_110010010011;
      patterns[51509] = 29'b1_100100100110_101_1_011001001001;
      patterns[51510] = 29'b1_100100100110_110_1_100100100110;
      patterns[51511] = 29'b1_100100100110_111_1_100100100110;
      patterns[51512] = 29'b1_100100100111_000_1_100100100111;
      patterns[51513] = 29'b1_100100100111_001_1_100111100100;
      patterns[51514] = 29'b1_100100100111_010_1_001001001111;
      patterns[51515] = 29'b1_100100100111_011_0_010010011111;
      patterns[51516] = 29'b1_100100100111_100_1_110010010011;
      patterns[51517] = 29'b1_100100100111_101_1_111001001001;
      patterns[51518] = 29'b1_100100100111_110_1_100100100111;
      patterns[51519] = 29'b1_100100100111_111_1_100100100111;
      patterns[51520] = 29'b1_100100101000_000_1_100100101000;
      patterns[51521] = 29'b1_100100101000_001_1_101000100100;
      patterns[51522] = 29'b1_100100101000_010_1_001001010001;
      patterns[51523] = 29'b1_100100101000_011_0_010010100011;
      patterns[51524] = 29'b1_100100101000_100_0_110010010100;
      patterns[51525] = 29'b1_100100101000_101_0_011001001010;
      patterns[51526] = 29'b1_100100101000_110_1_100100101000;
      patterns[51527] = 29'b1_100100101000_111_1_100100101000;
      patterns[51528] = 29'b1_100100101001_000_1_100100101001;
      patterns[51529] = 29'b1_100100101001_001_1_101001100100;
      patterns[51530] = 29'b1_100100101001_010_1_001001010011;
      patterns[51531] = 29'b1_100100101001_011_0_010010100111;
      patterns[51532] = 29'b1_100100101001_100_1_110010010100;
      patterns[51533] = 29'b1_100100101001_101_0_111001001010;
      patterns[51534] = 29'b1_100100101001_110_1_100100101001;
      patterns[51535] = 29'b1_100100101001_111_1_100100101001;
      patterns[51536] = 29'b1_100100101010_000_1_100100101010;
      patterns[51537] = 29'b1_100100101010_001_1_101010100100;
      patterns[51538] = 29'b1_100100101010_010_1_001001010101;
      patterns[51539] = 29'b1_100100101010_011_0_010010101011;
      patterns[51540] = 29'b1_100100101010_100_0_110010010101;
      patterns[51541] = 29'b1_100100101010_101_1_011001001010;
      patterns[51542] = 29'b1_100100101010_110_1_100100101010;
      patterns[51543] = 29'b1_100100101010_111_1_100100101010;
      patterns[51544] = 29'b1_100100101011_000_1_100100101011;
      patterns[51545] = 29'b1_100100101011_001_1_101011100100;
      patterns[51546] = 29'b1_100100101011_010_1_001001010111;
      patterns[51547] = 29'b1_100100101011_011_0_010010101111;
      patterns[51548] = 29'b1_100100101011_100_1_110010010101;
      patterns[51549] = 29'b1_100100101011_101_1_111001001010;
      patterns[51550] = 29'b1_100100101011_110_1_100100101011;
      patterns[51551] = 29'b1_100100101011_111_1_100100101011;
      patterns[51552] = 29'b1_100100101100_000_1_100100101100;
      patterns[51553] = 29'b1_100100101100_001_1_101100100100;
      patterns[51554] = 29'b1_100100101100_010_1_001001011001;
      patterns[51555] = 29'b1_100100101100_011_0_010010110011;
      patterns[51556] = 29'b1_100100101100_100_0_110010010110;
      patterns[51557] = 29'b1_100100101100_101_0_011001001011;
      patterns[51558] = 29'b1_100100101100_110_1_100100101100;
      patterns[51559] = 29'b1_100100101100_111_1_100100101100;
      patterns[51560] = 29'b1_100100101101_000_1_100100101101;
      patterns[51561] = 29'b1_100100101101_001_1_101101100100;
      patterns[51562] = 29'b1_100100101101_010_1_001001011011;
      patterns[51563] = 29'b1_100100101101_011_0_010010110111;
      patterns[51564] = 29'b1_100100101101_100_1_110010010110;
      patterns[51565] = 29'b1_100100101101_101_0_111001001011;
      patterns[51566] = 29'b1_100100101101_110_1_100100101101;
      patterns[51567] = 29'b1_100100101101_111_1_100100101101;
      patterns[51568] = 29'b1_100100101110_000_1_100100101110;
      patterns[51569] = 29'b1_100100101110_001_1_101110100100;
      patterns[51570] = 29'b1_100100101110_010_1_001001011101;
      patterns[51571] = 29'b1_100100101110_011_0_010010111011;
      patterns[51572] = 29'b1_100100101110_100_0_110010010111;
      patterns[51573] = 29'b1_100100101110_101_1_011001001011;
      patterns[51574] = 29'b1_100100101110_110_1_100100101110;
      patterns[51575] = 29'b1_100100101110_111_1_100100101110;
      patterns[51576] = 29'b1_100100101111_000_1_100100101111;
      patterns[51577] = 29'b1_100100101111_001_1_101111100100;
      patterns[51578] = 29'b1_100100101111_010_1_001001011111;
      patterns[51579] = 29'b1_100100101111_011_0_010010111111;
      patterns[51580] = 29'b1_100100101111_100_1_110010010111;
      patterns[51581] = 29'b1_100100101111_101_1_111001001011;
      patterns[51582] = 29'b1_100100101111_110_1_100100101111;
      patterns[51583] = 29'b1_100100101111_111_1_100100101111;
      patterns[51584] = 29'b1_100100110000_000_1_100100110000;
      patterns[51585] = 29'b1_100100110000_001_1_110000100100;
      patterns[51586] = 29'b1_100100110000_010_1_001001100001;
      patterns[51587] = 29'b1_100100110000_011_0_010011000011;
      patterns[51588] = 29'b1_100100110000_100_0_110010011000;
      patterns[51589] = 29'b1_100100110000_101_0_011001001100;
      patterns[51590] = 29'b1_100100110000_110_1_100100110000;
      patterns[51591] = 29'b1_100100110000_111_1_100100110000;
      patterns[51592] = 29'b1_100100110001_000_1_100100110001;
      patterns[51593] = 29'b1_100100110001_001_1_110001100100;
      patterns[51594] = 29'b1_100100110001_010_1_001001100011;
      patterns[51595] = 29'b1_100100110001_011_0_010011000111;
      patterns[51596] = 29'b1_100100110001_100_1_110010011000;
      patterns[51597] = 29'b1_100100110001_101_0_111001001100;
      patterns[51598] = 29'b1_100100110001_110_1_100100110001;
      patterns[51599] = 29'b1_100100110001_111_1_100100110001;
      patterns[51600] = 29'b1_100100110010_000_1_100100110010;
      patterns[51601] = 29'b1_100100110010_001_1_110010100100;
      patterns[51602] = 29'b1_100100110010_010_1_001001100101;
      patterns[51603] = 29'b1_100100110010_011_0_010011001011;
      patterns[51604] = 29'b1_100100110010_100_0_110010011001;
      patterns[51605] = 29'b1_100100110010_101_1_011001001100;
      patterns[51606] = 29'b1_100100110010_110_1_100100110010;
      patterns[51607] = 29'b1_100100110010_111_1_100100110010;
      patterns[51608] = 29'b1_100100110011_000_1_100100110011;
      patterns[51609] = 29'b1_100100110011_001_1_110011100100;
      patterns[51610] = 29'b1_100100110011_010_1_001001100111;
      patterns[51611] = 29'b1_100100110011_011_0_010011001111;
      patterns[51612] = 29'b1_100100110011_100_1_110010011001;
      patterns[51613] = 29'b1_100100110011_101_1_111001001100;
      patterns[51614] = 29'b1_100100110011_110_1_100100110011;
      patterns[51615] = 29'b1_100100110011_111_1_100100110011;
      patterns[51616] = 29'b1_100100110100_000_1_100100110100;
      patterns[51617] = 29'b1_100100110100_001_1_110100100100;
      patterns[51618] = 29'b1_100100110100_010_1_001001101001;
      patterns[51619] = 29'b1_100100110100_011_0_010011010011;
      patterns[51620] = 29'b1_100100110100_100_0_110010011010;
      patterns[51621] = 29'b1_100100110100_101_0_011001001101;
      patterns[51622] = 29'b1_100100110100_110_1_100100110100;
      patterns[51623] = 29'b1_100100110100_111_1_100100110100;
      patterns[51624] = 29'b1_100100110101_000_1_100100110101;
      patterns[51625] = 29'b1_100100110101_001_1_110101100100;
      patterns[51626] = 29'b1_100100110101_010_1_001001101011;
      patterns[51627] = 29'b1_100100110101_011_0_010011010111;
      patterns[51628] = 29'b1_100100110101_100_1_110010011010;
      patterns[51629] = 29'b1_100100110101_101_0_111001001101;
      patterns[51630] = 29'b1_100100110101_110_1_100100110101;
      patterns[51631] = 29'b1_100100110101_111_1_100100110101;
      patterns[51632] = 29'b1_100100110110_000_1_100100110110;
      patterns[51633] = 29'b1_100100110110_001_1_110110100100;
      patterns[51634] = 29'b1_100100110110_010_1_001001101101;
      patterns[51635] = 29'b1_100100110110_011_0_010011011011;
      patterns[51636] = 29'b1_100100110110_100_0_110010011011;
      patterns[51637] = 29'b1_100100110110_101_1_011001001101;
      patterns[51638] = 29'b1_100100110110_110_1_100100110110;
      patterns[51639] = 29'b1_100100110110_111_1_100100110110;
      patterns[51640] = 29'b1_100100110111_000_1_100100110111;
      patterns[51641] = 29'b1_100100110111_001_1_110111100100;
      patterns[51642] = 29'b1_100100110111_010_1_001001101111;
      patterns[51643] = 29'b1_100100110111_011_0_010011011111;
      patterns[51644] = 29'b1_100100110111_100_1_110010011011;
      patterns[51645] = 29'b1_100100110111_101_1_111001001101;
      patterns[51646] = 29'b1_100100110111_110_1_100100110111;
      patterns[51647] = 29'b1_100100110111_111_1_100100110111;
      patterns[51648] = 29'b1_100100111000_000_1_100100111000;
      patterns[51649] = 29'b1_100100111000_001_1_111000100100;
      patterns[51650] = 29'b1_100100111000_010_1_001001110001;
      patterns[51651] = 29'b1_100100111000_011_0_010011100011;
      patterns[51652] = 29'b1_100100111000_100_0_110010011100;
      patterns[51653] = 29'b1_100100111000_101_0_011001001110;
      patterns[51654] = 29'b1_100100111000_110_1_100100111000;
      patterns[51655] = 29'b1_100100111000_111_1_100100111000;
      patterns[51656] = 29'b1_100100111001_000_1_100100111001;
      patterns[51657] = 29'b1_100100111001_001_1_111001100100;
      patterns[51658] = 29'b1_100100111001_010_1_001001110011;
      patterns[51659] = 29'b1_100100111001_011_0_010011100111;
      patterns[51660] = 29'b1_100100111001_100_1_110010011100;
      patterns[51661] = 29'b1_100100111001_101_0_111001001110;
      patterns[51662] = 29'b1_100100111001_110_1_100100111001;
      patterns[51663] = 29'b1_100100111001_111_1_100100111001;
      patterns[51664] = 29'b1_100100111010_000_1_100100111010;
      patterns[51665] = 29'b1_100100111010_001_1_111010100100;
      patterns[51666] = 29'b1_100100111010_010_1_001001110101;
      patterns[51667] = 29'b1_100100111010_011_0_010011101011;
      patterns[51668] = 29'b1_100100111010_100_0_110010011101;
      patterns[51669] = 29'b1_100100111010_101_1_011001001110;
      patterns[51670] = 29'b1_100100111010_110_1_100100111010;
      patterns[51671] = 29'b1_100100111010_111_1_100100111010;
      patterns[51672] = 29'b1_100100111011_000_1_100100111011;
      patterns[51673] = 29'b1_100100111011_001_1_111011100100;
      patterns[51674] = 29'b1_100100111011_010_1_001001110111;
      patterns[51675] = 29'b1_100100111011_011_0_010011101111;
      patterns[51676] = 29'b1_100100111011_100_1_110010011101;
      patterns[51677] = 29'b1_100100111011_101_1_111001001110;
      patterns[51678] = 29'b1_100100111011_110_1_100100111011;
      patterns[51679] = 29'b1_100100111011_111_1_100100111011;
      patterns[51680] = 29'b1_100100111100_000_1_100100111100;
      patterns[51681] = 29'b1_100100111100_001_1_111100100100;
      patterns[51682] = 29'b1_100100111100_010_1_001001111001;
      patterns[51683] = 29'b1_100100111100_011_0_010011110011;
      patterns[51684] = 29'b1_100100111100_100_0_110010011110;
      patterns[51685] = 29'b1_100100111100_101_0_011001001111;
      patterns[51686] = 29'b1_100100111100_110_1_100100111100;
      patterns[51687] = 29'b1_100100111100_111_1_100100111100;
      patterns[51688] = 29'b1_100100111101_000_1_100100111101;
      patterns[51689] = 29'b1_100100111101_001_1_111101100100;
      patterns[51690] = 29'b1_100100111101_010_1_001001111011;
      patterns[51691] = 29'b1_100100111101_011_0_010011110111;
      patterns[51692] = 29'b1_100100111101_100_1_110010011110;
      patterns[51693] = 29'b1_100100111101_101_0_111001001111;
      patterns[51694] = 29'b1_100100111101_110_1_100100111101;
      patterns[51695] = 29'b1_100100111101_111_1_100100111101;
      patterns[51696] = 29'b1_100100111110_000_1_100100111110;
      patterns[51697] = 29'b1_100100111110_001_1_111110100100;
      patterns[51698] = 29'b1_100100111110_010_1_001001111101;
      patterns[51699] = 29'b1_100100111110_011_0_010011111011;
      patterns[51700] = 29'b1_100100111110_100_0_110010011111;
      patterns[51701] = 29'b1_100100111110_101_1_011001001111;
      patterns[51702] = 29'b1_100100111110_110_1_100100111110;
      patterns[51703] = 29'b1_100100111110_111_1_100100111110;
      patterns[51704] = 29'b1_100100111111_000_1_100100111111;
      patterns[51705] = 29'b1_100100111111_001_1_111111100100;
      patterns[51706] = 29'b1_100100111111_010_1_001001111111;
      patterns[51707] = 29'b1_100100111111_011_0_010011111111;
      patterns[51708] = 29'b1_100100111111_100_1_110010011111;
      patterns[51709] = 29'b1_100100111111_101_1_111001001111;
      patterns[51710] = 29'b1_100100111111_110_1_100100111111;
      patterns[51711] = 29'b1_100100111111_111_1_100100111111;
      patterns[51712] = 29'b1_100101000000_000_1_100101000000;
      patterns[51713] = 29'b1_100101000000_001_1_000000100101;
      patterns[51714] = 29'b1_100101000000_010_1_001010000001;
      patterns[51715] = 29'b1_100101000000_011_0_010100000011;
      patterns[51716] = 29'b1_100101000000_100_0_110010100000;
      patterns[51717] = 29'b1_100101000000_101_0_011001010000;
      patterns[51718] = 29'b1_100101000000_110_1_100101000000;
      patterns[51719] = 29'b1_100101000000_111_1_100101000000;
      patterns[51720] = 29'b1_100101000001_000_1_100101000001;
      patterns[51721] = 29'b1_100101000001_001_1_000001100101;
      patterns[51722] = 29'b1_100101000001_010_1_001010000011;
      patterns[51723] = 29'b1_100101000001_011_0_010100000111;
      patterns[51724] = 29'b1_100101000001_100_1_110010100000;
      patterns[51725] = 29'b1_100101000001_101_0_111001010000;
      patterns[51726] = 29'b1_100101000001_110_1_100101000001;
      patterns[51727] = 29'b1_100101000001_111_1_100101000001;
      patterns[51728] = 29'b1_100101000010_000_1_100101000010;
      patterns[51729] = 29'b1_100101000010_001_1_000010100101;
      patterns[51730] = 29'b1_100101000010_010_1_001010000101;
      patterns[51731] = 29'b1_100101000010_011_0_010100001011;
      patterns[51732] = 29'b1_100101000010_100_0_110010100001;
      patterns[51733] = 29'b1_100101000010_101_1_011001010000;
      patterns[51734] = 29'b1_100101000010_110_1_100101000010;
      patterns[51735] = 29'b1_100101000010_111_1_100101000010;
      patterns[51736] = 29'b1_100101000011_000_1_100101000011;
      patterns[51737] = 29'b1_100101000011_001_1_000011100101;
      patterns[51738] = 29'b1_100101000011_010_1_001010000111;
      patterns[51739] = 29'b1_100101000011_011_0_010100001111;
      patterns[51740] = 29'b1_100101000011_100_1_110010100001;
      patterns[51741] = 29'b1_100101000011_101_1_111001010000;
      patterns[51742] = 29'b1_100101000011_110_1_100101000011;
      patterns[51743] = 29'b1_100101000011_111_1_100101000011;
      patterns[51744] = 29'b1_100101000100_000_1_100101000100;
      patterns[51745] = 29'b1_100101000100_001_1_000100100101;
      patterns[51746] = 29'b1_100101000100_010_1_001010001001;
      patterns[51747] = 29'b1_100101000100_011_0_010100010011;
      patterns[51748] = 29'b1_100101000100_100_0_110010100010;
      patterns[51749] = 29'b1_100101000100_101_0_011001010001;
      patterns[51750] = 29'b1_100101000100_110_1_100101000100;
      patterns[51751] = 29'b1_100101000100_111_1_100101000100;
      patterns[51752] = 29'b1_100101000101_000_1_100101000101;
      patterns[51753] = 29'b1_100101000101_001_1_000101100101;
      patterns[51754] = 29'b1_100101000101_010_1_001010001011;
      patterns[51755] = 29'b1_100101000101_011_0_010100010111;
      patterns[51756] = 29'b1_100101000101_100_1_110010100010;
      patterns[51757] = 29'b1_100101000101_101_0_111001010001;
      patterns[51758] = 29'b1_100101000101_110_1_100101000101;
      patterns[51759] = 29'b1_100101000101_111_1_100101000101;
      patterns[51760] = 29'b1_100101000110_000_1_100101000110;
      patterns[51761] = 29'b1_100101000110_001_1_000110100101;
      patterns[51762] = 29'b1_100101000110_010_1_001010001101;
      patterns[51763] = 29'b1_100101000110_011_0_010100011011;
      patterns[51764] = 29'b1_100101000110_100_0_110010100011;
      patterns[51765] = 29'b1_100101000110_101_1_011001010001;
      patterns[51766] = 29'b1_100101000110_110_1_100101000110;
      patterns[51767] = 29'b1_100101000110_111_1_100101000110;
      patterns[51768] = 29'b1_100101000111_000_1_100101000111;
      patterns[51769] = 29'b1_100101000111_001_1_000111100101;
      patterns[51770] = 29'b1_100101000111_010_1_001010001111;
      patterns[51771] = 29'b1_100101000111_011_0_010100011111;
      patterns[51772] = 29'b1_100101000111_100_1_110010100011;
      patterns[51773] = 29'b1_100101000111_101_1_111001010001;
      patterns[51774] = 29'b1_100101000111_110_1_100101000111;
      patterns[51775] = 29'b1_100101000111_111_1_100101000111;
      patterns[51776] = 29'b1_100101001000_000_1_100101001000;
      patterns[51777] = 29'b1_100101001000_001_1_001000100101;
      patterns[51778] = 29'b1_100101001000_010_1_001010010001;
      patterns[51779] = 29'b1_100101001000_011_0_010100100011;
      patterns[51780] = 29'b1_100101001000_100_0_110010100100;
      patterns[51781] = 29'b1_100101001000_101_0_011001010010;
      patterns[51782] = 29'b1_100101001000_110_1_100101001000;
      patterns[51783] = 29'b1_100101001000_111_1_100101001000;
      patterns[51784] = 29'b1_100101001001_000_1_100101001001;
      patterns[51785] = 29'b1_100101001001_001_1_001001100101;
      patterns[51786] = 29'b1_100101001001_010_1_001010010011;
      patterns[51787] = 29'b1_100101001001_011_0_010100100111;
      patterns[51788] = 29'b1_100101001001_100_1_110010100100;
      patterns[51789] = 29'b1_100101001001_101_0_111001010010;
      patterns[51790] = 29'b1_100101001001_110_1_100101001001;
      patterns[51791] = 29'b1_100101001001_111_1_100101001001;
      patterns[51792] = 29'b1_100101001010_000_1_100101001010;
      patterns[51793] = 29'b1_100101001010_001_1_001010100101;
      patterns[51794] = 29'b1_100101001010_010_1_001010010101;
      patterns[51795] = 29'b1_100101001010_011_0_010100101011;
      patterns[51796] = 29'b1_100101001010_100_0_110010100101;
      patterns[51797] = 29'b1_100101001010_101_1_011001010010;
      patterns[51798] = 29'b1_100101001010_110_1_100101001010;
      patterns[51799] = 29'b1_100101001010_111_1_100101001010;
      patterns[51800] = 29'b1_100101001011_000_1_100101001011;
      patterns[51801] = 29'b1_100101001011_001_1_001011100101;
      patterns[51802] = 29'b1_100101001011_010_1_001010010111;
      patterns[51803] = 29'b1_100101001011_011_0_010100101111;
      patterns[51804] = 29'b1_100101001011_100_1_110010100101;
      patterns[51805] = 29'b1_100101001011_101_1_111001010010;
      patterns[51806] = 29'b1_100101001011_110_1_100101001011;
      patterns[51807] = 29'b1_100101001011_111_1_100101001011;
      patterns[51808] = 29'b1_100101001100_000_1_100101001100;
      patterns[51809] = 29'b1_100101001100_001_1_001100100101;
      patterns[51810] = 29'b1_100101001100_010_1_001010011001;
      patterns[51811] = 29'b1_100101001100_011_0_010100110011;
      patterns[51812] = 29'b1_100101001100_100_0_110010100110;
      patterns[51813] = 29'b1_100101001100_101_0_011001010011;
      patterns[51814] = 29'b1_100101001100_110_1_100101001100;
      patterns[51815] = 29'b1_100101001100_111_1_100101001100;
      patterns[51816] = 29'b1_100101001101_000_1_100101001101;
      patterns[51817] = 29'b1_100101001101_001_1_001101100101;
      patterns[51818] = 29'b1_100101001101_010_1_001010011011;
      patterns[51819] = 29'b1_100101001101_011_0_010100110111;
      patterns[51820] = 29'b1_100101001101_100_1_110010100110;
      patterns[51821] = 29'b1_100101001101_101_0_111001010011;
      patterns[51822] = 29'b1_100101001101_110_1_100101001101;
      patterns[51823] = 29'b1_100101001101_111_1_100101001101;
      patterns[51824] = 29'b1_100101001110_000_1_100101001110;
      patterns[51825] = 29'b1_100101001110_001_1_001110100101;
      patterns[51826] = 29'b1_100101001110_010_1_001010011101;
      patterns[51827] = 29'b1_100101001110_011_0_010100111011;
      patterns[51828] = 29'b1_100101001110_100_0_110010100111;
      patterns[51829] = 29'b1_100101001110_101_1_011001010011;
      patterns[51830] = 29'b1_100101001110_110_1_100101001110;
      patterns[51831] = 29'b1_100101001110_111_1_100101001110;
      patterns[51832] = 29'b1_100101001111_000_1_100101001111;
      patterns[51833] = 29'b1_100101001111_001_1_001111100101;
      patterns[51834] = 29'b1_100101001111_010_1_001010011111;
      patterns[51835] = 29'b1_100101001111_011_0_010100111111;
      patterns[51836] = 29'b1_100101001111_100_1_110010100111;
      patterns[51837] = 29'b1_100101001111_101_1_111001010011;
      patterns[51838] = 29'b1_100101001111_110_1_100101001111;
      patterns[51839] = 29'b1_100101001111_111_1_100101001111;
      patterns[51840] = 29'b1_100101010000_000_1_100101010000;
      patterns[51841] = 29'b1_100101010000_001_1_010000100101;
      patterns[51842] = 29'b1_100101010000_010_1_001010100001;
      patterns[51843] = 29'b1_100101010000_011_0_010101000011;
      patterns[51844] = 29'b1_100101010000_100_0_110010101000;
      patterns[51845] = 29'b1_100101010000_101_0_011001010100;
      patterns[51846] = 29'b1_100101010000_110_1_100101010000;
      patterns[51847] = 29'b1_100101010000_111_1_100101010000;
      patterns[51848] = 29'b1_100101010001_000_1_100101010001;
      patterns[51849] = 29'b1_100101010001_001_1_010001100101;
      patterns[51850] = 29'b1_100101010001_010_1_001010100011;
      patterns[51851] = 29'b1_100101010001_011_0_010101000111;
      patterns[51852] = 29'b1_100101010001_100_1_110010101000;
      patterns[51853] = 29'b1_100101010001_101_0_111001010100;
      patterns[51854] = 29'b1_100101010001_110_1_100101010001;
      patterns[51855] = 29'b1_100101010001_111_1_100101010001;
      patterns[51856] = 29'b1_100101010010_000_1_100101010010;
      patterns[51857] = 29'b1_100101010010_001_1_010010100101;
      patterns[51858] = 29'b1_100101010010_010_1_001010100101;
      patterns[51859] = 29'b1_100101010010_011_0_010101001011;
      patterns[51860] = 29'b1_100101010010_100_0_110010101001;
      patterns[51861] = 29'b1_100101010010_101_1_011001010100;
      patterns[51862] = 29'b1_100101010010_110_1_100101010010;
      patterns[51863] = 29'b1_100101010010_111_1_100101010010;
      patterns[51864] = 29'b1_100101010011_000_1_100101010011;
      patterns[51865] = 29'b1_100101010011_001_1_010011100101;
      patterns[51866] = 29'b1_100101010011_010_1_001010100111;
      patterns[51867] = 29'b1_100101010011_011_0_010101001111;
      patterns[51868] = 29'b1_100101010011_100_1_110010101001;
      patterns[51869] = 29'b1_100101010011_101_1_111001010100;
      patterns[51870] = 29'b1_100101010011_110_1_100101010011;
      patterns[51871] = 29'b1_100101010011_111_1_100101010011;
      patterns[51872] = 29'b1_100101010100_000_1_100101010100;
      patterns[51873] = 29'b1_100101010100_001_1_010100100101;
      patterns[51874] = 29'b1_100101010100_010_1_001010101001;
      patterns[51875] = 29'b1_100101010100_011_0_010101010011;
      patterns[51876] = 29'b1_100101010100_100_0_110010101010;
      patterns[51877] = 29'b1_100101010100_101_0_011001010101;
      patterns[51878] = 29'b1_100101010100_110_1_100101010100;
      patterns[51879] = 29'b1_100101010100_111_1_100101010100;
      patterns[51880] = 29'b1_100101010101_000_1_100101010101;
      patterns[51881] = 29'b1_100101010101_001_1_010101100101;
      patterns[51882] = 29'b1_100101010101_010_1_001010101011;
      patterns[51883] = 29'b1_100101010101_011_0_010101010111;
      patterns[51884] = 29'b1_100101010101_100_1_110010101010;
      patterns[51885] = 29'b1_100101010101_101_0_111001010101;
      patterns[51886] = 29'b1_100101010101_110_1_100101010101;
      patterns[51887] = 29'b1_100101010101_111_1_100101010101;
      patterns[51888] = 29'b1_100101010110_000_1_100101010110;
      patterns[51889] = 29'b1_100101010110_001_1_010110100101;
      patterns[51890] = 29'b1_100101010110_010_1_001010101101;
      patterns[51891] = 29'b1_100101010110_011_0_010101011011;
      patterns[51892] = 29'b1_100101010110_100_0_110010101011;
      patterns[51893] = 29'b1_100101010110_101_1_011001010101;
      patterns[51894] = 29'b1_100101010110_110_1_100101010110;
      patterns[51895] = 29'b1_100101010110_111_1_100101010110;
      patterns[51896] = 29'b1_100101010111_000_1_100101010111;
      patterns[51897] = 29'b1_100101010111_001_1_010111100101;
      patterns[51898] = 29'b1_100101010111_010_1_001010101111;
      patterns[51899] = 29'b1_100101010111_011_0_010101011111;
      patterns[51900] = 29'b1_100101010111_100_1_110010101011;
      patterns[51901] = 29'b1_100101010111_101_1_111001010101;
      patterns[51902] = 29'b1_100101010111_110_1_100101010111;
      patterns[51903] = 29'b1_100101010111_111_1_100101010111;
      patterns[51904] = 29'b1_100101011000_000_1_100101011000;
      patterns[51905] = 29'b1_100101011000_001_1_011000100101;
      patterns[51906] = 29'b1_100101011000_010_1_001010110001;
      patterns[51907] = 29'b1_100101011000_011_0_010101100011;
      patterns[51908] = 29'b1_100101011000_100_0_110010101100;
      patterns[51909] = 29'b1_100101011000_101_0_011001010110;
      patterns[51910] = 29'b1_100101011000_110_1_100101011000;
      patterns[51911] = 29'b1_100101011000_111_1_100101011000;
      patterns[51912] = 29'b1_100101011001_000_1_100101011001;
      patterns[51913] = 29'b1_100101011001_001_1_011001100101;
      patterns[51914] = 29'b1_100101011001_010_1_001010110011;
      patterns[51915] = 29'b1_100101011001_011_0_010101100111;
      patterns[51916] = 29'b1_100101011001_100_1_110010101100;
      patterns[51917] = 29'b1_100101011001_101_0_111001010110;
      patterns[51918] = 29'b1_100101011001_110_1_100101011001;
      patterns[51919] = 29'b1_100101011001_111_1_100101011001;
      patterns[51920] = 29'b1_100101011010_000_1_100101011010;
      patterns[51921] = 29'b1_100101011010_001_1_011010100101;
      patterns[51922] = 29'b1_100101011010_010_1_001010110101;
      patterns[51923] = 29'b1_100101011010_011_0_010101101011;
      patterns[51924] = 29'b1_100101011010_100_0_110010101101;
      patterns[51925] = 29'b1_100101011010_101_1_011001010110;
      patterns[51926] = 29'b1_100101011010_110_1_100101011010;
      patterns[51927] = 29'b1_100101011010_111_1_100101011010;
      patterns[51928] = 29'b1_100101011011_000_1_100101011011;
      patterns[51929] = 29'b1_100101011011_001_1_011011100101;
      patterns[51930] = 29'b1_100101011011_010_1_001010110111;
      patterns[51931] = 29'b1_100101011011_011_0_010101101111;
      patterns[51932] = 29'b1_100101011011_100_1_110010101101;
      patterns[51933] = 29'b1_100101011011_101_1_111001010110;
      patterns[51934] = 29'b1_100101011011_110_1_100101011011;
      patterns[51935] = 29'b1_100101011011_111_1_100101011011;
      patterns[51936] = 29'b1_100101011100_000_1_100101011100;
      patterns[51937] = 29'b1_100101011100_001_1_011100100101;
      patterns[51938] = 29'b1_100101011100_010_1_001010111001;
      patterns[51939] = 29'b1_100101011100_011_0_010101110011;
      patterns[51940] = 29'b1_100101011100_100_0_110010101110;
      patterns[51941] = 29'b1_100101011100_101_0_011001010111;
      patterns[51942] = 29'b1_100101011100_110_1_100101011100;
      patterns[51943] = 29'b1_100101011100_111_1_100101011100;
      patterns[51944] = 29'b1_100101011101_000_1_100101011101;
      patterns[51945] = 29'b1_100101011101_001_1_011101100101;
      patterns[51946] = 29'b1_100101011101_010_1_001010111011;
      patterns[51947] = 29'b1_100101011101_011_0_010101110111;
      patterns[51948] = 29'b1_100101011101_100_1_110010101110;
      patterns[51949] = 29'b1_100101011101_101_0_111001010111;
      patterns[51950] = 29'b1_100101011101_110_1_100101011101;
      patterns[51951] = 29'b1_100101011101_111_1_100101011101;
      patterns[51952] = 29'b1_100101011110_000_1_100101011110;
      patterns[51953] = 29'b1_100101011110_001_1_011110100101;
      patterns[51954] = 29'b1_100101011110_010_1_001010111101;
      patterns[51955] = 29'b1_100101011110_011_0_010101111011;
      patterns[51956] = 29'b1_100101011110_100_0_110010101111;
      patterns[51957] = 29'b1_100101011110_101_1_011001010111;
      patterns[51958] = 29'b1_100101011110_110_1_100101011110;
      patterns[51959] = 29'b1_100101011110_111_1_100101011110;
      patterns[51960] = 29'b1_100101011111_000_1_100101011111;
      patterns[51961] = 29'b1_100101011111_001_1_011111100101;
      patterns[51962] = 29'b1_100101011111_010_1_001010111111;
      patterns[51963] = 29'b1_100101011111_011_0_010101111111;
      patterns[51964] = 29'b1_100101011111_100_1_110010101111;
      patterns[51965] = 29'b1_100101011111_101_1_111001010111;
      patterns[51966] = 29'b1_100101011111_110_1_100101011111;
      patterns[51967] = 29'b1_100101011111_111_1_100101011111;
      patterns[51968] = 29'b1_100101100000_000_1_100101100000;
      patterns[51969] = 29'b1_100101100000_001_1_100000100101;
      patterns[51970] = 29'b1_100101100000_010_1_001011000001;
      patterns[51971] = 29'b1_100101100000_011_0_010110000011;
      patterns[51972] = 29'b1_100101100000_100_0_110010110000;
      patterns[51973] = 29'b1_100101100000_101_0_011001011000;
      patterns[51974] = 29'b1_100101100000_110_1_100101100000;
      patterns[51975] = 29'b1_100101100000_111_1_100101100000;
      patterns[51976] = 29'b1_100101100001_000_1_100101100001;
      patterns[51977] = 29'b1_100101100001_001_1_100001100101;
      patterns[51978] = 29'b1_100101100001_010_1_001011000011;
      patterns[51979] = 29'b1_100101100001_011_0_010110000111;
      patterns[51980] = 29'b1_100101100001_100_1_110010110000;
      patterns[51981] = 29'b1_100101100001_101_0_111001011000;
      patterns[51982] = 29'b1_100101100001_110_1_100101100001;
      patterns[51983] = 29'b1_100101100001_111_1_100101100001;
      patterns[51984] = 29'b1_100101100010_000_1_100101100010;
      patterns[51985] = 29'b1_100101100010_001_1_100010100101;
      patterns[51986] = 29'b1_100101100010_010_1_001011000101;
      patterns[51987] = 29'b1_100101100010_011_0_010110001011;
      patterns[51988] = 29'b1_100101100010_100_0_110010110001;
      patterns[51989] = 29'b1_100101100010_101_1_011001011000;
      patterns[51990] = 29'b1_100101100010_110_1_100101100010;
      patterns[51991] = 29'b1_100101100010_111_1_100101100010;
      patterns[51992] = 29'b1_100101100011_000_1_100101100011;
      patterns[51993] = 29'b1_100101100011_001_1_100011100101;
      patterns[51994] = 29'b1_100101100011_010_1_001011000111;
      patterns[51995] = 29'b1_100101100011_011_0_010110001111;
      patterns[51996] = 29'b1_100101100011_100_1_110010110001;
      patterns[51997] = 29'b1_100101100011_101_1_111001011000;
      patterns[51998] = 29'b1_100101100011_110_1_100101100011;
      patterns[51999] = 29'b1_100101100011_111_1_100101100011;
      patterns[52000] = 29'b1_100101100100_000_1_100101100100;
      patterns[52001] = 29'b1_100101100100_001_1_100100100101;
      patterns[52002] = 29'b1_100101100100_010_1_001011001001;
      patterns[52003] = 29'b1_100101100100_011_0_010110010011;
      patterns[52004] = 29'b1_100101100100_100_0_110010110010;
      patterns[52005] = 29'b1_100101100100_101_0_011001011001;
      patterns[52006] = 29'b1_100101100100_110_1_100101100100;
      patterns[52007] = 29'b1_100101100100_111_1_100101100100;
      patterns[52008] = 29'b1_100101100101_000_1_100101100101;
      patterns[52009] = 29'b1_100101100101_001_1_100101100101;
      patterns[52010] = 29'b1_100101100101_010_1_001011001011;
      patterns[52011] = 29'b1_100101100101_011_0_010110010111;
      patterns[52012] = 29'b1_100101100101_100_1_110010110010;
      patterns[52013] = 29'b1_100101100101_101_0_111001011001;
      patterns[52014] = 29'b1_100101100101_110_1_100101100101;
      patterns[52015] = 29'b1_100101100101_111_1_100101100101;
      patterns[52016] = 29'b1_100101100110_000_1_100101100110;
      patterns[52017] = 29'b1_100101100110_001_1_100110100101;
      patterns[52018] = 29'b1_100101100110_010_1_001011001101;
      patterns[52019] = 29'b1_100101100110_011_0_010110011011;
      patterns[52020] = 29'b1_100101100110_100_0_110010110011;
      patterns[52021] = 29'b1_100101100110_101_1_011001011001;
      patterns[52022] = 29'b1_100101100110_110_1_100101100110;
      patterns[52023] = 29'b1_100101100110_111_1_100101100110;
      patterns[52024] = 29'b1_100101100111_000_1_100101100111;
      patterns[52025] = 29'b1_100101100111_001_1_100111100101;
      patterns[52026] = 29'b1_100101100111_010_1_001011001111;
      patterns[52027] = 29'b1_100101100111_011_0_010110011111;
      patterns[52028] = 29'b1_100101100111_100_1_110010110011;
      patterns[52029] = 29'b1_100101100111_101_1_111001011001;
      patterns[52030] = 29'b1_100101100111_110_1_100101100111;
      patterns[52031] = 29'b1_100101100111_111_1_100101100111;
      patterns[52032] = 29'b1_100101101000_000_1_100101101000;
      patterns[52033] = 29'b1_100101101000_001_1_101000100101;
      patterns[52034] = 29'b1_100101101000_010_1_001011010001;
      patterns[52035] = 29'b1_100101101000_011_0_010110100011;
      patterns[52036] = 29'b1_100101101000_100_0_110010110100;
      patterns[52037] = 29'b1_100101101000_101_0_011001011010;
      patterns[52038] = 29'b1_100101101000_110_1_100101101000;
      patterns[52039] = 29'b1_100101101000_111_1_100101101000;
      patterns[52040] = 29'b1_100101101001_000_1_100101101001;
      patterns[52041] = 29'b1_100101101001_001_1_101001100101;
      patterns[52042] = 29'b1_100101101001_010_1_001011010011;
      patterns[52043] = 29'b1_100101101001_011_0_010110100111;
      patterns[52044] = 29'b1_100101101001_100_1_110010110100;
      patterns[52045] = 29'b1_100101101001_101_0_111001011010;
      patterns[52046] = 29'b1_100101101001_110_1_100101101001;
      patterns[52047] = 29'b1_100101101001_111_1_100101101001;
      patterns[52048] = 29'b1_100101101010_000_1_100101101010;
      patterns[52049] = 29'b1_100101101010_001_1_101010100101;
      patterns[52050] = 29'b1_100101101010_010_1_001011010101;
      patterns[52051] = 29'b1_100101101010_011_0_010110101011;
      patterns[52052] = 29'b1_100101101010_100_0_110010110101;
      patterns[52053] = 29'b1_100101101010_101_1_011001011010;
      patterns[52054] = 29'b1_100101101010_110_1_100101101010;
      patterns[52055] = 29'b1_100101101010_111_1_100101101010;
      patterns[52056] = 29'b1_100101101011_000_1_100101101011;
      patterns[52057] = 29'b1_100101101011_001_1_101011100101;
      patterns[52058] = 29'b1_100101101011_010_1_001011010111;
      patterns[52059] = 29'b1_100101101011_011_0_010110101111;
      patterns[52060] = 29'b1_100101101011_100_1_110010110101;
      patterns[52061] = 29'b1_100101101011_101_1_111001011010;
      patterns[52062] = 29'b1_100101101011_110_1_100101101011;
      patterns[52063] = 29'b1_100101101011_111_1_100101101011;
      patterns[52064] = 29'b1_100101101100_000_1_100101101100;
      patterns[52065] = 29'b1_100101101100_001_1_101100100101;
      patterns[52066] = 29'b1_100101101100_010_1_001011011001;
      patterns[52067] = 29'b1_100101101100_011_0_010110110011;
      patterns[52068] = 29'b1_100101101100_100_0_110010110110;
      patterns[52069] = 29'b1_100101101100_101_0_011001011011;
      patterns[52070] = 29'b1_100101101100_110_1_100101101100;
      patterns[52071] = 29'b1_100101101100_111_1_100101101100;
      patterns[52072] = 29'b1_100101101101_000_1_100101101101;
      patterns[52073] = 29'b1_100101101101_001_1_101101100101;
      patterns[52074] = 29'b1_100101101101_010_1_001011011011;
      patterns[52075] = 29'b1_100101101101_011_0_010110110111;
      patterns[52076] = 29'b1_100101101101_100_1_110010110110;
      patterns[52077] = 29'b1_100101101101_101_0_111001011011;
      patterns[52078] = 29'b1_100101101101_110_1_100101101101;
      patterns[52079] = 29'b1_100101101101_111_1_100101101101;
      patterns[52080] = 29'b1_100101101110_000_1_100101101110;
      patterns[52081] = 29'b1_100101101110_001_1_101110100101;
      patterns[52082] = 29'b1_100101101110_010_1_001011011101;
      patterns[52083] = 29'b1_100101101110_011_0_010110111011;
      patterns[52084] = 29'b1_100101101110_100_0_110010110111;
      patterns[52085] = 29'b1_100101101110_101_1_011001011011;
      patterns[52086] = 29'b1_100101101110_110_1_100101101110;
      patterns[52087] = 29'b1_100101101110_111_1_100101101110;
      patterns[52088] = 29'b1_100101101111_000_1_100101101111;
      patterns[52089] = 29'b1_100101101111_001_1_101111100101;
      patterns[52090] = 29'b1_100101101111_010_1_001011011111;
      patterns[52091] = 29'b1_100101101111_011_0_010110111111;
      patterns[52092] = 29'b1_100101101111_100_1_110010110111;
      patterns[52093] = 29'b1_100101101111_101_1_111001011011;
      patterns[52094] = 29'b1_100101101111_110_1_100101101111;
      patterns[52095] = 29'b1_100101101111_111_1_100101101111;
      patterns[52096] = 29'b1_100101110000_000_1_100101110000;
      patterns[52097] = 29'b1_100101110000_001_1_110000100101;
      patterns[52098] = 29'b1_100101110000_010_1_001011100001;
      patterns[52099] = 29'b1_100101110000_011_0_010111000011;
      patterns[52100] = 29'b1_100101110000_100_0_110010111000;
      patterns[52101] = 29'b1_100101110000_101_0_011001011100;
      patterns[52102] = 29'b1_100101110000_110_1_100101110000;
      patterns[52103] = 29'b1_100101110000_111_1_100101110000;
      patterns[52104] = 29'b1_100101110001_000_1_100101110001;
      patterns[52105] = 29'b1_100101110001_001_1_110001100101;
      patterns[52106] = 29'b1_100101110001_010_1_001011100011;
      patterns[52107] = 29'b1_100101110001_011_0_010111000111;
      patterns[52108] = 29'b1_100101110001_100_1_110010111000;
      patterns[52109] = 29'b1_100101110001_101_0_111001011100;
      patterns[52110] = 29'b1_100101110001_110_1_100101110001;
      patterns[52111] = 29'b1_100101110001_111_1_100101110001;
      patterns[52112] = 29'b1_100101110010_000_1_100101110010;
      patterns[52113] = 29'b1_100101110010_001_1_110010100101;
      patterns[52114] = 29'b1_100101110010_010_1_001011100101;
      patterns[52115] = 29'b1_100101110010_011_0_010111001011;
      patterns[52116] = 29'b1_100101110010_100_0_110010111001;
      patterns[52117] = 29'b1_100101110010_101_1_011001011100;
      patterns[52118] = 29'b1_100101110010_110_1_100101110010;
      patterns[52119] = 29'b1_100101110010_111_1_100101110010;
      patterns[52120] = 29'b1_100101110011_000_1_100101110011;
      patterns[52121] = 29'b1_100101110011_001_1_110011100101;
      patterns[52122] = 29'b1_100101110011_010_1_001011100111;
      patterns[52123] = 29'b1_100101110011_011_0_010111001111;
      patterns[52124] = 29'b1_100101110011_100_1_110010111001;
      patterns[52125] = 29'b1_100101110011_101_1_111001011100;
      patterns[52126] = 29'b1_100101110011_110_1_100101110011;
      patterns[52127] = 29'b1_100101110011_111_1_100101110011;
      patterns[52128] = 29'b1_100101110100_000_1_100101110100;
      patterns[52129] = 29'b1_100101110100_001_1_110100100101;
      patterns[52130] = 29'b1_100101110100_010_1_001011101001;
      patterns[52131] = 29'b1_100101110100_011_0_010111010011;
      patterns[52132] = 29'b1_100101110100_100_0_110010111010;
      patterns[52133] = 29'b1_100101110100_101_0_011001011101;
      patterns[52134] = 29'b1_100101110100_110_1_100101110100;
      patterns[52135] = 29'b1_100101110100_111_1_100101110100;
      patterns[52136] = 29'b1_100101110101_000_1_100101110101;
      patterns[52137] = 29'b1_100101110101_001_1_110101100101;
      patterns[52138] = 29'b1_100101110101_010_1_001011101011;
      patterns[52139] = 29'b1_100101110101_011_0_010111010111;
      patterns[52140] = 29'b1_100101110101_100_1_110010111010;
      patterns[52141] = 29'b1_100101110101_101_0_111001011101;
      patterns[52142] = 29'b1_100101110101_110_1_100101110101;
      patterns[52143] = 29'b1_100101110101_111_1_100101110101;
      patterns[52144] = 29'b1_100101110110_000_1_100101110110;
      patterns[52145] = 29'b1_100101110110_001_1_110110100101;
      patterns[52146] = 29'b1_100101110110_010_1_001011101101;
      patterns[52147] = 29'b1_100101110110_011_0_010111011011;
      patterns[52148] = 29'b1_100101110110_100_0_110010111011;
      patterns[52149] = 29'b1_100101110110_101_1_011001011101;
      patterns[52150] = 29'b1_100101110110_110_1_100101110110;
      patterns[52151] = 29'b1_100101110110_111_1_100101110110;
      patterns[52152] = 29'b1_100101110111_000_1_100101110111;
      patterns[52153] = 29'b1_100101110111_001_1_110111100101;
      patterns[52154] = 29'b1_100101110111_010_1_001011101111;
      patterns[52155] = 29'b1_100101110111_011_0_010111011111;
      patterns[52156] = 29'b1_100101110111_100_1_110010111011;
      patterns[52157] = 29'b1_100101110111_101_1_111001011101;
      patterns[52158] = 29'b1_100101110111_110_1_100101110111;
      patterns[52159] = 29'b1_100101110111_111_1_100101110111;
      patterns[52160] = 29'b1_100101111000_000_1_100101111000;
      patterns[52161] = 29'b1_100101111000_001_1_111000100101;
      patterns[52162] = 29'b1_100101111000_010_1_001011110001;
      patterns[52163] = 29'b1_100101111000_011_0_010111100011;
      patterns[52164] = 29'b1_100101111000_100_0_110010111100;
      patterns[52165] = 29'b1_100101111000_101_0_011001011110;
      patterns[52166] = 29'b1_100101111000_110_1_100101111000;
      patterns[52167] = 29'b1_100101111000_111_1_100101111000;
      patterns[52168] = 29'b1_100101111001_000_1_100101111001;
      patterns[52169] = 29'b1_100101111001_001_1_111001100101;
      patterns[52170] = 29'b1_100101111001_010_1_001011110011;
      patterns[52171] = 29'b1_100101111001_011_0_010111100111;
      patterns[52172] = 29'b1_100101111001_100_1_110010111100;
      patterns[52173] = 29'b1_100101111001_101_0_111001011110;
      patterns[52174] = 29'b1_100101111001_110_1_100101111001;
      patterns[52175] = 29'b1_100101111001_111_1_100101111001;
      patterns[52176] = 29'b1_100101111010_000_1_100101111010;
      patterns[52177] = 29'b1_100101111010_001_1_111010100101;
      patterns[52178] = 29'b1_100101111010_010_1_001011110101;
      patterns[52179] = 29'b1_100101111010_011_0_010111101011;
      patterns[52180] = 29'b1_100101111010_100_0_110010111101;
      patterns[52181] = 29'b1_100101111010_101_1_011001011110;
      patterns[52182] = 29'b1_100101111010_110_1_100101111010;
      patterns[52183] = 29'b1_100101111010_111_1_100101111010;
      patterns[52184] = 29'b1_100101111011_000_1_100101111011;
      patterns[52185] = 29'b1_100101111011_001_1_111011100101;
      patterns[52186] = 29'b1_100101111011_010_1_001011110111;
      patterns[52187] = 29'b1_100101111011_011_0_010111101111;
      patterns[52188] = 29'b1_100101111011_100_1_110010111101;
      patterns[52189] = 29'b1_100101111011_101_1_111001011110;
      patterns[52190] = 29'b1_100101111011_110_1_100101111011;
      patterns[52191] = 29'b1_100101111011_111_1_100101111011;
      patterns[52192] = 29'b1_100101111100_000_1_100101111100;
      patterns[52193] = 29'b1_100101111100_001_1_111100100101;
      patterns[52194] = 29'b1_100101111100_010_1_001011111001;
      patterns[52195] = 29'b1_100101111100_011_0_010111110011;
      patterns[52196] = 29'b1_100101111100_100_0_110010111110;
      patterns[52197] = 29'b1_100101111100_101_0_011001011111;
      patterns[52198] = 29'b1_100101111100_110_1_100101111100;
      patterns[52199] = 29'b1_100101111100_111_1_100101111100;
      patterns[52200] = 29'b1_100101111101_000_1_100101111101;
      patterns[52201] = 29'b1_100101111101_001_1_111101100101;
      patterns[52202] = 29'b1_100101111101_010_1_001011111011;
      patterns[52203] = 29'b1_100101111101_011_0_010111110111;
      patterns[52204] = 29'b1_100101111101_100_1_110010111110;
      patterns[52205] = 29'b1_100101111101_101_0_111001011111;
      patterns[52206] = 29'b1_100101111101_110_1_100101111101;
      patterns[52207] = 29'b1_100101111101_111_1_100101111101;
      patterns[52208] = 29'b1_100101111110_000_1_100101111110;
      patterns[52209] = 29'b1_100101111110_001_1_111110100101;
      patterns[52210] = 29'b1_100101111110_010_1_001011111101;
      patterns[52211] = 29'b1_100101111110_011_0_010111111011;
      patterns[52212] = 29'b1_100101111110_100_0_110010111111;
      patterns[52213] = 29'b1_100101111110_101_1_011001011111;
      patterns[52214] = 29'b1_100101111110_110_1_100101111110;
      patterns[52215] = 29'b1_100101111110_111_1_100101111110;
      patterns[52216] = 29'b1_100101111111_000_1_100101111111;
      patterns[52217] = 29'b1_100101111111_001_1_111111100101;
      patterns[52218] = 29'b1_100101111111_010_1_001011111111;
      patterns[52219] = 29'b1_100101111111_011_0_010111111111;
      patterns[52220] = 29'b1_100101111111_100_1_110010111111;
      patterns[52221] = 29'b1_100101111111_101_1_111001011111;
      patterns[52222] = 29'b1_100101111111_110_1_100101111111;
      patterns[52223] = 29'b1_100101111111_111_1_100101111111;
      patterns[52224] = 29'b1_100110000000_000_1_100110000000;
      patterns[52225] = 29'b1_100110000000_001_1_000000100110;
      patterns[52226] = 29'b1_100110000000_010_1_001100000001;
      patterns[52227] = 29'b1_100110000000_011_0_011000000011;
      patterns[52228] = 29'b1_100110000000_100_0_110011000000;
      patterns[52229] = 29'b1_100110000000_101_0_011001100000;
      patterns[52230] = 29'b1_100110000000_110_1_100110000000;
      patterns[52231] = 29'b1_100110000000_111_1_100110000000;
      patterns[52232] = 29'b1_100110000001_000_1_100110000001;
      patterns[52233] = 29'b1_100110000001_001_1_000001100110;
      patterns[52234] = 29'b1_100110000001_010_1_001100000011;
      patterns[52235] = 29'b1_100110000001_011_0_011000000111;
      patterns[52236] = 29'b1_100110000001_100_1_110011000000;
      patterns[52237] = 29'b1_100110000001_101_0_111001100000;
      patterns[52238] = 29'b1_100110000001_110_1_100110000001;
      patterns[52239] = 29'b1_100110000001_111_1_100110000001;
      patterns[52240] = 29'b1_100110000010_000_1_100110000010;
      patterns[52241] = 29'b1_100110000010_001_1_000010100110;
      patterns[52242] = 29'b1_100110000010_010_1_001100000101;
      patterns[52243] = 29'b1_100110000010_011_0_011000001011;
      patterns[52244] = 29'b1_100110000010_100_0_110011000001;
      patterns[52245] = 29'b1_100110000010_101_1_011001100000;
      patterns[52246] = 29'b1_100110000010_110_1_100110000010;
      patterns[52247] = 29'b1_100110000010_111_1_100110000010;
      patterns[52248] = 29'b1_100110000011_000_1_100110000011;
      patterns[52249] = 29'b1_100110000011_001_1_000011100110;
      patterns[52250] = 29'b1_100110000011_010_1_001100000111;
      patterns[52251] = 29'b1_100110000011_011_0_011000001111;
      patterns[52252] = 29'b1_100110000011_100_1_110011000001;
      patterns[52253] = 29'b1_100110000011_101_1_111001100000;
      patterns[52254] = 29'b1_100110000011_110_1_100110000011;
      patterns[52255] = 29'b1_100110000011_111_1_100110000011;
      patterns[52256] = 29'b1_100110000100_000_1_100110000100;
      patterns[52257] = 29'b1_100110000100_001_1_000100100110;
      patterns[52258] = 29'b1_100110000100_010_1_001100001001;
      patterns[52259] = 29'b1_100110000100_011_0_011000010011;
      patterns[52260] = 29'b1_100110000100_100_0_110011000010;
      patterns[52261] = 29'b1_100110000100_101_0_011001100001;
      patterns[52262] = 29'b1_100110000100_110_1_100110000100;
      patterns[52263] = 29'b1_100110000100_111_1_100110000100;
      patterns[52264] = 29'b1_100110000101_000_1_100110000101;
      patterns[52265] = 29'b1_100110000101_001_1_000101100110;
      patterns[52266] = 29'b1_100110000101_010_1_001100001011;
      patterns[52267] = 29'b1_100110000101_011_0_011000010111;
      patterns[52268] = 29'b1_100110000101_100_1_110011000010;
      patterns[52269] = 29'b1_100110000101_101_0_111001100001;
      patterns[52270] = 29'b1_100110000101_110_1_100110000101;
      patterns[52271] = 29'b1_100110000101_111_1_100110000101;
      patterns[52272] = 29'b1_100110000110_000_1_100110000110;
      patterns[52273] = 29'b1_100110000110_001_1_000110100110;
      patterns[52274] = 29'b1_100110000110_010_1_001100001101;
      patterns[52275] = 29'b1_100110000110_011_0_011000011011;
      patterns[52276] = 29'b1_100110000110_100_0_110011000011;
      patterns[52277] = 29'b1_100110000110_101_1_011001100001;
      patterns[52278] = 29'b1_100110000110_110_1_100110000110;
      patterns[52279] = 29'b1_100110000110_111_1_100110000110;
      patterns[52280] = 29'b1_100110000111_000_1_100110000111;
      patterns[52281] = 29'b1_100110000111_001_1_000111100110;
      patterns[52282] = 29'b1_100110000111_010_1_001100001111;
      patterns[52283] = 29'b1_100110000111_011_0_011000011111;
      patterns[52284] = 29'b1_100110000111_100_1_110011000011;
      patterns[52285] = 29'b1_100110000111_101_1_111001100001;
      patterns[52286] = 29'b1_100110000111_110_1_100110000111;
      patterns[52287] = 29'b1_100110000111_111_1_100110000111;
      patterns[52288] = 29'b1_100110001000_000_1_100110001000;
      patterns[52289] = 29'b1_100110001000_001_1_001000100110;
      patterns[52290] = 29'b1_100110001000_010_1_001100010001;
      patterns[52291] = 29'b1_100110001000_011_0_011000100011;
      patterns[52292] = 29'b1_100110001000_100_0_110011000100;
      patterns[52293] = 29'b1_100110001000_101_0_011001100010;
      patterns[52294] = 29'b1_100110001000_110_1_100110001000;
      patterns[52295] = 29'b1_100110001000_111_1_100110001000;
      patterns[52296] = 29'b1_100110001001_000_1_100110001001;
      patterns[52297] = 29'b1_100110001001_001_1_001001100110;
      patterns[52298] = 29'b1_100110001001_010_1_001100010011;
      patterns[52299] = 29'b1_100110001001_011_0_011000100111;
      patterns[52300] = 29'b1_100110001001_100_1_110011000100;
      patterns[52301] = 29'b1_100110001001_101_0_111001100010;
      patterns[52302] = 29'b1_100110001001_110_1_100110001001;
      patterns[52303] = 29'b1_100110001001_111_1_100110001001;
      patterns[52304] = 29'b1_100110001010_000_1_100110001010;
      patterns[52305] = 29'b1_100110001010_001_1_001010100110;
      patterns[52306] = 29'b1_100110001010_010_1_001100010101;
      patterns[52307] = 29'b1_100110001010_011_0_011000101011;
      patterns[52308] = 29'b1_100110001010_100_0_110011000101;
      patterns[52309] = 29'b1_100110001010_101_1_011001100010;
      patterns[52310] = 29'b1_100110001010_110_1_100110001010;
      patterns[52311] = 29'b1_100110001010_111_1_100110001010;
      patterns[52312] = 29'b1_100110001011_000_1_100110001011;
      patterns[52313] = 29'b1_100110001011_001_1_001011100110;
      patterns[52314] = 29'b1_100110001011_010_1_001100010111;
      patterns[52315] = 29'b1_100110001011_011_0_011000101111;
      patterns[52316] = 29'b1_100110001011_100_1_110011000101;
      patterns[52317] = 29'b1_100110001011_101_1_111001100010;
      patterns[52318] = 29'b1_100110001011_110_1_100110001011;
      patterns[52319] = 29'b1_100110001011_111_1_100110001011;
      patterns[52320] = 29'b1_100110001100_000_1_100110001100;
      patterns[52321] = 29'b1_100110001100_001_1_001100100110;
      patterns[52322] = 29'b1_100110001100_010_1_001100011001;
      patterns[52323] = 29'b1_100110001100_011_0_011000110011;
      patterns[52324] = 29'b1_100110001100_100_0_110011000110;
      patterns[52325] = 29'b1_100110001100_101_0_011001100011;
      patterns[52326] = 29'b1_100110001100_110_1_100110001100;
      patterns[52327] = 29'b1_100110001100_111_1_100110001100;
      patterns[52328] = 29'b1_100110001101_000_1_100110001101;
      patterns[52329] = 29'b1_100110001101_001_1_001101100110;
      patterns[52330] = 29'b1_100110001101_010_1_001100011011;
      patterns[52331] = 29'b1_100110001101_011_0_011000110111;
      patterns[52332] = 29'b1_100110001101_100_1_110011000110;
      patterns[52333] = 29'b1_100110001101_101_0_111001100011;
      patterns[52334] = 29'b1_100110001101_110_1_100110001101;
      patterns[52335] = 29'b1_100110001101_111_1_100110001101;
      patterns[52336] = 29'b1_100110001110_000_1_100110001110;
      patterns[52337] = 29'b1_100110001110_001_1_001110100110;
      patterns[52338] = 29'b1_100110001110_010_1_001100011101;
      patterns[52339] = 29'b1_100110001110_011_0_011000111011;
      patterns[52340] = 29'b1_100110001110_100_0_110011000111;
      patterns[52341] = 29'b1_100110001110_101_1_011001100011;
      patterns[52342] = 29'b1_100110001110_110_1_100110001110;
      patterns[52343] = 29'b1_100110001110_111_1_100110001110;
      patterns[52344] = 29'b1_100110001111_000_1_100110001111;
      patterns[52345] = 29'b1_100110001111_001_1_001111100110;
      patterns[52346] = 29'b1_100110001111_010_1_001100011111;
      patterns[52347] = 29'b1_100110001111_011_0_011000111111;
      patterns[52348] = 29'b1_100110001111_100_1_110011000111;
      patterns[52349] = 29'b1_100110001111_101_1_111001100011;
      patterns[52350] = 29'b1_100110001111_110_1_100110001111;
      patterns[52351] = 29'b1_100110001111_111_1_100110001111;
      patterns[52352] = 29'b1_100110010000_000_1_100110010000;
      patterns[52353] = 29'b1_100110010000_001_1_010000100110;
      patterns[52354] = 29'b1_100110010000_010_1_001100100001;
      patterns[52355] = 29'b1_100110010000_011_0_011001000011;
      patterns[52356] = 29'b1_100110010000_100_0_110011001000;
      patterns[52357] = 29'b1_100110010000_101_0_011001100100;
      patterns[52358] = 29'b1_100110010000_110_1_100110010000;
      patterns[52359] = 29'b1_100110010000_111_1_100110010000;
      patterns[52360] = 29'b1_100110010001_000_1_100110010001;
      patterns[52361] = 29'b1_100110010001_001_1_010001100110;
      patterns[52362] = 29'b1_100110010001_010_1_001100100011;
      patterns[52363] = 29'b1_100110010001_011_0_011001000111;
      patterns[52364] = 29'b1_100110010001_100_1_110011001000;
      patterns[52365] = 29'b1_100110010001_101_0_111001100100;
      patterns[52366] = 29'b1_100110010001_110_1_100110010001;
      patterns[52367] = 29'b1_100110010001_111_1_100110010001;
      patterns[52368] = 29'b1_100110010010_000_1_100110010010;
      patterns[52369] = 29'b1_100110010010_001_1_010010100110;
      patterns[52370] = 29'b1_100110010010_010_1_001100100101;
      patterns[52371] = 29'b1_100110010010_011_0_011001001011;
      patterns[52372] = 29'b1_100110010010_100_0_110011001001;
      patterns[52373] = 29'b1_100110010010_101_1_011001100100;
      patterns[52374] = 29'b1_100110010010_110_1_100110010010;
      patterns[52375] = 29'b1_100110010010_111_1_100110010010;
      patterns[52376] = 29'b1_100110010011_000_1_100110010011;
      patterns[52377] = 29'b1_100110010011_001_1_010011100110;
      patterns[52378] = 29'b1_100110010011_010_1_001100100111;
      patterns[52379] = 29'b1_100110010011_011_0_011001001111;
      patterns[52380] = 29'b1_100110010011_100_1_110011001001;
      patterns[52381] = 29'b1_100110010011_101_1_111001100100;
      patterns[52382] = 29'b1_100110010011_110_1_100110010011;
      patterns[52383] = 29'b1_100110010011_111_1_100110010011;
      patterns[52384] = 29'b1_100110010100_000_1_100110010100;
      patterns[52385] = 29'b1_100110010100_001_1_010100100110;
      patterns[52386] = 29'b1_100110010100_010_1_001100101001;
      patterns[52387] = 29'b1_100110010100_011_0_011001010011;
      patterns[52388] = 29'b1_100110010100_100_0_110011001010;
      patterns[52389] = 29'b1_100110010100_101_0_011001100101;
      patterns[52390] = 29'b1_100110010100_110_1_100110010100;
      patterns[52391] = 29'b1_100110010100_111_1_100110010100;
      patterns[52392] = 29'b1_100110010101_000_1_100110010101;
      patterns[52393] = 29'b1_100110010101_001_1_010101100110;
      patterns[52394] = 29'b1_100110010101_010_1_001100101011;
      patterns[52395] = 29'b1_100110010101_011_0_011001010111;
      patterns[52396] = 29'b1_100110010101_100_1_110011001010;
      patterns[52397] = 29'b1_100110010101_101_0_111001100101;
      patterns[52398] = 29'b1_100110010101_110_1_100110010101;
      patterns[52399] = 29'b1_100110010101_111_1_100110010101;
      patterns[52400] = 29'b1_100110010110_000_1_100110010110;
      patterns[52401] = 29'b1_100110010110_001_1_010110100110;
      patterns[52402] = 29'b1_100110010110_010_1_001100101101;
      patterns[52403] = 29'b1_100110010110_011_0_011001011011;
      patterns[52404] = 29'b1_100110010110_100_0_110011001011;
      patterns[52405] = 29'b1_100110010110_101_1_011001100101;
      patterns[52406] = 29'b1_100110010110_110_1_100110010110;
      patterns[52407] = 29'b1_100110010110_111_1_100110010110;
      patterns[52408] = 29'b1_100110010111_000_1_100110010111;
      patterns[52409] = 29'b1_100110010111_001_1_010111100110;
      patterns[52410] = 29'b1_100110010111_010_1_001100101111;
      patterns[52411] = 29'b1_100110010111_011_0_011001011111;
      patterns[52412] = 29'b1_100110010111_100_1_110011001011;
      patterns[52413] = 29'b1_100110010111_101_1_111001100101;
      patterns[52414] = 29'b1_100110010111_110_1_100110010111;
      patterns[52415] = 29'b1_100110010111_111_1_100110010111;
      patterns[52416] = 29'b1_100110011000_000_1_100110011000;
      patterns[52417] = 29'b1_100110011000_001_1_011000100110;
      patterns[52418] = 29'b1_100110011000_010_1_001100110001;
      patterns[52419] = 29'b1_100110011000_011_0_011001100011;
      patterns[52420] = 29'b1_100110011000_100_0_110011001100;
      patterns[52421] = 29'b1_100110011000_101_0_011001100110;
      patterns[52422] = 29'b1_100110011000_110_1_100110011000;
      patterns[52423] = 29'b1_100110011000_111_1_100110011000;
      patterns[52424] = 29'b1_100110011001_000_1_100110011001;
      patterns[52425] = 29'b1_100110011001_001_1_011001100110;
      patterns[52426] = 29'b1_100110011001_010_1_001100110011;
      patterns[52427] = 29'b1_100110011001_011_0_011001100111;
      patterns[52428] = 29'b1_100110011001_100_1_110011001100;
      patterns[52429] = 29'b1_100110011001_101_0_111001100110;
      patterns[52430] = 29'b1_100110011001_110_1_100110011001;
      patterns[52431] = 29'b1_100110011001_111_1_100110011001;
      patterns[52432] = 29'b1_100110011010_000_1_100110011010;
      patterns[52433] = 29'b1_100110011010_001_1_011010100110;
      patterns[52434] = 29'b1_100110011010_010_1_001100110101;
      patterns[52435] = 29'b1_100110011010_011_0_011001101011;
      patterns[52436] = 29'b1_100110011010_100_0_110011001101;
      patterns[52437] = 29'b1_100110011010_101_1_011001100110;
      patterns[52438] = 29'b1_100110011010_110_1_100110011010;
      patterns[52439] = 29'b1_100110011010_111_1_100110011010;
      patterns[52440] = 29'b1_100110011011_000_1_100110011011;
      patterns[52441] = 29'b1_100110011011_001_1_011011100110;
      patterns[52442] = 29'b1_100110011011_010_1_001100110111;
      patterns[52443] = 29'b1_100110011011_011_0_011001101111;
      patterns[52444] = 29'b1_100110011011_100_1_110011001101;
      patterns[52445] = 29'b1_100110011011_101_1_111001100110;
      patterns[52446] = 29'b1_100110011011_110_1_100110011011;
      patterns[52447] = 29'b1_100110011011_111_1_100110011011;
      patterns[52448] = 29'b1_100110011100_000_1_100110011100;
      patterns[52449] = 29'b1_100110011100_001_1_011100100110;
      patterns[52450] = 29'b1_100110011100_010_1_001100111001;
      patterns[52451] = 29'b1_100110011100_011_0_011001110011;
      patterns[52452] = 29'b1_100110011100_100_0_110011001110;
      patterns[52453] = 29'b1_100110011100_101_0_011001100111;
      patterns[52454] = 29'b1_100110011100_110_1_100110011100;
      patterns[52455] = 29'b1_100110011100_111_1_100110011100;
      patterns[52456] = 29'b1_100110011101_000_1_100110011101;
      patterns[52457] = 29'b1_100110011101_001_1_011101100110;
      patterns[52458] = 29'b1_100110011101_010_1_001100111011;
      patterns[52459] = 29'b1_100110011101_011_0_011001110111;
      patterns[52460] = 29'b1_100110011101_100_1_110011001110;
      patterns[52461] = 29'b1_100110011101_101_0_111001100111;
      patterns[52462] = 29'b1_100110011101_110_1_100110011101;
      patterns[52463] = 29'b1_100110011101_111_1_100110011101;
      patterns[52464] = 29'b1_100110011110_000_1_100110011110;
      patterns[52465] = 29'b1_100110011110_001_1_011110100110;
      patterns[52466] = 29'b1_100110011110_010_1_001100111101;
      patterns[52467] = 29'b1_100110011110_011_0_011001111011;
      patterns[52468] = 29'b1_100110011110_100_0_110011001111;
      patterns[52469] = 29'b1_100110011110_101_1_011001100111;
      patterns[52470] = 29'b1_100110011110_110_1_100110011110;
      patterns[52471] = 29'b1_100110011110_111_1_100110011110;
      patterns[52472] = 29'b1_100110011111_000_1_100110011111;
      patterns[52473] = 29'b1_100110011111_001_1_011111100110;
      patterns[52474] = 29'b1_100110011111_010_1_001100111111;
      patterns[52475] = 29'b1_100110011111_011_0_011001111111;
      patterns[52476] = 29'b1_100110011111_100_1_110011001111;
      patterns[52477] = 29'b1_100110011111_101_1_111001100111;
      patterns[52478] = 29'b1_100110011111_110_1_100110011111;
      patterns[52479] = 29'b1_100110011111_111_1_100110011111;
      patterns[52480] = 29'b1_100110100000_000_1_100110100000;
      patterns[52481] = 29'b1_100110100000_001_1_100000100110;
      patterns[52482] = 29'b1_100110100000_010_1_001101000001;
      patterns[52483] = 29'b1_100110100000_011_0_011010000011;
      patterns[52484] = 29'b1_100110100000_100_0_110011010000;
      patterns[52485] = 29'b1_100110100000_101_0_011001101000;
      patterns[52486] = 29'b1_100110100000_110_1_100110100000;
      patterns[52487] = 29'b1_100110100000_111_1_100110100000;
      patterns[52488] = 29'b1_100110100001_000_1_100110100001;
      patterns[52489] = 29'b1_100110100001_001_1_100001100110;
      patterns[52490] = 29'b1_100110100001_010_1_001101000011;
      patterns[52491] = 29'b1_100110100001_011_0_011010000111;
      patterns[52492] = 29'b1_100110100001_100_1_110011010000;
      patterns[52493] = 29'b1_100110100001_101_0_111001101000;
      patterns[52494] = 29'b1_100110100001_110_1_100110100001;
      patterns[52495] = 29'b1_100110100001_111_1_100110100001;
      patterns[52496] = 29'b1_100110100010_000_1_100110100010;
      patterns[52497] = 29'b1_100110100010_001_1_100010100110;
      patterns[52498] = 29'b1_100110100010_010_1_001101000101;
      patterns[52499] = 29'b1_100110100010_011_0_011010001011;
      patterns[52500] = 29'b1_100110100010_100_0_110011010001;
      patterns[52501] = 29'b1_100110100010_101_1_011001101000;
      patterns[52502] = 29'b1_100110100010_110_1_100110100010;
      patterns[52503] = 29'b1_100110100010_111_1_100110100010;
      patterns[52504] = 29'b1_100110100011_000_1_100110100011;
      patterns[52505] = 29'b1_100110100011_001_1_100011100110;
      patterns[52506] = 29'b1_100110100011_010_1_001101000111;
      patterns[52507] = 29'b1_100110100011_011_0_011010001111;
      patterns[52508] = 29'b1_100110100011_100_1_110011010001;
      patterns[52509] = 29'b1_100110100011_101_1_111001101000;
      patterns[52510] = 29'b1_100110100011_110_1_100110100011;
      patterns[52511] = 29'b1_100110100011_111_1_100110100011;
      patterns[52512] = 29'b1_100110100100_000_1_100110100100;
      patterns[52513] = 29'b1_100110100100_001_1_100100100110;
      patterns[52514] = 29'b1_100110100100_010_1_001101001001;
      patterns[52515] = 29'b1_100110100100_011_0_011010010011;
      patterns[52516] = 29'b1_100110100100_100_0_110011010010;
      patterns[52517] = 29'b1_100110100100_101_0_011001101001;
      patterns[52518] = 29'b1_100110100100_110_1_100110100100;
      patterns[52519] = 29'b1_100110100100_111_1_100110100100;
      patterns[52520] = 29'b1_100110100101_000_1_100110100101;
      patterns[52521] = 29'b1_100110100101_001_1_100101100110;
      patterns[52522] = 29'b1_100110100101_010_1_001101001011;
      patterns[52523] = 29'b1_100110100101_011_0_011010010111;
      patterns[52524] = 29'b1_100110100101_100_1_110011010010;
      patterns[52525] = 29'b1_100110100101_101_0_111001101001;
      patterns[52526] = 29'b1_100110100101_110_1_100110100101;
      patterns[52527] = 29'b1_100110100101_111_1_100110100101;
      patterns[52528] = 29'b1_100110100110_000_1_100110100110;
      patterns[52529] = 29'b1_100110100110_001_1_100110100110;
      patterns[52530] = 29'b1_100110100110_010_1_001101001101;
      patterns[52531] = 29'b1_100110100110_011_0_011010011011;
      patterns[52532] = 29'b1_100110100110_100_0_110011010011;
      patterns[52533] = 29'b1_100110100110_101_1_011001101001;
      patterns[52534] = 29'b1_100110100110_110_1_100110100110;
      patterns[52535] = 29'b1_100110100110_111_1_100110100110;
      patterns[52536] = 29'b1_100110100111_000_1_100110100111;
      patterns[52537] = 29'b1_100110100111_001_1_100111100110;
      patterns[52538] = 29'b1_100110100111_010_1_001101001111;
      patterns[52539] = 29'b1_100110100111_011_0_011010011111;
      patterns[52540] = 29'b1_100110100111_100_1_110011010011;
      patterns[52541] = 29'b1_100110100111_101_1_111001101001;
      patterns[52542] = 29'b1_100110100111_110_1_100110100111;
      patterns[52543] = 29'b1_100110100111_111_1_100110100111;
      patterns[52544] = 29'b1_100110101000_000_1_100110101000;
      patterns[52545] = 29'b1_100110101000_001_1_101000100110;
      patterns[52546] = 29'b1_100110101000_010_1_001101010001;
      patterns[52547] = 29'b1_100110101000_011_0_011010100011;
      patterns[52548] = 29'b1_100110101000_100_0_110011010100;
      patterns[52549] = 29'b1_100110101000_101_0_011001101010;
      patterns[52550] = 29'b1_100110101000_110_1_100110101000;
      patterns[52551] = 29'b1_100110101000_111_1_100110101000;
      patterns[52552] = 29'b1_100110101001_000_1_100110101001;
      patterns[52553] = 29'b1_100110101001_001_1_101001100110;
      patterns[52554] = 29'b1_100110101001_010_1_001101010011;
      patterns[52555] = 29'b1_100110101001_011_0_011010100111;
      patterns[52556] = 29'b1_100110101001_100_1_110011010100;
      patterns[52557] = 29'b1_100110101001_101_0_111001101010;
      patterns[52558] = 29'b1_100110101001_110_1_100110101001;
      patterns[52559] = 29'b1_100110101001_111_1_100110101001;
      patterns[52560] = 29'b1_100110101010_000_1_100110101010;
      patterns[52561] = 29'b1_100110101010_001_1_101010100110;
      patterns[52562] = 29'b1_100110101010_010_1_001101010101;
      patterns[52563] = 29'b1_100110101010_011_0_011010101011;
      patterns[52564] = 29'b1_100110101010_100_0_110011010101;
      patterns[52565] = 29'b1_100110101010_101_1_011001101010;
      patterns[52566] = 29'b1_100110101010_110_1_100110101010;
      patterns[52567] = 29'b1_100110101010_111_1_100110101010;
      patterns[52568] = 29'b1_100110101011_000_1_100110101011;
      patterns[52569] = 29'b1_100110101011_001_1_101011100110;
      patterns[52570] = 29'b1_100110101011_010_1_001101010111;
      patterns[52571] = 29'b1_100110101011_011_0_011010101111;
      patterns[52572] = 29'b1_100110101011_100_1_110011010101;
      patterns[52573] = 29'b1_100110101011_101_1_111001101010;
      patterns[52574] = 29'b1_100110101011_110_1_100110101011;
      patterns[52575] = 29'b1_100110101011_111_1_100110101011;
      patterns[52576] = 29'b1_100110101100_000_1_100110101100;
      patterns[52577] = 29'b1_100110101100_001_1_101100100110;
      patterns[52578] = 29'b1_100110101100_010_1_001101011001;
      patterns[52579] = 29'b1_100110101100_011_0_011010110011;
      patterns[52580] = 29'b1_100110101100_100_0_110011010110;
      patterns[52581] = 29'b1_100110101100_101_0_011001101011;
      patterns[52582] = 29'b1_100110101100_110_1_100110101100;
      patterns[52583] = 29'b1_100110101100_111_1_100110101100;
      patterns[52584] = 29'b1_100110101101_000_1_100110101101;
      patterns[52585] = 29'b1_100110101101_001_1_101101100110;
      patterns[52586] = 29'b1_100110101101_010_1_001101011011;
      patterns[52587] = 29'b1_100110101101_011_0_011010110111;
      patterns[52588] = 29'b1_100110101101_100_1_110011010110;
      patterns[52589] = 29'b1_100110101101_101_0_111001101011;
      patterns[52590] = 29'b1_100110101101_110_1_100110101101;
      patterns[52591] = 29'b1_100110101101_111_1_100110101101;
      patterns[52592] = 29'b1_100110101110_000_1_100110101110;
      patterns[52593] = 29'b1_100110101110_001_1_101110100110;
      patterns[52594] = 29'b1_100110101110_010_1_001101011101;
      patterns[52595] = 29'b1_100110101110_011_0_011010111011;
      patterns[52596] = 29'b1_100110101110_100_0_110011010111;
      patterns[52597] = 29'b1_100110101110_101_1_011001101011;
      patterns[52598] = 29'b1_100110101110_110_1_100110101110;
      patterns[52599] = 29'b1_100110101110_111_1_100110101110;
      patterns[52600] = 29'b1_100110101111_000_1_100110101111;
      patterns[52601] = 29'b1_100110101111_001_1_101111100110;
      patterns[52602] = 29'b1_100110101111_010_1_001101011111;
      patterns[52603] = 29'b1_100110101111_011_0_011010111111;
      patterns[52604] = 29'b1_100110101111_100_1_110011010111;
      patterns[52605] = 29'b1_100110101111_101_1_111001101011;
      patterns[52606] = 29'b1_100110101111_110_1_100110101111;
      patterns[52607] = 29'b1_100110101111_111_1_100110101111;
      patterns[52608] = 29'b1_100110110000_000_1_100110110000;
      patterns[52609] = 29'b1_100110110000_001_1_110000100110;
      patterns[52610] = 29'b1_100110110000_010_1_001101100001;
      patterns[52611] = 29'b1_100110110000_011_0_011011000011;
      patterns[52612] = 29'b1_100110110000_100_0_110011011000;
      patterns[52613] = 29'b1_100110110000_101_0_011001101100;
      patterns[52614] = 29'b1_100110110000_110_1_100110110000;
      patterns[52615] = 29'b1_100110110000_111_1_100110110000;
      patterns[52616] = 29'b1_100110110001_000_1_100110110001;
      patterns[52617] = 29'b1_100110110001_001_1_110001100110;
      patterns[52618] = 29'b1_100110110001_010_1_001101100011;
      patterns[52619] = 29'b1_100110110001_011_0_011011000111;
      patterns[52620] = 29'b1_100110110001_100_1_110011011000;
      patterns[52621] = 29'b1_100110110001_101_0_111001101100;
      patterns[52622] = 29'b1_100110110001_110_1_100110110001;
      patterns[52623] = 29'b1_100110110001_111_1_100110110001;
      patterns[52624] = 29'b1_100110110010_000_1_100110110010;
      patterns[52625] = 29'b1_100110110010_001_1_110010100110;
      patterns[52626] = 29'b1_100110110010_010_1_001101100101;
      patterns[52627] = 29'b1_100110110010_011_0_011011001011;
      patterns[52628] = 29'b1_100110110010_100_0_110011011001;
      patterns[52629] = 29'b1_100110110010_101_1_011001101100;
      patterns[52630] = 29'b1_100110110010_110_1_100110110010;
      patterns[52631] = 29'b1_100110110010_111_1_100110110010;
      patterns[52632] = 29'b1_100110110011_000_1_100110110011;
      patterns[52633] = 29'b1_100110110011_001_1_110011100110;
      patterns[52634] = 29'b1_100110110011_010_1_001101100111;
      patterns[52635] = 29'b1_100110110011_011_0_011011001111;
      patterns[52636] = 29'b1_100110110011_100_1_110011011001;
      patterns[52637] = 29'b1_100110110011_101_1_111001101100;
      patterns[52638] = 29'b1_100110110011_110_1_100110110011;
      patterns[52639] = 29'b1_100110110011_111_1_100110110011;
      patterns[52640] = 29'b1_100110110100_000_1_100110110100;
      patterns[52641] = 29'b1_100110110100_001_1_110100100110;
      patterns[52642] = 29'b1_100110110100_010_1_001101101001;
      patterns[52643] = 29'b1_100110110100_011_0_011011010011;
      patterns[52644] = 29'b1_100110110100_100_0_110011011010;
      patterns[52645] = 29'b1_100110110100_101_0_011001101101;
      patterns[52646] = 29'b1_100110110100_110_1_100110110100;
      patterns[52647] = 29'b1_100110110100_111_1_100110110100;
      patterns[52648] = 29'b1_100110110101_000_1_100110110101;
      patterns[52649] = 29'b1_100110110101_001_1_110101100110;
      patterns[52650] = 29'b1_100110110101_010_1_001101101011;
      patterns[52651] = 29'b1_100110110101_011_0_011011010111;
      patterns[52652] = 29'b1_100110110101_100_1_110011011010;
      patterns[52653] = 29'b1_100110110101_101_0_111001101101;
      patterns[52654] = 29'b1_100110110101_110_1_100110110101;
      patterns[52655] = 29'b1_100110110101_111_1_100110110101;
      patterns[52656] = 29'b1_100110110110_000_1_100110110110;
      patterns[52657] = 29'b1_100110110110_001_1_110110100110;
      patterns[52658] = 29'b1_100110110110_010_1_001101101101;
      patterns[52659] = 29'b1_100110110110_011_0_011011011011;
      patterns[52660] = 29'b1_100110110110_100_0_110011011011;
      patterns[52661] = 29'b1_100110110110_101_1_011001101101;
      patterns[52662] = 29'b1_100110110110_110_1_100110110110;
      patterns[52663] = 29'b1_100110110110_111_1_100110110110;
      patterns[52664] = 29'b1_100110110111_000_1_100110110111;
      patterns[52665] = 29'b1_100110110111_001_1_110111100110;
      patterns[52666] = 29'b1_100110110111_010_1_001101101111;
      patterns[52667] = 29'b1_100110110111_011_0_011011011111;
      patterns[52668] = 29'b1_100110110111_100_1_110011011011;
      patterns[52669] = 29'b1_100110110111_101_1_111001101101;
      patterns[52670] = 29'b1_100110110111_110_1_100110110111;
      patterns[52671] = 29'b1_100110110111_111_1_100110110111;
      patterns[52672] = 29'b1_100110111000_000_1_100110111000;
      patterns[52673] = 29'b1_100110111000_001_1_111000100110;
      patterns[52674] = 29'b1_100110111000_010_1_001101110001;
      patterns[52675] = 29'b1_100110111000_011_0_011011100011;
      patterns[52676] = 29'b1_100110111000_100_0_110011011100;
      patterns[52677] = 29'b1_100110111000_101_0_011001101110;
      patterns[52678] = 29'b1_100110111000_110_1_100110111000;
      patterns[52679] = 29'b1_100110111000_111_1_100110111000;
      patterns[52680] = 29'b1_100110111001_000_1_100110111001;
      patterns[52681] = 29'b1_100110111001_001_1_111001100110;
      patterns[52682] = 29'b1_100110111001_010_1_001101110011;
      patterns[52683] = 29'b1_100110111001_011_0_011011100111;
      patterns[52684] = 29'b1_100110111001_100_1_110011011100;
      patterns[52685] = 29'b1_100110111001_101_0_111001101110;
      patterns[52686] = 29'b1_100110111001_110_1_100110111001;
      patterns[52687] = 29'b1_100110111001_111_1_100110111001;
      patterns[52688] = 29'b1_100110111010_000_1_100110111010;
      patterns[52689] = 29'b1_100110111010_001_1_111010100110;
      patterns[52690] = 29'b1_100110111010_010_1_001101110101;
      patterns[52691] = 29'b1_100110111010_011_0_011011101011;
      patterns[52692] = 29'b1_100110111010_100_0_110011011101;
      patterns[52693] = 29'b1_100110111010_101_1_011001101110;
      patterns[52694] = 29'b1_100110111010_110_1_100110111010;
      patterns[52695] = 29'b1_100110111010_111_1_100110111010;
      patterns[52696] = 29'b1_100110111011_000_1_100110111011;
      patterns[52697] = 29'b1_100110111011_001_1_111011100110;
      patterns[52698] = 29'b1_100110111011_010_1_001101110111;
      patterns[52699] = 29'b1_100110111011_011_0_011011101111;
      patterns[52700] = 29'b1_100110111011_100_1_110011011101;
      patterns[52701] = 29'b1_100110111011_101_1_111001101110;
      patterns[52702] = 29'b1_100110111011_110_1_100110111011;
      patterns[52703] = 29'b1_100110111011_111_1_100110111011;
      patterns[52704] = 29'b1_100110111100_000_1_100110111100;
      patterns[52705] = 29'b1_100110111100_001_1_111100100110;
      patterns[52706] = 29'b1_100110111100_010_1_001101111001;
      patterns[52707] = 29'b1_100110111100_011_0_011011110011;
      patterns[52708] = 29'b1_100110111100_100_0_110011011110;
      patterns[52709] = 29'b1_100110111100_101_0_011001101111;
      patterns[52710] = 29'b1_100110111100_110_1_100110111100;
      patterns[52711] = 29'b1_100110111100_111_1_100110111100;
      patterns[52712] = 29'b1_100110111101_000_1_100110111101;
      patterns[52713] = 29'b1_100110111101_001_1_111101100110;
      patterns[52714] = 29'b1_100110111101_010_1_001101111011;
      patterns[52715] = 29'b1_100110111101_011_0_011011110111;
      patterns[52716] = 29'b1_100110111101_100_1_110011011110;
      patterns[52717] = 29'b1_100110111101_101_0_111001101111;
      patterns[52718] = 29'b1_100110111101_110_1_100110111101;
      patterns[52719] = 29'b1_100110111101_111_1_100110111101;
      patterns[52720] = 29'b1_100110111110_000_1_100110111110;
      patterns[52721] = 29'b1_100110111110_001_1_111110100110;
      patterns[52722] = 29'b1_100110111110_010_1_001101111101;
      patterns[52723] = 29'b1_100110111110_011_0_011011111011;
      patterns[52724] = 29'b1_100110111110_100_0_110011011111;
      patterns[52725] = 29'b1_100110111110_101_1_011001101111;
      patterns[52726] = 29'b1_100110111110_110_1_100110111110;
      patterns[52727] = 29'b1_100110111110_111_1_100110111110;
      patterns[52728] = 29'b1_100110111111_000_1_100110111111;
      patterns[52729] = 29'b1_100110111111_001_1_111111100110;
      patterns[52730] = 29'b1_100110111111_010_1_001101111111;
      patterns[52731] = 29'b1_100110111111_011_0_011011111111;
      patterns[52732] = 29'b1_100110111111_100_1_110011011111;
      patterns[52733] = 29'b1_100110111111_101_1_111001101111;
      patterns[52734] = 29'b1_100110111111_110_1_100110111111;
      patterns[52735] = 29'b1_100110111111_111_1_100110111111;
      patterns[52736] = 29'b1_100111000000_000_1_100111000000;
      patterns[52737] = 29'b1_100111000000_001_1_000000100111;
      patterns[52738] = 29'b1_100111000000_010_1_001110000001;
      patterns[52739] = 29'b1_100111000000_011_0_011100000011;
      patterns[52740] = 29'b1_100111000000_100_0_110011100000;
      patterns[52741] = 29'b1_100111000000_101_0_011001110000;
      patterns[52742] = 29'b1_100111000000_110_1_100111000000;
      patterns[52743] = 29'b1_100111000000_111_1_100111000000;
      patterns[52744] = 29'b1_100111000001_000_1_100111000001;
      patterns[52745] = 29'b1_100111000001_001_1_000001100111;
      patterns[52746] = 29'b1_100111000001_010_1_001110000011;
      patterns[52747] = 29'b1_100111000001_011_0_011100000111;
      patterns[52748] = 29'b1_100111000001_100_1_110011100000;
      patterns[52749] = 29'b1_100111000001_101_0_111001110000;
      patterns[52750] = 29'b1_100111000001_110_1_100111000001;
      patterns[52751] = 29'b1_100111000001_111_1_100111000001;
      patterns[52752] = 29'b1_100111000010_000_1_100111000010;
      patterns[52753] = 29'b1_100111000010_001_1_000010100111;
      patterns[52754] = 29'b1_100111000010_010_1_001110000101;
      patterns[52755] = 29'b1_100111000010_011_0_011100001011;
      patterns[52756] = 29'b1_100111000010_100_0_110011100001;
      patterns[52757] = 29'b1_100111000010_101_1_011001110000;
      patterns[52758] = 29'b1_100111000010_110_1_100111000010;
      patterns[52759] = 29'b1_100111000010_111_1_100111000010;
      patterns[52760] = 29'b1_100111000011_000_1_100111000011;
      patterns[52761] = 29'b1_100111000011_001_1_000011100111;
      patterns[52762] = 29'b1_100111000011_010_1_001110000111;
      patterns[52763] = 29'b1_100111000011_011_0_011100001111;
      patterns[52764] = 29'b1_100111000011_100_1_110011100001;
      patterns[52765] = 29'b1_100111000011_101_1_111001110000;
      patterns[52766] = 29'b1_100111000011_110_1_100111000011;
      patterns[52767] = 29'b1_100111000011_111_1_100111000011;
      patterns[52768] = 29'b1_100111000100_000_1_100111000100;
      patterns[52769] = 29'b1_100111000100_001_1_000100100111;
      patterns[52770] = 29'b1_100111000100_010_1_001110001001;
      patterns[52771] = 29'b1_100111000100_011_0_011100010011;
      patterns[52772] = 29'b1_100111000100_100_0_110011100010;
      patterns[52773] = 29'b1_100111000100_101_0_011001110001;
      patterns[52774] = 29'b1_100111000100_110_1_100111000100;
      patterns[52775] = 29'b1_100111000100_111_1_100111000100;
      patterns[52776] = 29'b1_100111000101_000_1_100111000101;
      patterns[52777] = 29'b1_100111000101_001_1_000101100111;
      patterns[52778] = 29'b1_100111000101_010_1_001110001011;
      patterns[52779] = 29'b1_100111000101_011_0_011100010111;
      patterns[52780] = 29'b1_100111000101_100_1_110011100010;
      patterns[52781] = 29'b1_100111000101_101_0_111001110001;
      patterns[52782] = 29'b1_100111000101_110_1_100111000101;
      patterns[52783] = 29'b1_100111000101_111_1_100111000101;
      patterns[52784] = 29'b1_100111000110_000_1_100111000110;
      patterns[52785] = 29'b1_100111000110_001_1_000110100111;
      patterns[52786] = 29'b1_100111000110_010_1_001110001101;
      patterns[52787] = 29'b1_100111000110_011_0_011100011011;
      patterns[52788] = 29'b1_100111000110_100_0_110011100011;
      patterns[52789] = 29'b1_100111000110_101_1_011001110001;
      patterns[52790] = 29'b1_100111000110_110_1_100111000110;
      patterns[52791] = 29'b1_100111000110_111_1_100111000110;
      patterns[52792] = 29'b1_100111000111_000_1_100111000111;
      patterns[52793] = 29'b1_100111000111_001_1_000111100111;
      patterns[52794] = 29'b1_100111000111_010_1_001110001111;
      patterns[52795] = 29'b1_100111000111_011_0_011100011111;
      patterns[52796] = 29'b1_100111000111_100_1_110011100011;
      patterns[52797] = 29'b1_100111000111_101_1_111001110001;
      patterns[52798] = 29'b1_100111000111_110_1_100111000111;
      patterns[52799] = 29'b1_100111000111_111_1_100111000111;
      patterns[52800] = 29'b1_100111001000_000_1_100111001000;
      patterns[52801] = 29'b1_100111001000_001_1_001000100111;
      patterns[52802] = 29'b1_100111001000_010_1_001110010001;
      patterns[52803] = 29'b1_100111001000_011_0_011100100011;
      patterns[52804] = 29'b1_100111001000_100_0_110011100100;
      patterns[52805] = 29'b1_100111001000_101_0_011001110010;
      patterns[52806] = 29'b1_100111001000_110_1_100111001000;
      patterns[52807] = 29'b1_100111001000_111_1_100111001000;
      patterns[52808] = 29'b1_100111001001_000_1_100111001001;
      patterns[52809] = 29'b1_100111001001_001_1_001001100111;
      patterns[52810] = 29'b1_100111001001_010_1_001110010011;
      patterns[52811] = 29'b1_100111001001_011_0_011100100111;
      patterns[52812] = 29'b1_100111001001_100_1_110011100100;
      patterns[52813] = 29'b1_100111001001_101_0_111001110010;
      patterns[52814] = 29'b1_100111001001_110_1_100111001001;
      patterns[52815] = 29'b1_100111001001_111_1_100111001001;
      patterns[52816] = 29'b1_100111001010_000_1_100111001010;
      patterns[52817] = 29'b1_100111001010_001_1_001010100111;
      patterns[52818] = 29'b1_100111001010_010_1_001110010101;
      patterns[52819] = 29'b1_100111001010_011_0_011100101011;
      patterns[52820] = 29'b1_100111001010_100_0_110011100101;
      patterns[52821] = 29'b1_100111001010_101_1_011001110010;
      patterns[52822] = 29'b1_100111001010_110_1_100111001010;
      patterns[52823] = 29'b1_100111001010_111_1_100111001010;
      patterns[52824] = 29'b1_100111001011_000_1_100111001011;
      patterns[52825] = 29'b1_100111001011_001_1_001011100111;
      patterns[52826] = 29'b1_100111001011_010_1_001110010111;
      patterns[52827] = 29'b1_100111001011_011_0_011100101111;
      patterns[52828] = 29'b1_100111001011_100_1_110011100101;
      patterns[52829] = 29'b1_100111001011_101_1_111001110010;
      patterns[52830] = 29'b1_100111001011_110_1_100111001011;
      patterns[52831] = 29'b1_100111001011_111_1_100111001011;
      patterns[52832] = 29'b1_100111001100_000_1_100111001100;
      patterns[52833] = 29'b1_100111001100_001_1_001100100111;
      patterns[52834] = 29'b1_100111001100_010_1_001110011001;
      patterns[52835] = 29'b1_100111001100_011_0_011100110011;
      patterns[52836] = 29'b1_100111001100_100_0_110011100110;
      patterns[52837] = 29'b1_100111001100_101_0_011001110011;
      patterns[52838] = 29'b1_100111001100_110_1_100111001100;
      patterns[52839] = 29'b1_100111001100_111_1_100111001100;
      patterns[52840] = 29'b1_100111001101_000_1_100111001101;
      patterns[52841] = 29'b1_100111001101_001_1_001101100111;
      patterns[52842] = 29'b1_100111001101_010_1_001110011011;
      patterns[52843] = 29'b1_100111001101_011_0_011100110111;
      patterns[52844] = 29'b1_100111001101_100_1_110011100110;
      patterns[52845] = 29'b1_100111001101_101_0_111001110011;
      patterns[52846] = 29'b1_100111001101_110_1_100111001101;
      patterns[52847] = 29'b1_100111001101_111_1_100111001101;
      patterns[52848] = 29'b1_100111001110_000_1_100111001110;
      patterns[52849] = 29'b1_100111001110_001_1_001110100111;
      patterns[52850] = 29'b1_100111001110_010_1_001110011101;
      patterns[52851] = 29'b1_100111001110_011_0_011100111011;
      patterns[52852] = 29'b1_100111001110_100_0_110011100111;
      patterns[52853] = 29'b1_100111001110_101_1_011001110011;
      patterns[52854] = 29'b1_100111001110_110_1_100111001110;
      patterns[52855] = 29'b1_100111001110_111_1_100111001110;
      patterns[52856] = 29'b1_100111001111_000_1_100111001111;
      patterns[52857] = 29'b1_100111001111_001_1_001111100111;
      patterns[52858] = 29'b1_100111001111_010_1_001110011111;
      patterns[52859] = 29'b1_100111001111_011_0_011100111111;
      patterns[52860] = 29'b1_100111001111_100_1_110011100111;
      patterns[52861] = 29'b1_100111001111_101_1_111001110011;
      patterns[52862] = 29'b1_100111001111_110_1_100111001111;
      patterns[52863] = 29'b1_100111001111_111_1_100111001111;
      patterns[52864] = 29'b1_100111010000_000_1_100111010000;
      patterns[52865] = 29'b1_100111010000_001_1_010000100111;
      patterns[52866] = 29'b1_100111010000_010_1_001110100001;
      patterns[52867] = 29'b1_100111010000_011_0_011101000011;
      patterns[52868] = 29'b1_100111010000_100_0_110011101000;
      patterns[52869] = 29'b1_100111010000_101_0_011001110100;
      patterns[52870] = 29'b1_100111010000_110_1_100111010000;
      patterns[52871] = 29'b1_100111010000_111_1_100111010000;
      patterns[52872] = 29'b1_100111010001_000_1_100111010001;
      patterns[52873] = 29'b1_100111010001_001_1_010001100111;
      patterns[52874] = 29'b1_100111010001_010_1_001110100011;
      patterns[52875] = 29'b1_100111010001_011_0_011101000111;
      patterns[52876] = 29'b1_100111010001_100_1_110011101000;
      patterns[52877] = 29'b1_100111010001_101_0_111001110100;
      patterns[52878] = 29'b1_100111010001_110_1_100111010001;
      patterns[52879] = 29'b1_100111010001_111_1_100111010001;
      patterns[52880] = 29'b1_100111010010_000_1_100111010010;
      patterns[52881] = 29'b1_100111010010_001_1_010010100111;
      patterns[52882] = 29'b1_100111010010_010_1_001110100101;
      patterns[52883] = 29'b1_100111010010_011_0_011101001011;
      patterns[52884] = 29'b1_100111010010_100_0_110011101001;
      patterns[52885] = 29'b1_100111010010_101_1_011001110100;
      patterns[52886] = 29'b1_100111010010_110_1_100111010010;
      patterns[52887] = 29'b1_100111010010_111_1_100111010010;
      patterns[52888] = 29'b1_100111010011_000_1_100111010011;
      patterns[52889] = 29'b1_100111010011_001_1_010011100111;
      patterns[52890] = 29'b1_100111010011_010_1_001110100111;
      patterns[52891] = 29'b1_100111010011_011_0_011101001111;
      patterns[52892] = 29'b1_100111010011_100_1_110011101001;
      patterns[52893] = 29'b1_100111010011_101_1_111001110100;
      patterns[52894] = 29'b1_100111010011_110_1_100111010011;
      patterns[52895] = 29'b1_100111010011_111_1_100111010011;
      patterns[52896] = 29'b1_100111010100_000_1_100111010100;
      patterns[52897] = 29'b1_100111010100_001_1_010100100111;
      patterns[52898] = 29'b1_100111010100_010_1_001110101001;
      patterns[52899] = 29'b1_100111010100_011_0_011101010011;
      patterns[52900] = 29'b1_100111010100_100_0_110011101010;
      patterns[52901] = 29'b1_100111010100_101_0_011001110101;
      patterns[52902] = 29'b1_100111010100_110_1_100111010100;
      patterns[52903] = 29'b1_100111010100_111_1_100111010100;
      patterns[52904] = 29'b1_100111010101_000_1_100111010101;
      patterns[52905] = 29'b1_100111010101_001_1_010101100111;
      patterns[52906] = 29'b1_100111010101_010_1_001110101011;
      patterns[52907] = 29'b1_100111010101_011_0_011101010111;
      patterns[52908] = 29'b1_100111010101_100_1_110011101010;
      patterns[52909] = 29'b1_100111010101_101_0_111001110101;
      patterns[52910] = 29'b1_100111010101_110_1_100111010101;
      patterns[52911] = 29'b1_100111010101_111_1_100111010101;
      patterns[52912] = 29'b1_100111010110_000_1_100111010110;
      patterns[52913] = 29'b1_100111010110_001_1_010110100111;
      patterns[52914] = 29'b1_100111010110_010_1_001110101101;
      patterns[52915] = 29'b1_100111010110_011_0_011101011011;
      patterns[52916] = 29'b1_100111010110_100_0_110011101011;
      patterns[52917] = 29'b1_100111010110_101_1_011001110101;
      patterns[52918] = 29'b1_100111010110_110_1_100111010110;
      patterns[52919] = 29'b1_100111010110_111_1_100111010110;
      patterns[52920] = 29'b1_100111010111_000_1_100111010111;
      patterns[52921] = 29'b1_100111010111_001_1_010111100111;
      patterns[52922] = 29'b1_100111010111_010_1_001110101111;
      patterns[52923] = 29'b1_100111010111_011_0_011101011111;
      patterns[52924] = 29'b1_100111010111_100_1_110011101011;
      patterns[52925] = 29'b1_100111010111_101_1_111001110101;
      patterns[52926] = 29'b1_100111010111_110_1_100111010111;
      patterns[52927] = 29'b1_100111010111_111_1_100111010111;
      patterns[52928] = 29'b1_100111011000_000_1_100111011000;
      patterns[52929] = 29'b1_100111011000_001_1_011000100111;
      patterns[52930] = 29'b1_100111011000_010_1_001110110001;
      patterns[52931] = 29'b1_100111011000_011_0_011101100011;
      patterns[52932] = 29'b1_100111011000_100_0_110011101100;
      patterns[52933] = 29'b1_100111011000_101_0_011001110110;
      patterns[52934] = 29'b1_100111011000_110_1_100111011000;
      patterns[52935] = 29'b1_100111011000_111_1_100111011000;
      patterns[52936] = 29'b1_100111011001_000_1_100111011001;
      patterns[52937] = 29'b1_100111011001_001_1_011001100111;
      patterns[52938] = 29'b1_100111011001_010_1_001110110011;
      patterns[52939] = 29'b1_100111011001_011_0_011101100111;
      patterns[52940] = 29'b1_100111011001_100_1_110011101100;
      patterns[52941] = 29'b1_100111011001_101_0_111001110110;
      patterns[52942] = 29'b1_100111011001_110_1_100111011001;
      patterns[52943] = 29'b1_100111011001_111_1_100111011001;
      patterns[52944] = 29'b1_100111011010_000_1_100111011010;
      patterns[52945] = 29'b1_100111011010_001_1_011010100111;
      patterns[52946] = 29'b1_100111011010_010_1_001110110101;
      patterns[52947] = 29'b1_100111011010_011_0_011101101011;
      patterns[52948] = 29'b1_100111011010_100_0_110011101101;
      patterns[52949] = 29'b1_100111011010_101_1_011001110110;
      patterns[52950] = 29'b1_100111011010_110_1_100111011010;
      patterns[52951] = 29'b1_100111011010_111_1_100111011010;
      patterns[52952] = 29'b1_100111011011_000_1_100111011011;
      patterns[52953] = 29'b1_100111011011_001_1_011011100111;
      patterns[52954] = 29'b1_100111011011_010_1_001110110111;
      patterns[52955] = 29'b1_100111011011_011_0_011101101111;
      patterns[52956] = 29'b1_100111011011_100_1_110011101101;
      patterns[52957] = 29'b1_100111011011_101_1_111001110110;
      patterns[52958] = 29'b1_100111011011_110_1_100111011011;
      patterns[52959] = 29'b1_100111011011_111_1_100111011011;
      patterns[52960] = 29'b1_100111011100_000_1_100111011100;
      patterns[52961] = 29'b1_100111011100_001_1_011100100111;
      patterns[52962] = 29'b1_100111011100_010_1_001110111001;
      patterns[52963] = 29'b1_100111011100_011_0_011101110011;
      patterns[52964] = 29'b1_100111011100_100_0_110011101110;
      patterns[52965] = 29'b1_100111011100_101_0_011001110111;
      patterns[52966] = 29'b1_100111011100_110_1_100111011100;
      patterns[52967] = 29'b1_100111011100_111_1_100111011100;
      patterns[52968] = 29'b1_100111011101_000_1_100111011101;
      patterns[52969] = 29'b1_100111011101_001_1_011101100111;
      patterns[52970] = 29'b1_100111011101_010_1_001110111011;
      patterns[52971] = 29'b1_100111011101_011_0_011101110111;
      patterns[52972] = 29'b1_100111011101_100_1_110011101110;
      patterns[52973] = 29'b1_100111011101_101_0_111001110111;
      patterns[52974] = 29'b1_100111011101_110_1_100111011101;
      patterns[52975] = 29'b1_100111011101_111_1_100111011101;
      patterns[52976] = 29'b1_100111011110_000_1_100111011110;
      patterns[52977] = 29'b1_100111011110_001_1_011110100111;
      patterns[52978] = 29'b1_100111011110_010_1_001110111101;
      patterns[52979] = 29'b1_100111011110_011_0_011101111011;
      patterns[52980] = 29'b1_100111011110_100_0_110011101111;
      patterns[52981] = 29'b1_100111011110_101_1_011001110111;
      patterns[52982] = 29'b1_100111011110_110_1_100111011110;
      patterns[52983] = 29'b1_100111011110_111_1_100111011110;
      patterns[52984] = 29'b1_100111011111_000_1_100111011111;
      patterns[52985] = 29'b1_100111011111_001_1_011111100111;
      patterns[52986] = 29'b1_100111011111_010_1_001110111111;
      patterns[52987] = 29'b1_100111011111_011_0_011101111111;
      patterns[52988] = 29'b1_100111011111_100_1_110011101111;
      patterns[52989] = 29'b1_100111011111_101_1_111001110111;
      patterns[52990] = 29'b1_100111011111_110_1_100111011111;
      patterns[52991] = 29'b1_100111011111_111_1_100111011111;
      patterns[52992] = 29'b1_100111100000_000_1_100111100000;
      patterns[52993] = 29'b1_100111100000_001_1_100000100111;
      patterns[52994] = 29'b1_100111100000_010_1_001111000001;
      patterns[52995] = 29'b1_100111100000_011_0_011110000011;
      patterns[52996] = 29'b1_100111100000_100_0_110011110000;
      patterns[52997] = 29'b1_100111100000_101_0_011001111000;
      patterns[52998] = 29'b1_100111100000_110_1_100111100000;
      patterns[52999] = 29'b1_100111100000_111_1_100111100000;
      patterns[53000] = 29'b1_100111100001_000_1_100111100001;
      patterns[53001] = 29'b1_100111100001_001_1_100001100111;
      patterns[53002] = 29'b1_100111100001_010_1_001111000011;
      patterns[53003] = 29'b1_100111100001_011_0_011110000111;
      patterns[53004] = 29'b1_100111100001_100_1_110011110000;
      patterns[53005] = 29'b1_100111100001_101_0_111001111000;
      patterns[53006] = 29'b1_100111100001_110_1_100111100001;
      patterns[53007] = 29'b1_100111100001_111_1_100111100001;
      patterns[53008] = 29'b1_100111100010_000_1_100111100010;
      patterns[53009] = 29'b1_100111100010_001_1_100010100111;
      patterns[53010] = 29'b1_100111100010_010_1_001111000101;
      patterns[53011] = 29'b1_100111100010_011_0_011110001011;
      patterns[53012] = 29'b1_100111100010_100_0_110011110001;
      patterns[53013] = 29'b1_100111100010_101_1_011001111000;
      patterns[53014] = 29'b1_100111100010_110_1_100111100010;
      patterns[53015] = 29'b1_100111100010_111_1_100111100010;
      patterns[53016] = 29'b1_100111100011_000_1_100111100011;
      patterns[53017] = 29'b1_100111100011_001_1_100011100111;
      patterns[53018] = 29'b1_100111100011_010_1_001111000111;
      patterns[53019] = 29'b1_100111100011_011_0_011110001111;
      patterns[53020] = 29'b1_100111100011_100_1_110011110001;
      patterns[53021] = 29'b1_100111100011_101_1_111001111000;
      patterns[53022] = 29'b1_100111100011_110_1_100111100011;
      patterns[53023] = 29'b1_100111100011_111_1_100111100011;
      patterns[53024] = 29'b1_100111100100_000_1_100111100100;
      patterns[53025] = 29'b1_100111100100_001_1_100100100111;
      patterns[53026] = 29'b1_100111100100_010_1_001111001001;
      patterns[53027] = 29'b1_100111100100_011_0_011110010011;
      patterns[53028] = 29'b1_100111100100_100_0_110011110010;
      patterns[53029] = 29'b1_100111100100_101_0_011001111001;
      patterns[53030] = 29'b1_100111100100_110_1_100111100100;
      patterns[53031] = 29'b1_100111100100_111_1_100111100100;
      patterns[53032] = 29'b1_100111100101_000_1_100111100101;
      patterns[53033] = 29'b1_100111100101_001_1_100101100111;
      patterns[53034] = 29'b1_100111100101_010_1_001111001011;
      patterns[53035] = 29'b1_100111100101_011_0_011110010111;
      patterns[53036] = 29'b1_100111100101_100_1_110011110010;
      patterns[53037] = 29'b1_100111100101_101_0_111001111001;
      patterns[53038] = 29'b1_100111100101_110_1_100111100101;
      patterns[53039] = 29'b1_100111100101_111_1_100111100101;
      patterns[53040] = 29'b1_100111100110_000_1_100111100110;
      patterns[53041] = 29'b1_100111100110_001_1_100110100111;
      patterns[53042] = 29'b1_100111100110_010_1_001111001101;
      patterns[53043] = 29'b1_100111100110_011_0_011110011011;
      patterns[53044] = 29'b1_100111100110_100_0_110011110011;
      patterns[53045] = 29'b1_100111100110_101_1_011001111001;
      patterns[53046] = 29'b1_100111100110_110_1_100111100110;
      patterns[53047] = 29'b1_100111100110_111_1_100111100110;
      patterns[53048] = 29'b1_100111100111_000_1_100111100111;
      patterns[53049] = 29'b1_100111100111_001_1_100111100111;
      patterns[53050] = 29'b1_100111100111_010_1_001111001111;
      patterns[53051] = 29'b1_100111100111_011_0_011110011111;
      patterns[53052] = 29'b1_100111100111_100_1_110011110011;
      patterns[53053] = 29'b1_100111100111_101_1_111001111001;
      patterns[53054] = 29'b1_100111100111_110_1_100111100111;
      patterns[53055] = 29'b1_100111100111_111_1_100111100111;
      patterns[53056] = 29'b1_100111101000_000_1_100111101000;
      patterns[53057] = 29'b1_100111101000_001_1_101000100111;
      patterns[53058] = 29'b1_100111101000_010_1_001111010001;
      patterns[53059] = 29'b1_100111101000_011_0_011110100011;
      patterns[53060] = 29'b1_100111101000_100_0_110011110100;
      patterns[53061] = 29'b1_100111101000_101_0_011001111010;
      patterns[53062] = 29'b1_100111101000_110_1_100111101000;
      patterns[53063] = 29'b1_100111101000_111_1_100111101000;
      patterns[53064] = 29'b1_100111101001_000_1_100111101001;
      patterns[53065] = 29'b1_100111101001_001_1_101001100111;
      patterns[53066] = 29'b1_100111101001_010_1_001111010011;
      patterns[53067] = 29'b1_100111101001_011_0_011110100111;
      patterns[53068] = 29'b1_100111101001_100_1_110011110100;
      patterns[53069] = 29'b1_100111101001_101_0_111001111010;
      patterns[53070] = 29'b1_100111101001_110_1_100111101001;
      patterns[53071] = 29'b1_100111101001_111_1_100111101001;
      patterns[53072] = 29'b1_100111101010_000_1_100111101010;
      patterns[53073] = 29'b1_100111101010_001_1_101010100111;
      patterns[53074] = 29'b1_100111101010_010_1_001111010101;
      patterns[53075] = 29'b1_100111101010_011_0_011110101011;
      patterns[53076] = 29'b1_100111101010_100_0_110011110101;
      patterns[53077] = 29'b1_100111101010_101_1_011001111010;
      patterns[53078] = 29'b1_100111101010_110_1_100111101010;
      patterns[53079] = 29'b1_100111101010_111_1_100111101010;
      patterns[53080] = 29'b1_100111101011_000_1_100111101011;
      patterns[53081] = 29'b1_100111101011_001_1_101011100111;
      patterns[53082] = 29'b1_100111101011_010_1_001111010111;
      patterns[53083] = 29'b1_100111101011_011_0_011110101111;
      patterns[53084] = 29'b1_100111101011_100_1_110011110101;
      patterns[53085] = 29'b1_100111101011_101_1_111001111010;
      patterns[53086] = 29'b1_100111101011_110_1_100111101011;
      patterns[53087] = 29'b1_100111101011_111_1_100111101011;
      patterns[53088] = 29'b1_100111101100_000_1_100111101100;
      patterns[53089] = 29'b1_100111101100_001_1_101100100111;
      patterns[53090] = 29'b1_100111101100_010_1_001111011001;
      patterns[53091] = 29'b1_100111101100_011_0_011110110011;
      patterns[53092] = 29'b1_100111101100_100_0_110011110110;
      patterns[53093] = 29'b1_100111101100_101_0_011001111011;
      patterns[53094] = 29'b1_100111101100_110_1_100111101100;
      patterns[53095] = 29'b1_100111101100_111_1_100111101100;
      patterns[53096] = 29'b1_100111101101_000_1_100111101101;
      patterns[53097] = 29'b1_100111101101_001_1_101101100111;
      patterns[53098] = 29'b1_100111101101_010_1_001111011011;
      patterns[53099] = 29'b1_100111101101_011_0_011110110111;
      patterns[53100] = 29'b1_100111101101_100_1_110011110110;
      patterns[53101] = 29'b1_100111101101_101_0_111001111011;
      patterns[53102] = 29'b1_100111101101_110_1_100111101101;
      patterns[53103] = 29'b1_100111101101_111_1_100111101101;
      patterns[53104] = 29'b1_100111101110_000_1_100111101110;
      patterns[53105] = 29'b1_100111101110_001_1_101110100111;
      patterns[53106] = 29'b1_100111101110_010_1_001111011101;
      patterns[53107] = 29'b1_100111101110_011_0_011110111011;
      patterns[53108] = 29'b1_100111101110_100_0_110011110111;
      patterns[53109] = 29'b1_100111101110_101_1_011001111011;
      patterns[53110] = 29'b1_100111101110_110_1_100111101110;
      patterns[53111] = 29'b1_100111101110_111_1_100111101110;
      patterns[53112] = 29'b1_100111101111_000_1_100111101111;
      patterns[53113] = 29'b1_100111101111_001_1_101111100111;
      patterns[53114] = 29'b1_100111101111_010_1_001111011111;
      patterns[53115] = 29'b1_100111101111_011_0_011110111111;
      patterns[53116] = 29'b1_100111101111_100_1_110011110111;
      patterns[53117] = 29'b1_100111101111_101_1_111001111011;
      patterns[53118] = 29'b1_100111101111_110_1_100111101111;
      patterns[53119] = 29'b1_100111101111_111_1_100111101111;
      patterns[53120] = 29'b1_100111110000_000_1_100111110000;
      patterns[53121] = 29'b1_100111110000_001_1_110000100111;
      patterns[53122] = 29'b1_100111110000_010_1_001111100001;
      patterns[53123] = 29'b1_100111110000_011_0_011111000011;
      patterns[53124] = 29'b1_100111110000_100_0_110011111000;
      patterns[53125] = 29'b1_100111110000_101_0_011001111100;
      patterns[53126] = 29'b1_100111110000_110_1_100111110000;
      patterns[53127] = 29'b1_100111110000_111_1_100111110000;
      patterns[53128] = 29'b1_100111110001_000_1_100111110001;
      patterns[53129] = 29'b1_100111110001_001_1_110001100111;
      patterns[53130] = 29'b1_100111110001_010_1_001111100011;
      patterns[53131] = 29'b1_100111110001_011_0_011111000111;
      patterns[53132] = 29'b1_100111110001_100_1_110011111000;
      patterns[53133] = 29'b1_100111110001_101_0_111001111100;
      patterns[53134] = 29'b1_100111110001_110_1_100111110001;
      patterns[53135] = 29'b1_100111110001_111_1_100111110001;
      patterns[53136] = 29'b1_100111110010_000_1_100111110010;
      patterns[53137] = 29'b1_100111110010_001_1_110010100111;
      patterns[53138] = 29'b1_100111110010_010_1_001111100101;
      patterns[53139] = 29'b1_100111110010_011_0_011111001011;
      patterns[53140] = 29'b1_100111110010_100_0_110011111001;
      patterns[53141] = 29'b1_100111110010_101_1_011001111100;
      patterns[53142] = 29'b1_100111110010_110_1_100111110010;
      patterns[53143] = 29'b1_100111110010_111_1_100111110010;
      patterns[53144] = 29'b1_100111110011_000_1_100111110011;
      patterns[53145] = 29'b1_100111110011_001_1_110011100111;
      patterns[53146] = 29'b1_100111110011_010_1_001111100111;
      patterns[53147] = 29'b1_100111110011_011_0_011111001111;
      patterns[53148] = 29'b1_100111110011_100_1_110011111001;
      patterns[53149] = 29'b1_100111110011_101_1_111001111100;
      patterns[53150] = 29'b1_100111110011_110_1_100111110011;
      patterns[53151] = 29'b1_100111110011_111_1_100111110011;
      patterns[53152] = 29'b1_100111110100_000_1_100111110100;
      patterns[53153] = 29'b1_100111110100_001_1_110100100111;
      patterns[53154] = 29'b1_100111110100_010_1_001111101001;
      patterns[53155] = 29'b1_100111110100_011_0_011111010011;
      patterns[53156] = 29'b1_100111110100_100_0_110011111010;
      patterns[53157] = 29'b1_100111110100_101_0_011001111101;
      patterns[53158] = 29'b1_100111110100_110_1_100111110100;
      patterns[53159] = 29'b1_100111110100_111_1_100111110100;
      patterns[53160] = 29'b1_100111110101_000_1_100111110101;
      patterns[53161] = 29'b1_100111110101_001_1_110101100111;
      patterns[53162] = 29'b1_100111110101_010_1_001111101011;
      patterns[53163] = 29'b1_100111110101_011_0_011111010111;
      patterns[53164] = 29'b1_100111110101_100_1_110011111010;
      patterns[53165] = 29'b1_100111110101_101_0_111001111101;
      patterns[53166] = 29'b1_100111110101_110_1_100111110101;
      patterns[53167] = 29'b1_100111110101_111_1_100111110101;
      patterns[53168] = 29'b1_100111110110_000_1_100111110110;
      patterns[53169] = 29'b1_100111110110_001_1_110110100111;
      patterns[53170] = 29'b1_100111110110_010_1_001111101101;
      patterns[53171] = 29'b1_100111110110_011_0_011111011011;
      patterns[53172] = 29'b1_100111110110_100_0_110011111011;
      patterns[53173] = 29'b1_100111110110_101_1_011001111101;
      patterns[53174] = 29'b1_100111110110_110_1_100111110110;
      patterns[53175] = 29'b1_100111110110_111_1_100111110110;
      patterns[53176] = 29'b1_100111110111_000_1_100111110111;
      patterns[53177] = 29'b1_100111110111_001_1_110111100111;
      patterns[53178] = 29'b1_100111110111_010_1_001111101111;
      patterns[53179] = 29'b1_100111110111_011_0_011111011111;
      patterns[53180] = 29'b1_100111110111_100_1_110011111011;
      patterns[53181] = 29'b1_100111110111_101_1_111001111101;
      patterns[53182] = 29'b1_100111110111_110_1_100111110111;
      patterns[53183] = 29'b1_100111110111_111_1_100111110111;
      patterns[53184] = 29'b1_100111111000_000_1_100111111000;
      patterns[53185] = 29'b1_100111111000_001_1_111000100111;
      patterns[53186] = 29'b1_100111111000_010_1_001111110001;
      patterns[53187] = 29'b1_100111111000_011_0_011111100011;
      patterns[53188] = 29'b1_100111111000_100_0_110011111100;
      patterns[53189] = 29'b1_100111111000_101_0_011001111110;
      patterns[53190] = 29'b1_100111111000_110_1_100111111000;
      patterns[53191] = 29'b1_100111111000_111_1_100111111000;
      patterns[53192] = 29'b1_100111111001_000_1_100111111001;
      patterns[53193] = 29'b1_100111111001_001_1_111001100111;
      patterns[53194] = 29'b1_100111111001_010_1_001111110011;
      patterns[53195] = 29'b1_100111111001_011_0_011111100111;
      patterns[53196] = 29'b1_100111111001_100_1_110011111100;
      patterns[53197] = 29'b1_100111111001_101_0_111001111110;
      patterns[53198] = 29'b1_100111111001_110_1_100111111001;
      patterns[53199] = 29'b1_100111111001_111_1_100111111001;
      patterns[53200] = 29'b1_100111111010_000_1_100111111010;
      patterns[53201] = 29'b1_100111111010_001_1_111010100111;
      patterns[53202] = 29'b1_100111111010_010_1_001111110101;
      patterns[53203] = 29'b1_100111111010_011_0_011111101011;
      patterns[53204] = 29'b1_100111111010_100_0_110011111101;
      patterns[53205] = 29'b1_100111111010_101_1_011001111110;
      patterns[53206] = 29'b1_100111111010_110_1_100111111010;
      patterns[53207] = 29'b1_100111111010_111_1_100111111010;
      patterns[53208] = 29'b1_100111111011_000_1_100111111011;
      patterns[53209] = 29'b1_100111111011_001_1_111011100111;
      patterns[53210] = 29'b1_100111111011_010_1_001111110111;
      patterns[53211] = 29'b1_100111111011_011_0_011111101111;
      patterns[53212] = 29'b1_100111111011_100_1_110011111101;
      patterns[53213] = 29'b1_100111111011_101_1_111001111110;
      patterns[53214] = 29'b1_100111111011_110_1_100111111011;
      patterns[53215] = 29'b1_100111111011_111_1_100111111011;
      patterns[53216] = 29'b1_100111111100_000_1_100111111100;
      patterns[53217] = 29'b1_100111111100_001_1_111100100111;
      patterns[53218] = 29'b1_100111111100_010_1_001111111001;
      patterns[53219] = 29'b1_100111111100_011_0_011111110011;
      patterns[53220] = 29'b1_100111111100_100_0_110011111110;
      patterns[53221] = 29'b1_100111111100_101_0_011001111111;
      patterns[53222] = 29'b1_100111111100_110_1_100111111100;
      patterns[53223] = 29'b1_100111111100_111_1_100111111100;
      patterns[53224] = 29'b1_100111111101_000_1_100111111101;
      patterns[53225] = 29'b1_100111111101_001_1_111101100111;
      patterns[53226] = 29'b1_100111111101_010_1_001111111011;
      patterns[53227] = 29'b1_100111111101_011_0_011111110111;
      patterns[53228] = 29'b1_100111111101_100_1_110011111110;
      patterns[53229] = 29'b1_100111111101_101_0_111001111111;
      patterns[53230] = 29'b1_100111111101_110_1_100111111101;
      patterns[53231] = 29'b1_100111111101_111_1_100111111101;
      patterns[53232] = 29'b1_100111111110_000_1_100111111110;
      patterns[53233] = 29'b1_100111111110_001_1_111110100111;
      patterns[53234] = 29'b1_100111111110_010_1_001111111101;
      patterns[53235] = 29'b1_100111111110_011_0_011111111011;
      patterns[53236] = 29'b1_100111111110_100_0_110011111111;
      patterns[53237] = 29'b1_100111111110_101_1_011001111111;
      patterns[53238] = 29'b1_100111111110_110_1_100111111110;
      patterns[53239] = 29'b1_100111111110_111_1_100111111110;
      patterns[53240] = 29'b1_100111111111_000_1_100111111111;
      patterns[53241] = 29'b1_100111111111_001_1_111111100111;
      patterns[53242] = 29'b1_100111111111_010_1_001111111111;
      patterns[53243] = 29'b1_100111111111_011_0_011111111111;
      patterns[53244] = 29'b1_100111111111_100_1_110011111111;
      patterns[53245] = 29'b1_100111111111_101_1_111001111111;
      patterns[53246] = 29'b1_100111111111_110_1_100111111111;
      patterns[53247] = 29'b1_100111111111_111_1_100111111111;
      patterns[53248] = 29'b1_101000000000_000_1_101000000000;
      patterns[53249] = 29'b1_101000000000_001_1_000000101000;
      patterns[53250] = 29'b1_101000000000_010_1_010000000001;
      patterns[53251] = 29'b1_101000000000_011_0_100000000011;
      patterns[53252] = 29'b1_101000000000_100_0_110100000000;
      patterns[53253] = 29'b1_101000000000_101_0_011010000000;
      patterns[53254] = 29'b1_101000000000_110_1_101000000000;
      patterns[53255] = 29'b1_101000000000_111_1_101000000000;
      patterns[53256] = 29'b1_101000000001_000_1_101000000001;
      patterns[53257] = 29'b1_101000000001_001_1_000001101000;
      patterns[53258] = 29'b1_101000000001_010_1_010000000011;
      patterns[53259] = 29'b1_101000000001_011_0_100000000111;
      patterns[53260] = 29'b1_101000000001_100_1_110100000000;
      patterns[53261] = 29'b1_101000000001_101_0_111010000000;
      patterns[53262] = 29'b1_101000000001_110_1_101000000001;
      patterns[53263] = 29'b1_101000000001_111_1_101000000001;
      patterns[53264] = 29'b1_101000000010_000_1_101000000010;
      patterns[53265] = 29'b1_101000000010_001_1_000010101000;
      patterns[53266] = 29'b1_101000000010_010_1_010000000101;
      patterns[53267] = 29'b1_101000000010_011_0_100000001011;
      patterns[53268] = 29'b1_101000000010_100_0_110100000001;
      patterns[53269] = 29'b1_101000000010_101_1_011010000000;
      patterns[53270] = 29'b1_101000000010_110_1_101000000010;
      patterns[53271] = 29'b1_101000000010_111_1_101000000010;
      patterns[53272] = 29'b1_101000000011_000_1_101000000011;
      patterns[53273] = 29'b1_101000000011_001_1_000011101000;
      patterns[53274] = 29'b1_101000000011_010_1_010000000111;
      patterns[53275] = 29'b1_101000000011_011_0_100000001111;
      patterns[53276] = 29'b1_101000000011_100_1_110100000001;
      patterns[53277] = 29'b1_101000000011_101_1_111010000000;
      patterns[53278] = 29'b1_101000000011_110_1_101000000011;
      patterns[53279] = 29'b1_101000000011_111_1_101000000011;
      patterns[53280] = 29'b1_101000000100_000_1_101000000100;
      patterns[53281] = 29'b1_101000000100_001_1_000100101000;
      patterns[53282] = 29'b1_101000000100_010_1_010000001001;
      patterns[53283] = 29'b1_101000000100_011_0_100000010011;
      patterns[53284] = 29'b1_101000000100_100_0_110100000010;
      patterns[53285] = 29'b1_101000000100_101_0_011010000001;
      patterns[53286] = 29'b1_101000000100_110_1_101000000100;
      patterns[53287] = 29'b1_101000000100_111_1_101000000100;
      patterns[53288] = 29'b1_101000000101_000_1_101000000101;
      patterns[53289] = 29'b1_101000000101_001_1_000101101000;
      patterns[53290] = 29'b1_101000000101_010_1_010000001011;
      patterns[53291] = 29'b1_101000000101_011_0_100000010111;
      patterns[53292] = 29'b1_101000000101_100_1_110100000010;
      patterns[53293] = 29'b1_101000000101_101_0_111010000001;
      patterns[53294] = 29'b1_101000000101_110_1_101000000101;
      patterns[53295] = 29'b1_101000000101_111_1_101000000101;
      patterns[53296] = 29'b1_101000000110_000_1_101000000110;
      patterns[53297] = 29'b1_101000000110_001_1_000110101000;
      patterns[53298] = 29'b1_101000000110_010_1_010000001101;
      patterns[53299] = 29'b1_101000000110_011_0_100000011011;
      patterns[53300] = 29'b1_101000000110_100_0_110100000011;
      patterns[53301] = 29'b1_101000000110_101_1_011010000001;
      patterns[53302] = 29'b1_101000000110_110_1_101000000110;
      patterns[53303] = 29'b1_101000000110_111_1_101000000110;
      patterns[53304] = 29'b1_101000000111_000_1_101000000111;
      patterns[53305] = 29'b1_101000000111_001_1_000111101000;
      patterns[53306] = 29'b1_101000000111_010_1_010000001111;
      patterns[53307] = 29'b1_101000000111_011_0_100000011111;
      patterns[53308] = 29'b1_101000000111_100_1_110100000011;
      patterns[53309] = 29'b1_101000000111_101_1_111010000001;
      patterns[53310] = 29'b1_101000000111_110_1_101000000111;
      patterns[53311] = 29'b1_101000000111_111_1_101000000111;
      patterns[53312] = 29'b1_101000001000_000_1_101000001000;
      patterns[53313] = 29'b1_101000001000_001_1_001000101000;
      patterns[53314] = 29'b1_101000001000_010_1_010000010001;
      patterns[53315] = 29'b1_101000001000_011_0_100000100011;
      patterns[53316] = 29'b1_101000001000_100_0_110100000100;
      patterns[53317] = 29'b1_101000001000_101_0_011010000010;
      patterns[53318] = 29'b1_101000001000_110_1_101000001000;
      patterns[53319] = 29'b1_101000001000_111_1_101000001000;
      patterns[53320] = 29'b1_101000001001_000_1_101000001001;
      patterns[53321] = 29'b1_101000001001_001_1_001001101000;
      patterns[53322] = 29'b1_101000001001_010_1_010000010011;
      patterns[53323] = 29'b1_101000001001_011_0_100000100111;
      patterns[53324] = 29'b1_101000001001_100_1_110100000100;
      patterns[53325] = 29'b1_101000001001_101_0_111010000010;
      patterns[53326] = 29'b1_101000001001_110_1_101000001001;
      patterns[53327] = 29'b1_101000001001_111_1_101000001001;
      patterns[53328] = 29'b1_101000001010_000_1_101000001010;
      patterns[53329] = 29'b1_101000001010_001_1_001010101000;
      patterns[53330] = 29'b1_101000001010_010_1_010000010101;
      patterns[53331] = 29'b1_101000001010_011_0_100000101011;
      patterns[53332] = 29'b1_101000001010_100_0_110100000101;
      patterns[53333] = 29'b1_101000001010_101_1_011010000010;
      patterns[53334] = 29'b1_101000001010_110_1_101000001010;
      patterns[53335] = 29'b1_101000001010_111_1_101000001010;
      patterns[53336] = 29'b1_101000001011_000_1_101000001011;
      patterns[53337] = 29'b1_101000001011_001_1_001011101000;
      patterns[53338] = 29'b1_101000001011_010_1_010000010111;
      patterns[53339] = 29'b1_101000001011_011_0_100000101111;
      patterns[53340] = 29'b1_101000001011_100_1_110100000101;
      patterns[53341] = 29'b1_101000001011_101_1_111010000010;
      patterns[53342] = 29'b1_101000001011_110_1_101000001011;
      patterns[53343] = 29'b1_101000001011_111_1_101000001011;
      patterns[53344] = 29'b1_101000001100_000_1_101000001100;
      patterns[53345] = 29'b1_101000001100_001_1_001100101000;
      patterns[53346] = 29'b1_101000001100_010_1_010000011001;
      patterns[53347] = 29'b1_101000001100_011_0_100000110011;
      patterns[53348] = 29'b1_101000001100_100_0_110100000110;
      patterns[53349] = 29'b1_101000001100_101_0_011010000011;
      patterns[53350] = 29'b1_101000001100_110_1_101000001100;
      patterns[53351] = 29'b1_101000001100_111_1_101000001100;
      patterns[53352] = 29'b1_101000001101_000_1_101000001101;
      patterns[53353] = 29'b1_101000001101_001_1_001101101000;
      patterns[53354] = 29'b1_101000001101_010_1_010000011011;
      patterns[53355] = 29'b1_101000001101_011_0_100000110111;
      patterns[53356] = 29'b1_101000001101_100_1_110100000110;
      patterns[53357] = 29'b1_101000001101_101_0_111010000011;
      patterns[53358] = 29'b1_101000001101_110_1_101000001101;
      patterns[53359] = 29'b1_101000001101_111_1_101000001101;
      patterns[53360] = 29'b1_101000001110_000_1_101000001110;
      patterns[53361] = 29'b1_101000001110_001_1_001110101000;
      patterns[53362] = 29'b1_101000001110_010_1_010000011101;
      patterns[53363] = 29'b1_101000001110_011_0_100000111011;
      patterns[53364] = 29'b1_101000001110_100_0_110100000111;
      patterns[53365] = 29'b1_101000001110_101_1_011010000011;
      patterns[53366] = 29'b1_101000001110_110_1_101000001110;
      patterns[53367] = 29'b1_101000001110_111_1_101000001110;
      patterns[53368] = 29'b1_101000001111_000_1_101000001111;
      patterns[53369] = 29'b1_101000001111_001_1_001111101000;
      patterns[53370] = 29'b1_101000001111_010_1_010000011111;
      patterns[53371] = 29'b1_101000001111_011_0_100000111111;
      patterns[53372] = 29'b1_101000001111_100_1_110100000111;
      patterns[53373] = 29'b1_101000001111_101_1_111010000011;
      patterns[53374] = 29'b1_101000001111_110_1_101000001111;
      patterns[53375] = 29'b1_101000001111_111_1_101000001111;
      patterns[53376] = 29'b1_101000010000_000_1_101000010000;
      patterns[53377] = 29'b1_101000010000_001_1_010000101000;
      patterns[53378] = 29'b1_101000010000_010_1_010000100001;
      patterns[53379] = 29'b1_101000010000_011_0_100001000011;
      patterns[53380] = 29'b1_101000010000_100_0_110100001000;
      patterns[53381] = 29'b1_101000010000_101_0_011010000100;
      patterns[53382] = 29'b1_101000010000_110_1_101000010000;
      patterns[53383] = 29'b1_101000010000_111_1_101000010000;
      patterns[53384] = 29'b1_101000010001_000_1_101000010001;
      patterns[53385] = 29'b1_101000010001_001_1_010001101000;
      patterns[53386] = 29'b1_101000010001_010_1_010000100011;
      patterns[53387] = 29'b1_101000010001_011_0_100001000111;
      patterns[53388] = 29'b1_101000010001_100_1_110100001000;
      patterns[53389] = 29'b1_101000010001_101_0_111010000100;
      patterns[53390] = 29'b1_101000010001_110_1_101000010001;
      patterns[53391] = 29'b1_101000010001_111_1_101000010001;
      patterns[53392] = 29'b1_101000010010_000_1_101000010010;
      patterns[53393] = 29'b1_101000010010_001_1_010010101000;
      patterns[53394] = 29'b1_101000010010_010_1_010000100101;
      patterns[53395] = 29'b1_101000010010_011_0_100001001011;
      patterns[53396] = 29'b1_101000010010_100_0_110100001001;
      patterns[53397] = 29'b1_101000010010_101_1_011010000100;
      patterns[53398] = 29'b1_101000010010_110_1_101000010010;
      patterns[53399] = 29'b1_101000010010_111_1_101000010010;
      patterns[53400] = 29'b1_101000010011_000_1_101000010011;
      patterns[53401] = 29'b1_101000010011_001_1_010011101000;
      patterns[53402] = 29'b1_101000010011_010_1_010000100111;
      patterns[53403] = 29'b1_101000010011_011_0_100001001111;
      patterns[53404] = 29'b1_101000010011_100_1_110100001001;
      patterns[53405] = 29'b1_101000010011_101_1_111010000100;
      patterns[53406] = 29'b1_101000010011_110_1_101000010011;
      patterns[53407] = 29'b1_101000010011_111_1_101000010011;
      patterns[53408] = 29'b1_101000010100_000_1_101000010100;
      patterns[53409] = 29'b1_101000010100_001_1_010100101000;
      patterns[53410] = 29'b1_101000010100_010_1_010000101001;
      patterns[53411] = 29'b1_101000010100_011_0_100001010011;
      patterns[53412] = 29'b1_101000010100_100_0_110100001010;
      patterns[53413] = 29'b1_101000010100_101_0_011010000101;
      patterns[53414] = 29'b1_101000010100_110_1_101000010100;
      patterns[53415] = 29'b1_101000010100_111_1_101000010100;
      patterns[53416] = 29'b1_101000010101_000_1_101000010101;
      patterns[53417] = 29'b1_101000010101_001_1_010101101000;
      patterns[53418] = 29'b1_101000010101_010_1_010000101011;
      patterns[53419] = 29'b1_101000010101_011_0_100001010111;
      patterns[53420] = 29'b1_101000010101_100_1_110100001010;
      patterns[53421] = 29'b1_101000010101_101_0_111010000101;
      patterns[53422] = 29'b1_101000010101_110_1_101000010101;
      patterns[53423] = 29'b1_101000010101_111_1_101000010101;
      patterns[53424] = 29'b1_101000010110_000_1_101000010110;
      patterns[53425] = 29'b1_101000010110_001_1_010110101000;
      patterns[53426] = 29'b1_101000010110_010_1_010000101101;
      patterns[53427] = 29'b1_101000010110_011_0_100001011011;
      patterns[53428] = 29'b1_101000010110_100_0_110100001011;
      patterns[53429] = 29'b1_101000010110_101_1_011010000101;
      patterns[53430] = 29'b1_101000010110_110_1_101000010110;
      patterns[53431] = 29'b1_101000010110_111_1_101000010110;
      patterns[53432] = 29'b1_101000010111_000_1_101000010111;
      patterns[53433] = 29'b1_101000010111_001_1_010111101000;
      patterns[53434] = 29'b1_101000010111_010_1_010000101111;
      patterns[53435] = 29'b1_101000010111_011_0_100001011111;
      patterns[53436] = 29'b1_101000010111_100_1_110100001011;
      patterns[53437] = 29'b1_101000010111_101_1_111010000101;
      patterns[53438] = 29'b1_101000010111_110_1_101000010111;
      patterns[53439] = 29'b1_101000010111_111_1_101000010111;
      patterns[53440] = 29'b1_101000011000_000_1_101000011000;
      patterns[53441] = 29'b1_101000011000_001_1_011000101000;
      patterns[53442] = 29'b1_101000011000_010_1_010000110001;
      patterns[53443] = 29'b1_101000011000_011_0_100001100011;
      patterns[53444] = 29'b1_101000011000_100_0_110100001100;
      patterns[53445] = 29'b1_101000011000_101_0_011010000110;
      patterns[53446] = 29'b1_101000011000_110_1_101000011000;
      patterns[53447] = 29'b1_101000011000_111_1_101000011000;
      patterns[53448] = 29'b1_101000011001_000_1_101000011001;
      patterns[53449] = 29'b1_101000011001_001_1_011001101000;
      patterns[53450] = 29'b1_101000011001_010_1_010000110011;
      patterns[53451] = 29'b1_101000011001_011_0_100001100111;
      patterns[53452] = 29'b1_101000011001_100_1_110100001100;
      patterns[53453] = 29'b1_101000011001_101_0_111010000110;
      patterns[53454] = 29'b1_101000011001_110_1_101000011001;
      patterns[53455] = 29'b1_101000011001_111_1_101000011001;
      patterns[53456] = 29'b1_101000011010_000_1_101000011010;
      patterns[53457] = 29'b1_101000011010_001_1_011010101000;
      patterns[53458] = 29'b1_101000011010_010_1_010000110101;
      patterns[53459] = 29'b1_101000011010_011_0_100001101011;
      patterns[53460] = 29'b1_101000011010_100_0_110100001101;
      patterns[53461] = 29'b1_101000011010_101_1_011010000110;
      patterns[53462] = 29'b1_101000011010_110_1_101000011010;
      patterns[53463] = 29'b1_101000011010_111_1_101000011010;
      patterns[53464] = 29'b1_101000011011_000_1_101000011011;
      patterns[53465] = 29'b1_101000011011_001_1_011011101000;
      patterns[53466] = 29'b1_101000011011_010_1_010000110111;
      patterns[53467] = 29'b1_101000011011_011_0_100001101111;
      patterns[53468] = 29'b1_101000011011_100_1_110100001101;
      patterns[53469] = 29'b1_101000011011_101_1_111010000110;
      patterns[53470] = 29'b1_101000011011_110_1_101000011011;
      patterns[53471] = 29'b1_101000011011_111_1_101000011011;
      patterns[53472] = 29'b1_101000011100_000_1_101000011100;
      patterns[53473] = 29'b1_101000011100_001_1_011100101000;
      patterns[53474] = 29'b1_101000011100_010_1_010000111001;
      patterns[53475] = 29'b1_101000011100_011_0_100001110011;
      patterns[53476] = 29'b1_101000011100_100_0_110100001110;
      patterns[53477] = 29'b1_101000011100_101_0_011010000111;
      patterns[53478] = 29'b1_101000011100_110_1_101000011100;
      patterns[53479] = 29'b1_101000011100_111_1_101000011100;
      patterns[53480] = 29'b1_101000011101_000_1_101000011101;
      patterns[53481] = 29'b1_101000011101_001_1_011101101000;
      patterns[53482] = 29'b1_101000011101_010_1_010000111011;
      patterns[53483] = 29'b1_101000011101_011_0_100001110111;
      patterns[53484] = 29'b1_101000011101_100_1_110100001110;
      patterns[53485] = 29'b1_101000011101_101_0_111010000111;
      patterns[53486] = 29'b1_101000011101_110_1_101000011101;
      patterns[53487] = 29'b1_101000011101_111_1_101000011101;
      patterns[53488] = 29'b1_101000011110_000_1_101000011110;
      patterns[53489] = 29'b1_101000011110_001_1_011110101000;
      patterns[53490] = 29'b1_101000011110_010_1_010000111101;
      patterns[53491] = 29'b1_101000011110_011_0_100001111011;
      patterns[53492] = 29'b1_101000011110_100_0_110100001111;
      patterns[53493] = 29'b1_101000011110_101_1_011010000111;
      patterns[53494] = 29'b1_101000011110_110_1_101000011110;
      patterns[53495] = 29'b1_101000011110_111_1_101000011110;
      patterns[53496] = 29'b1_101000011111_000_1_101000011111;
      patterns[53497] = 29'b1_101000011111_001_1_011111101000;
      patterns[53498] = 29'b1_101000011111_010_1_010000111111;
      patterns[53499] = 29'b1_101000011111_011_0_100001111111;
      patterns[53500] = 29'b1_101000011111_100_1_110100001111;
      patterns[53501] = 29'b1_101000011111_101_1_111010000111;
      patterns[53502] = 29'b1_101000011111_110_1_101000011111;
      patterns[53503] = 29'b1_101000011111_111_1_101000011111;
      patterns[53504] = 29'b1_101000100000_000_1_101000100000;
      patterns[53505] = 29'b1_101000100000_001_1_100000101000;
      patterns[53506] = 29'b1_101000100000_010_1_010001000001;
      patterns[53507] = 29'b1_101000100000_011_0_100010000011;
      patterns[53508] = 29'b1_101000100000_100_0_110100010000;
      patterns[53509] = 29'b1_101000100000_101_0_011010001000;
      patterns[53510] = 29'b1_101000100000_110_1_101000100000;
      patterns[53511] = 29'b1_101000100000_111_1_101000100000;
      patterns[53512] = 29'b1_101000100001_000_1_101000100001;
      patterns[53513] = 29'b1_101000100001_001_1_100001101000;
      patterns[53514] = 29'b1_101000100001_010_1_010001000011;
      patterns[53515] = 29'b1_101000100001_011_0_100010000111;
      patterns[53516] = 29'b1_101000100001_100_1_110100010000;
      patterns[53517] = 29'b1_101000100001_101_0_111010001000;
      patterns[53518] = 29'b1_101000100001_110_1_101000100001;
      patterns[53519] = 29'b1_101000100001_111_1_101000100001;
      patterns[53520] = 29'b1_101000100010_000_1_101000100010;
      patterns[53521] = 29'b1_101000100010_001_1_100010101000;
      patterns[53522] = 29'b1_101000100010_010_1_010001000101;
      patterns[53523] = 29'b1_101000100010_011_0_100010001011;
      patterns[53524] = 29'b1_101000100010_100_0_110100010001;
      patterns[53525] = 29'b1_101000100010_101_1_011010001000;
      patterns[53526] = 29'b1_101000100010_110_1_101000100010;
      patterns[53527] = 29'b1_101000100010_111_1_101000100010;
      patterns[53528] = 29'b1_101000100011_000_1_101000100011;
      patterns[53529] = 29'b1_101000100011_001_1_100011101000;
      patterns[53530] = 29'b1_101000100011_010_1_010001000111;
      patterns[53531] = 29'b1_101000100011_011_0_100010001111;
      patterns[53532] = 29'b1_101000100011_100_1_110100010001;
      patterns[53533] = 29'b1_101000100011_101_1_111010001000;
      patterns[53534] = 29'b1_101000100011_110_1_101000100011;
      patterns[53535] = 29'b1_101000100011_111_1_101000100011;
      patterns[53536] = 29'b1_101000100100_000_1_101000100100;
      patterns[53537] = 29'b1_101000100100_001_1_100100101000;
      patterns[53538] = 29'b1_101000100100_010_1_010001001001;
      patterns[53539] = 29'b1_101000100100_011_0_100010010011;
      patterns[53540] = 29'b1_101000100100_100_0_110100010010;
      patterns[53541] = 29'b1_101000100100_101_0_011010001001;
      patterns[53542] = 29'b1_101000100100_110_1_101000100100;
      patterns[53543] = 29'b1_101000100100_111_1_101000100100;
      patterns[53544] = 29'b1_101000100101_000_1_101000100101;
      patterns[53545] = 29'b1_101000100101_001_1_100101101000;
      patterns[53546] = 29'b1_101000100101_010_1_010001001011;
      patterns[53547] = 29'b1_101000100101_011_0_100010010111;
      patterns[53548] = 29'b1_101000100101_100_1_110100010010;
      patterns[53549] = 29'b1_101000100101_101_0_111010001001;
      patterns[53550] = 29'b1_101000100101_110_1_101000100101;
      patterns[53551] = 29'b1_101000100101_111_1_101000100101;
      patterns[53552] = 29'b1_101000100110_000_1_101000100110;
      patterns[53553] = 29'b1_101000100110_001_1_100110101000;
      patterns[53554] = 29'b1_101000100110_010_1_010001001101;
      patterns[53555] = 29'b1_101000100110_011_0_100010011011;
      patterns[53556] = 29'b1_101000100110_100_0_110100010011;
      patterns[53557] = 29'b1_101000100110_101_1_011010001001;
      patterns[53558] = 29'b1_101000100110_110_1_101000100110;
      patterns[53559] = 29'b1_101000100110_111_1_101000100110;
      patterns[53560] = 29'b1_101000100111_000_1_101000100111;
      patterns[53561] = 29'b1_101000100111_001_1_100111101000;
      patterns[53562] = 29'b1_101000100111_010_1_010001001111;
      patterns[53563] = 29'b1_101000100111_011_0_100010011111;
      patterns[53564] = 29'b1_101000100111_100_1_110100010011;
      patterns[53565] = 29'b1_101000100111_101_1_111010001001;
      patterns[53566] = 29'b1_101000100111_110_1_101000100111;
      patterns[53567] = 29'b1_101000100111_111_1_101000100111;
      patterns[53568] = 29'b1_101000101000_000_1_101000101000;
      patterns[53569] = 29'b1_101000101000_001_1_101000101000;
      patterns[53570] = 29'b1_101000101000_010_1_010001010001;
      patterns[53571] = 29'b1_101000101000_011_0_100010100011;
      patterns[53572] = 29'b1_101000101000_100_0_110100010100;
      patterns[53573] = 29'b1_101000101000_101_0_011010001010;
      patterns[53574] = 29'b1_101000101000_110_1_101000101000;
      patterns[53575] = 29'b1_101000101000_111_1_101000101000;
      patterns[53576] = 29'b1_101000101001_000_1_101000101001;
      patterns[53577] = 29'b1_101000101001_001_1_101001101000;
      patterns[53578] = 29'b1_101000101001_010_1_010001010011;
      patterns[53579] = 29'b1_101000101001_011_0_100010100111;
      patterns[53580] = 29'b1_101000101001_100_1_110100010100;
      patterns[53581] = 29'b1_101000101001_101_0_111010001010;
      patterns[53582] = 29'b1_101000101001_110_1_101000101001;
      patterns[53583] = 29'b1_101000101001_111_1_101000101001;
      patterns[53584] = 29'b1_101000101010_000_1_101000101010;
      patterns[53585] = 29'b1_101000101010_001_1_101010101000;
      patterns[53586] = 29'b1_101000101010_010_1_010001010101;
      patterns[53587] = 29'b1_101000101010_011_0_100010101011;
      patterns[53588] = 29'b1_101000101010_100_0_110100010101;
      patterns[53589] = 29'b1_101000101010_101_1_011010001010;
      patterns[53590] = 29'b1_101000101010_110_1_101000101010;
      patterns[53591] = 29'b1_101000101010_111_1_101000101010;
      patterns[53592] = 29'b1_101000101011_000_1_101000101011;
      patterns[53593] = 29'b1_101000101011_001_1_101011101000;
      patterns[53594] = 29'b1_101000101011_010_1_010001010111;
      patterns[53595] = 29'b1_101000101011_011_0_100010101111;
      patterns[53596] = 29'b1_101000101011_100_1_110100010101;
      patterns[53597] = 29'b1_101000101011_101_1_111010001010;
      patterns[53598] = 29'b1_101000101011_110_1_101000101011;
      patterns[53599] = 29'b1_101000101011_111_1_101000101011;
      patterns[53600] = 29'b1_101000101100_000_1_101000101100;
      patterns[53601] = 29'b1_101000101100_001_1_101100101000;
      patterns[53602] = 29'b1_101000101100_010_1_010001011001;
      patterns[53603] = 29'b1_101000101100_011_0_100010110011;
      patterns[53604] = 29'b1_101000101100_100_0_110100010110;
      patterns[53605] = 29'b1_101000101100_101_0_011010001011;
      patterns[53606] = 29'b1_101000101100_110_1_101000101100;
      patterns[53607] = 29'b1_101000101100_111_1_101000101100;
      patterns[53608] = 29'b1_101000101101_000_1_101000101101;
      patterns[53609] = 29'b1_101000101101_001_1_101101101000;
      patterns[53610] = 29'b1_101000101101_010_1_010001011011;
      patterns[53611] = 29'b1_101000101101_011_0_100010110111;
      patterns[53612] = 29'b1_101000101101_100_1_110100010110;
      patterns[53613] = 29'b1_101000101101_101_0_111010001011;
      patterns[53614] = 29'b1_101000101101_110_1_101000101101;
      patterns[53615] = 29'b1_101000101101_111_1_101000101101;
      patterns[53616] = 29'b1_101000101110_000_1_101000101110;
      patterns[53617] = 29'b1_101000101110_001_1_101110101000;
      patterns[53618] = 29'b1_101000101110_010_1_010001011101;
      patterns[53619] = 29'b1_101000101110_011_0_100010111011;
      patterns[53620] = 29'b1_101000101110_100_0_110100010111;
      patterns[53621] = 29'b1_101000101110_101_1_011010001011;
      patterns[53622] = 29'b1_101000101110_110_1_101000101110;
      patterns[53623] = 29'b1_101000101110_111_1_101000101110;
      patterns[53624] = 29'b1_101000101111_000_1_101000101111;
      patterns[53625] = 29'b1_101000101111_001_1_101111101000;
      patterns[53626] = 29'b1_101000101111_010_1_010001011111;
      patterns[53627] = 29'b1_101000101111_011_0_100010111111;
      patterns[53628] = 29'b1_101000101111_100_1_110100010111;
      patterns[53629] = 29'b1_101000101111_101_1_111010001011;
      patterns[53630] = 29'b1_101000101111_110_1_101000101111;
      patterns[53631] = 29'b1_101000101111_111_1_101000101111;
      patterns[53632] = 29'b1_101000110000_000_1_101000110000;
      patterns[53633] = 29'b1_101000110000_001_1_110000101000;
      patterns[53634] = 29'b1_101000110000_010_1_010001100001;
      patterns[53635] = 29'b1_101000110000_011_0_100011000011;
      patterns[53636] = 29'b1_101000110000_100_0_110100011000;
      patterns[53637] = 29'b1_101000110000_101_0_011010001100;
      patterns[53638] = 29'b1_101000110000_110_1_101000110000;
      patterns[53639] = 29'b1_101000110000_111_1_101000110000;
      patterns[53640] = 29'b1_101000110001_000_1_101000110001;
      patterns[53641] = 29'b1_101000110001_001_1_110001101000;
      patterns[53642] = 29'b1_101000110001_010_1_010001100011;
      patterns[53643] = 29'b1_101000110001_011_0_100011000111;
      patterns[53644] = 29'b1_101000110001_100_1_110100011000;
      patterns[53645] = 29'b1_101000110001_101_0_111010001100;
      patterns[53646] = 29'b1_101000110001_110_1_101000110001;
      patterns[53647] = 29'b1_101000110001_111_1_101000110001;
      patterns[53648] = 29'b1_101000110010_000_1_101000110010;
      patterns[53649] = 29'b1_101000110010_001_1_110010101000;
      patterns[53650] = 29'b1_101000110010_010_1_010001100101;
      patterns[53651] = 29'b1_101000110010_011_0_100011001011;
      patterns[53652] = 29'b1_101000110010_100_0_110100011001;
      patterns[53653] = 29'b1_101000110010_101_1_011010001100;
      patterns[53654] = 29'b1_101000110010_110_1_101000110010;
      patterns[53655] = 29'b1_101000110010_111_1_101000110010;
      patterns[53656] = 29'b1_101000110011_000_1_101000110011;
      patterns[53657] = 29'b1_101000110011_001_1_110011101000;
      patterns[53658] = 29'b1_101000110011_010_1_010001100111;
      patterns[53659] = 29'b1_101000110011_011_0_100011001111;
      patterns[53660] = 29'b1_101000110011_100_1_110100011001;
      patterns[53661] = 29'b1_101000110011_101_1_111010001100;
      patterns[53662] = 29'b1_101000110011_110_1_101000110011;
      patterns[53663] = 29'b1_101000110011_111_1_101000110011;
      patterns[53664] = 29'b1_101000110100_000_1_101000110100;
      patterns[53665] = 29'b1_101000110100_001_1_110100101000;
      patterns[53666] = 29'b1_101000110100_010_1_010001101001;
      patterns[53667] = 29'b1_101000110100_011_0_100011010011;
      patterns[53668] = 29'b1_101000110100_100_0_110100011010;
      patterns[53669] = 29'b1_101000110100_101_0_011010001101;
      patterns[53670] = 29'b1_101000110100_110_1_101000110100;
      patterns[53671] = 29'b1_101000110100_111_1_101000110100;
      patterns[53672] = 29'b1_101000110101_000_1_101000110101;
      patterns[53673] = 29'b1_101000110101_001_1_110101101000;
      patterns[53674] = 29'b1_101000110101_010_1_010001101011;
      patterns[53675] = 29'b1_101000110101_011_0_100011010111;
      patterns[53676] = 29'b1_101000110101_100_1_110100011010;
      patterns[53677] = 29'b1_101000110101_101_0_111010001101;
      patterns[53678] = 29'b1_101000110101_110_1_101000110101;
      patterns[53679] = 29'b1_101000110101_111_1_101000110101;
      patterns[53680] = 29'b1_101000110110_000_1_101000110110;
      patterns[53681] = 29'b1_101000110110_001_1_110110101000;
      patterns[53682] = 29'b1_101000110110_010_1_010001101101;
      patterns[53683] = 29'b1_101000110110_011_0_100011011011;
      patterns[53684] = 29'b1_101000110110_100_0_110100011011;
      patterns[53685] = 29'b1_101000110110_101_1_011010001101;
      patterns[53686] = 29'b1_101000110110_110_1_101000110110;
      patterns[53687] = 29'b1_101000110110_111_1_101000110110;
      patterns[53688] = 29'b1_101000110111_000_1_101000110111;
      patterns[53689] = 29'b1_101000110111_001_1_110111101000;
      patterns[53690] = 29'b1_101000110111_010_1_010001101111;
      patterns[53691] = 29'b1_101000110111_011_0_100011011111;
      patterns[53692] = 29'b1_101000110111_100_1_110100011011;
      patterns[53693] = 29'b1_101000110111_101_1_111010001101;
      patterns[53694] = 29'b1_101000110111_110_1_101000110111;
      patterns[53695] = 29'b1_101000110111_111_1_101000110111;
      patterns[53696] = 29'b1_101000111000_000_1_101000111000;
      patterns[53697] = 29'b1_101000111000_001_1_111000101000;
      patterns[53698] = 29'b1_101000111000_010_1_010001110001;
      patterns[53699] = 29'b1_101000111000_011_0_100011100011;
      patterns[53700] = 29'b1_101000111000_100_0_110100011100;
      patterns[53701] = 29'b1_101000111000_101_0_011010001110;
      patterns[53702] = 29'b1_101000111000_110_1_101000111000;
      patterns[53703] = 29'b1_101000111000_111_1_101000111000;
      patterns[53704] = 29'b1_101000111001_000_1_101000111001;
      patterns[53705] = 29'b1_101000111001_001_1_111001101000;
      patterns[53706] = 29'b1_101000111001_010_1_010001110011;
      patterns[53707] = 29'b1_101000111001_011_0_100011100111;
      patterns[53708] = 29'b1_101000111001_100_1_110100011100;
      patterns[53709] = 29'b1_101000111001_101_0_111010001110;
      patterns[53710] = 29'b1_101000111001_110_1_101000111001;
      patterns[53711] = 29'b1_101000111001_111_1_101000111001;
      patterns[53712] = 29'b1_101000111010_000_1_101000111010;
      patterns[53713] = 29'b1_101000111010_001_1_111010101000;
      patterns[53714] = 29'b1_101000111010_010_1_010001110101;
      patterns[53715] = 29'b1_101000111010_011_0_100011101011;
      patterns[53716] = 29'b1_101000111010_100_0_110100011101;
      patterns[53717] = 29'b1_101000111010_101_1_011010001110;
      patterns[53718] = 29'b1_101000111010_110_1_101000111010;
      patterns[53719] = 29'b1_101000111010_111_1_101000111010;
      patterns[53720] = 29'b1_101000111011_000_1_101000111011;
      patterns[53721] = 29'b1_101000111011_001_1_111011101000;
      patterns[53722] = 29'b1_101000111011_010_1_010001110111;
      patterns[53723] = 29'b1_101000111011_011_0_100011101111;
      patterns[53724] = 29'b1_101000111011_100_1_110100011101;
      patterns[53725] = 29'b1_101000111011_101_1_111010001110;
      patterns[53726] = 29'b1_101000111011_110_1_101000111011;
      patterns[53727] = 29'b1_101000111011_111_1_101000111011;
      patterns[53728] = 29'b1_101000111100_000_1_101000111100;
      patterns[53729] = 29'b1_101000111100_001_1_111100101000;
      patterns[53730] = 29'b1_101000111100_010_1_010001111001;
      patterns[53731] = 29'b1_101000111100_011_0_100011110011;
      patterns[53732] = 29'b1_101000111100_100_0_110100011110;
      patterns[53733] = 29'b1_101000111100_101_0_011010001111;
      patterns[53734] = 29'b1_101000111100_110_1_101000111100;
      patterns[53735] = 29'b1_101000111100_111_1_101000111100;
      patterns[53736] = 29'b1_101000111101_000_1_101000111101;
      patterns[53737] = 29'b1_101000111101_001_1_111101101000;
      patterns[53738] = 29'b1_101000111101_010_1_010001111011;
      patterns[53739] = 29'b1_101000111101_011_0_100011110111;
      patterns[53740] = 29'b1_101000111101_100_1_110100011110;
      patterns[53741] = 29'b1_101000111101_101_0_111010001111;
      patterns[53742] = 29'b1_101000111101_110_1_101000111101;
      patterns[53743] = 29'b1_101000111101_111_1_101000111101;
      patterns[53744] = 29'b1_101000111110_000_1_101000111110;
      patterns[53745] = 29'b1_101000111110_001_1_111110101000;
      patterns[53746] = 29'b1_101000111110_010_1_010001111101;
      patterns[53747] = 29'b1_101000111110_011_0_100011111011;
      patterns[53748] = 29'b1_101000111110_100_0_110100011111;
      patterns[53749] = 29'b1_101000111110_101_1_011010001111;
      patterns[53750] = 29'b1_101000111110_110_1_101000111110;
      patterns[53751] = 29'b1_101000111110_111_1_101000111110;
      patterns[53752] = 29'b1_101000111111_000_1_101000111111;
      patterns[53753] = 29'b1_101000111111_001_1_111111101000;
      patterns[53754] = 29'b1_101000111111_010_1_010001111111;
      patterns[53755] = 29'b1_101000111111_011_0_100011111111;
      patterns[53756] = 29'b1_101000111111_100_1_110100011111;
      patterns[53757] = 29'b1_101000111111_101_1_111010001111;
      patterns[53758] = 29'b1_101000111111_110_1_101000111111;
      patterns[53759] = 29'b1_101000111111_111_1_101000111111;
      patterns[53760] = 29'b1_101001000000_000_1_101001000000;
      patterns[53761] = 29'b1_101001000000_001_1_000000101001;
      patterns[53762] = 29'b1_101001000000_010_1_010010000001;
      patterns[53763] = 29'b1_101001000000_011_0_100100000011;
      patterns[53764] = 29'b1_101001000000_100_0_110100100000;
      patterns[53765] = 29'b1_101001000000_101_0_011010010000;
      patterns[53766] = 29'b1_101001000000_110_1_101001000000;
      patterns[53767] = 29'b1_101001000000_111_1_101001000000;
      patterns[53768] = 29'b1_101001000001_000_1_101001000001;
      patterns[53769] = 29'b1_101001000001_001_1_000001101001;
      patterns[53770] = 29'b1_101001000001_010_1_010010000011;
      patterns[53771] = 29'b1_101001000001_011_0_100100000111;
      patterns[53772] = 29'b1_101001000001_100_1_110100100000;
      patterns[53773] = 29'b1_101001000001_101_0_111010010000;
      patterns[53774] = 29'b1_101001000001_110_1_101001000001;
      patterns[53775] = 29'b1_101001000001_111_1_101001000001;
      patterns[53776] = 29'b1_101001000010_000_1_101001000010;
      patterns[53777] = 29'b1_101001000010_001_1_000010101001;
      patterns[53778] = 29'b1_101001000010_010_1_010010000101;
      patterns[53779] = 29'b1_101001000010_011_0_100100001011;
      patterns[53780] = 29'b1_101001000010_100_0_110100100001;
      patterns[53781] = 29'b1_101001000010_101_1_011010010000;
      patterns[53782] = 29'b1_101001000010_110_1_101001000010;
      patterns[53783] = 29'b1_101001000010_111_1_101001000010;
      patterns[53784] = 29'b1_101001000011_000_1_101001000011;
      patterns[53785] = 29'b1_101001000011_001_1_000011101001;
      patterns[53786] = 29'b1_101001000011_010_1_010010000111;
      patterns[53787] = 29'b1_101001000011_011_0_100100001111;
      patterns[53788] = 29'b1_101001000011_100_1_110100100001;
      patterns[53789] = 29'b1_101001000011_101_1_111010010000;
      patterns[53790] = 29'b1_101001000011_110_1_101001000011;
      patterns[53791] = 29'b1_101001000011_111_1_101001000011;
      patterns[53792] = 29'b1_101001000100_000_1_101001000100;
      patterns[53793] = 29'b1_101001000100_001_1_000100101001;
      patterns[53794] = 29'b1_101001000100_010_1_010010001001;
      patterns[53795] = 29'b1_101001000100_011_0_100100010011;
      patterns[53796] = 29'b1_101001000100_100_0_110100100010;
      patterns[53797] = 29'b1_101001000100_101_0_011010010001;
      patterns[53798] = 29'b1_101001000100_110_1_101001000100;
      patterns[53799] = 29'b1_101001000100_111_1_101001000100;
      patterns[53800] = 29'b1_101001000101_000_1_101001000101;
      patterns[53801] = 29'b1_101001000101_001_1_000101101001;
      patterns[53802] = 29'b1_101001000101_010_1_010010001011;
      patterns[53803] = 29'b1_101001000101_011_0_100100010111;
      patterns[53804] = 29'b1_101001000101_100_1_110100100010;
      patterns[53805] = 29'b1_101001000101_101_0_111010010001;
      patterns[53806] = 29'b1_101001000101_110_1_101001000101;
      patterns[53807] = 29'b1_101001000101_111_1_101001000101;
      patterns[53808] = 29'b1_101001000110_000_1_101001000110;
      patterns[53809] = 29'b1_101001000110_001_1_000110101001;
      patterns[53810] = 29'b1_101001000110_010_1_010010001101;
      patterns[53811] = 29'b1_101001000110_011_0_100100011011;
      patterns[53812] = 29'b1_101001000110_100_0_110100100011;
      patterns[53813] = 29'b1_101001000110_101_1_011010010001;
      patterns[53814] = 29'b1_101001000110_110_1_101001000110;
      patterns[53815] = 29'b1_101001000110_111_1_101001000110;
      patterns[53816] = 29'b1_101001000111_000_1_101001000111;
      patterns[53817] = 29'b1_101001000111_001_1_000111101001;
      patterns[53818] = 29'b1_101001000111_010_1_010010001111;
      patterns[53819] = 29'b1_101001000111_011_0_100100011111;
      patterns[53820] = 29'b1_101001000111_100_1_110100100011;
      patterns[53821] = 29'b1_101001000111_101_1_111010010001;
      patterns[53822] = 29'b1_101001000111_110_1_101001000111;
      patterns[53823] = 29'b1_101001000111_111_1_101001000111;
      patterns[53824] = 29'b1_101001001000_000_1_101001001000;
      patterns[53825] = 29'b1_101001001000_001_1_001000101001;
      patterns[53826] = 29'b1_101001001000_010_1_010010010001;
      patterns[53827] = 29'b1_101001001000_011_0_100100100011;
      patterns[53828] = 29'b1_101001001000_100_0_110100100100;
      patterns[53829] = 29'b1_101001001000_101_0_011010010010;
      patterns[53830] = 29'b1_101001001000_110_1_101001001000;
      patterns[53831] = 29'b1_101001001000_111_1_101001001000;
      patterns[53832] = 29'b1_101001001001_000_1_101001001001;
      patterns[53833] = 29'b1_101001001001_001_1_001001101001;
      patterns[53834] = 29'b1_101001001001_010_1_010010010011;
      patterns[53835] = 29'b1_101001001001_011_0_100100100111;
      patterns[53836] = 29'b1_101001001001_100_1_110100100100;
      patterns[53837] = 29'b1_101001001001_101_0_111010010010;
      patterns[53838] = 29'b1_101001001001_110_1_101001001001;
      patterns[53839] = 29'b1_101001001001_111_1_101001001001;
      patterns[53840] = 29'b1_101001001010_000_1_101001001010;
      patterns[53841] = 29'b1_101001001010_001_1_001010101001;
      patterns[53842] = 29'b1_101001001010_010_1_010010010101;
      patterns[53843] = 29'b1_101001001010_011_0_100100101011;
      patterns[53844] = 29'b1_101001001010_100_0_110100100101;
      patterns[53845] = 29'b1_101001001010_101_1_011010010010;
      patterns[53846] = 29'b1_101001001010_110_1_101001001010;
      patterns[53847] = 29'b1_101001001010_111_1_101001001010;
      patterns[53848] = 29'b1_101001001011_000_1_101001001011;
      patterns[53849] = 29'b1_101001001011_001_1_001011101001;
      patterns[53850] = 29'b1_101001001011_010_1_010010010111;
      patterns[53851] = 29'b1_101001001011_011_0_100100101111;
      patterns[53852] = 29'b1_101001001011_100_1_110100100101;
      patterns[53853] = 29'b1_101001001011_101_1_111010010010;
      patterns[53854] = 29'b1_101001001011_110_1_101001001011;
      patterns[53855] = 29'b1_101001001011_111_1_101001001011;
      patterns[53856] = 29'b1_101001001100_000_1_101001001100;
      patterns[53857] = 29'b1_101001001100_001_1_001100101001;
      patterns[53858] = 29'b1_101001001100_010_1_010010011001;
      patterns[53859] = 29'b1_101001001100_011_0_100100110011;
      patterns[53860] = 29'b1_101001001100_100_0_110100100110;
      patterns[53861] = 29'b1_101001001100_101_0_011010010011;
      patterns[53862] = 29'b1_101001001100_110_1_101001001100;
      patterns[53863] = 29'b1_101001001100_111_1_101001001100;
      patterns[53864] = 29'b1_101001001101_000_1_101001001101;
      patterns[53865] = 29'b1_101001001101_001_1_001101101001;
      patterns[53866] = 29'b1_101001001101_010_1_010010011011;
      patterns[53867] = 29'b1_101001001101_011_0_100100110111;
      patterns[53868] = 29'b1_101001001101_100_1_110100100110;
      patterns[53869] = 29'b1_101001001101_101_0_111010010011;
      patterns[53870] = 29'b1_101001001101_110_1_101001001101;
      patterns[53871] = 29'b1_101001001101_111_1_101001001101;
      patterns[53872] = 29'b1_101001001110_000_1_101001001110;
      patterns[53873] = 29'b1_101001001110_001_1_001110101001;
      patterns[53874] = 29'b1_101001001110_010_1_010010011101;
      patterns[53875] = 29'b1_101001001110_011_0_100100111011;
      patterns[53876] = 29'b1_101001001110_100_0_110100100111;
      patterns[53877] = 29'b1_101001001110_101_1_011010010011;
      patterns[53878] = 29'b1_101001001110_110_1_101001001110;
      patterns[53879] = 29'b1_101001001110_111_1_101001001110;
      patterns[53880] = 29'b1_101001001111_000_1_101001001111;
      patterns[53881] = 29'b1_101001001111_001_1_001111101001;
      patterns[53882] = 29'b1_101001001111_010_1_010010011111;
      patterns[53883] = 29'b1_101001001111_011_0_100100111111;
      patterns[53884] = 29'b1_101001001111_100_1_110100100111;
      patterns[53885] = 29'b1_101001001111_101_1_111010010011;
      patterns[53886] = 29'b1_101001001111_110_1_101001001111;
      patterns[53887] = 29'b1_101001001111_111_1_101001001111;
      patterns[53888] = 29'b1_101001010000_000_1_101001010000;
      patterns[53889] = 29'b1_101001010000_001_1_010000101001;
      patterns[53890] = 29'b1_101001010000_010_1_010010100001;
      patterns[53891] = 29'b1_101001010000_011_0_100101000011;
      patterns[53892] = 29'b1_101001010000_100_0_110100101000;
      patterns[53893] = 29'b1_101001010000_101_0_011010010100;
      patterns[53894] = 29'b1_101001010000_110_1_101001010000;
      patterns[53895] = 29'b1_101001010000_111_1_101001010000;
      patterns[53896] = 29'b1_101001010001_000_1_101001010001;
      patterns[53897] = 29'b1_101001010001_001_1_010001101001;
      patterns[53898] = 29'b1_101001010001_010_1_010010100011;
      patterns[53899] = 29'b1_101001010001_011_0_100101000111;
      patterns[53900] = 29'b1_101001010001_100_1_110100101000;
      patterns[53901] = 29'b1_101001010001_101_0_111010010100;
      patterns[53902] = 29'b1_101001010001_110_1_101001010001;
      patterns[53903] = 29'b1_101001010001_111_1_101001010001;
      patterns[53904] = 29'b1_101001010010_000_1_101001010010;
      patterns[53905] = 29'b1_101001010010_001_1_010010101001;
      patterns[53906] = 29'b1_101001010010_010_1_010010100101;
      patterns[53907] = 29'b1_101001010010_011_0_100101001011;
      patterns[53908] = 29'b1_101001010010_100_0_110100101001;
      patterns[53909] = 29'b1_101001010010_101_1_011010010100;
      patterns[53910] = 29'b1_101001010010_110_1_101001010010;
      patterns[53911] = 29'b1_101001010010_111_1_101001010010;
      patterns[53912] = 29'b1_101001010011_000_1_101001010011;
      patterns[53913] = 29'b1_101001010011_001_1_010011101001;
      patterns[53914] = 29'b1_101001010011_010_1_010010100111;
      patterns[53915] = 29'b1_101001010011_011_0_100101001111;
      patterns[53916] = 29'b1_101001010011_100_1_110100101001;
      patterns[53917] = 29'b1_101001010011_101_1_111010010100;
      patterns[53918] = 29'b1_101001010011_110_1_101001010011;
      patterns[53919] = 29'b1_101001010011_111_1_101001010011;
      patterns[53920] = 29'b1_101001010100_000_1_101001010100;
      patterns[53921] = 29'b1_101001010100_001_1_010100101001;
      patterns[53922] = 29'b1_101001010100_010_1_010010101001;
      patterns[53923] = 29'b1_101001010100_011_0_100101010011;
      patterns[53924] = 29'b1_101001010100_100_0_110100101010;
      patterns[53925] = 29'b1_101001010100_101_0_011010010101;
      patterns[53926] = 29'b1_101001010100_110_1_101001010100;
      patterns[53927] = 29'b1_101001010100_111_1_101001010100;
      patterns[53928] = 29'b1_101001010101_000_1_101001010101;
      patterns[53929] = 29'b1_101001010101_001_1_010101101001;
      patterns[53930] = 29'b1_101001010101_010_1_010010101011;
      patterns[53931] = 29'b1_101001010101_011_0_100101010111;
      patterns[53932] = 29'b1_101001010101_100_1_110100101010;
      patterns[53933] = 29'b1_101001010101_101_0_111010010101;
      patterns[53934] = 29'b1_101001010101_110_1_101001010101;
      patterns[53935] = 29'b1_101001010101_111_1_101001010101;
      patterns[53936] = 29'b1_101001010110_000_1_101001010110;
      patterns[53937] = 29'b1_101001010110_001_1_010110101001;
      patterns[53938] = 29'b1_101001010110_010_1_010010101101;
      patterns[53939] = 29'b1_101001010110_011_0_100101011011;
      patterns[53940] = 29'b1_101001010110_100_0_110100101011;
      patterns[53941] = 29'b1_101001010110_101_1_011010010101;
      patterns[53942] = 29'b1_101001010110_110_1_101001010110;
      patterns[53943] = 29'b1_101001010110_111_1_101001010110;
      patterns[53944] = 29'b1_101001010111_000_1_101001010111;
      patterns[53945] = 29'b1_101001010111_001_1_010111101001;
      patterns[53946] = 29'b1_101001010111_010_1_010010101111;
      patterns[53947] = 29'b1_101001010111_011_0_100101011111;
      patterns[53948] = 29'b1_101001010111_100_1_110100101011;
      patterns[53949] = 29'b1_101001010111_101_1_111010010101;
      patterns[53950] = 29'b1_101001010111_110_1_101001010111;
      patterns[53951] = 29'b1_101001010111_111_1_101001010111;
      patterns[53952] = 29'b1_101001011000_000_1_101001011000;
      patterns[53953] = 29'b1_101001011000_001_1_011000101001;
      patterns[53954] = 29'b1_101001011000_010_1_010010110001;
      patterns[53955] = 29'b1_101001011000_011_0_100101100011;
      patterns[53956] = 29'b1_101001011000_100_0_110100101100;
      patterns[53957] = 29'b1_101001011000_101_0_011010010110;
      patterns[53958] = 29'b1_101001011000_110_1_101001011000;
      patterns[53959] = 29'b1_101001011000_111_1_101001011000;
      patterns[53960] = 29'b1_101001011001_000_1_101001011001;
      patterns[53961] = 29'b1_101001011001_001_1_011001101001;
      patterns[53962] = 29'b1_101001011001_010_1_010010110011;
      patterns[53963] = 29'b1_101001011001_011_0_100101100111;
      patterns[53964] = 29'b1_101001011001_100_1_110100101100;
      patterns[53965] = 29'b1_101001011001_101_0_111010010110;
      patterns[53966] = 29'b1_101001011001_110_1_101001011001;
      patterns[53967] = 29'b1_101001011001_111_1_101001011001;
      patterns[53968] = 29'b1_101001011010_000_1_101001011010;
      patterns[53969] = 29'b1_101001011010_001_1_011010101001;
      patterns[53970] = 29'b1_101001011010_010_1_010010110101;
      patterns[53971] = 29'b1_101001011010_011_0_100101101011;
      patterns[53972] = 29'b1_101001011010_100_0_110100101101;
      patterns[53973] = 29'b1_101001011010_101_1_011010010110;
      patterns[53974] = 29'b1_101001011010_110_1_101001011010;
      patterns[53975] = 29'b1_101001011010_111_1_101001011010;
      patterns[53976] = 29'b1_101001011011_000_1_101001011011;
      patterns[53977] = 29'b1_101001011011_001_1_011011101001;
      patterns[53978] = 29'b1_101001011011_010_1_010010110111;
      patterns[53979] = 29'b1_101001011011_011_0_100101101111;
      patterns[53980] = 29'b1_101001011011_100_1_110100101101;
      patterns[53981] = 29'b1_101001011011_101_1_111010010110;
      patterns[53982] = 29'b1_101001011011_110_1_101001011011;
      patterns[53983] = 29'b1_101001011011_111_1_101001011011;
      patterns[53984] = 29'b1_101001011100_000_1_101001011100;
      patterns[53985] = 29'b1_101001011100_001_1_011100101001;
      patterns[53986] = 29'b1_101001011100_010_1_010010111001;
      patterns[53987] = 29'b1_101001011100_011_0_100101110011;
      patterns[53988] = 29'b1_101001011100_100_0_110100101110;
      patterns[53989] = 29'b1_101001011100_101_0_011010010111;
      patterns[53990] = 29'b1_101001011100_110_1_101001011100;
      patterns[53991] = 29'b1_101001011100_111_1_101001011100;
      patterns[53992] = 29'b1_101001011101_000_1_101001011101;
      patterns[53993] = 29'b1_101001011101_001_1_011101101001;
      patterns[53994] = 29'b1_101001011101_010_1_010010111011;
      patterns[53995] = 29'b1_101001011101_011_0_100101110111;
      patterns[53996] = 29'b1_101001011101_100_1_110100101110;
      patterns[53997] = 29'b1_101001011101_101_0_111010010111;
      patterns[53998] = 29'b1_101001011101_110_1_101001011101;
      patterns[53999] = 29'b1_101001011101_111_1_101001011101;
      patterns[54000] = 29'b1_101001011110_000_1_101001011110;
      patterns[54001] = 29'b1_101001011110_001_1_011110101001;
      patterns[54002] = 29'b1_101001011110_010_1_010010111101;
      patterns[54003] = 29'b1_101001011110_011_0_100101111011;
      patterns[54004] = 29'b1_101001011110_100_0_110100101111;
      patterns[54005] = 29'b1_101001011110_101_1_011010010111;
      patterns[54006] = 29'b1_101001011110_110_1_101001011110;
      patterns[54007] = 29'b1_101001011110_111_1_101001011110;
      patterns[54008] = 29'b1_101001011111_000_1_101001011111;
      patterns[54009] = 29'b1_101001011111_001_1_011111101001;
      patterns[54010] = 29'b1_101001011111_010_1_010010111111;
      patterns[54011] = 29'b1_101001011111_011_0_100101111111;
      patterns[54012] = 29'b1_101001011111_100_1_110100101111;
      patterns[54013] = 29'b1_101001011111_101_1_111010010111;
      patterns[54014] = 29'b1_101001011111_110_1_101001011111;
      patterns[54015] = 29'b1_101001011111_111_1_101001011111;
      patterns[54016] = 29'b1_101001100000_000_1_101001100000;
      patterns[54017] = 29'b1_101001100000_001_1_100000101001;
      patterns[54018] = 29'b1_101001100000_010_1_010011000001;
      patterns[54019] = 29'b1_101001100000_011_0_100110000011;
      patterns[54020] = 29'b1_101001100000_100_0_110100110000;
      patterns[54021] = 29'b1_101001100000_101_0_011010011000;
      patterns[54022] = 29'b1_101001100000_110_1_101001100000;
      patterns[54023] = 29'b1_101001100000_111_1_101001100000;
      patterns[54024] = 29'b1_101001100001_000_1_101001100001;
      patterns[54025] = 29'b1_101001100001_001_1_100001101001;
      patterns[54026] = 29'b1_101001100001_010_1_010011000011;
      patterns[54027] = 29'b1_101001100001_011_0_100110000111;
      patterns[54028] = 29'b1_101001100001_100_1_110100110000;
      patterns[54029] = 29'b1_101001100001_101_0_111010011000;
      patterns[54030] = 29'b1_101001100001_110_1_101001100001;
      patterns[54031] = 29'b1_101001100001_111_1_101001100001;
      patterns[54032] = 29'b1_101001100010_000_1_101001100010;
      patterns[54033] = 29'b1_101001100010_001_1_100010101001;
      patterns[54034] = 29'b1_101001100010_010_1_010011000101;
      patterns[54035] = 29'b1_101001100010_011_0_100110001011;
      patterns[54036] = 29'b1_101001100010_100_0_110100110001;
      patterns[54037] = 29'b1_101001100010_101_1_011010011000;
      patterns[54038] = 29'b1_101001100010_110_1_101001100010;
      patterns[54039] = 29'b1_101001100010_111_1_101001100010;
      patterns[54040] = 29'b1_101001100011_000_1_101001100011;
      patterns[54041] = 29'b1_101001100011_001_1_100011101001;
      patterns[54042] = 29'b1_101001100011_010_1_010011000111;
      patterns[54043] = 29'b1_101001100011_011_0_100110001111;
      patterns[54044] = 29'b1_101001100011_100_1_110100110001;
      patterns[54045] = 29'b1_101001100011_101_1_111010011000;
      patterns[54046] = 29'b1_101001100011_110_1_101001100011;
      patterns[54047] = 29'b1_101001100011_111_1_101001100011;
      patterns[54048] = 29'b1_101001100100_000_1_101001100100;
      patterns[54049] = 29'b1_101001100100_001_1_100100101001;
      patterns[54050] = 29'b1_101001100100_010_1_010011001001;
      patterns[54051] = 29'b1_101001100100_011_0_100110010011;
      patterns[54052] = 29'b1_101001100100_100_0_110100110010;
      patterns[54053] = 29'b1_101001100100_101_0_011010011001;
      patterns[54054] = 29'b1_101001100100_110_1_101001100100;
      patterns[54055] = 29'b1_101001100100_111_1_101001100100;
      patterns[54056] = 29'b1_101001100101_000_1_101001100101;
      patterns[54057] = 29'b1_101001100101_001_1_100101101001;
      patterns[54058] = 29'b1_101001100101_010_1_010011001011;
      patterns[54059] = 29'b1_101001100101_011_0_100110010111;
      patterns[54060] = 29'b1_101001100101_100_1_110100110010;
      patterns[54061] = 29'b1_101001100101_101_0_111010011001;
      patterns[54062] = 29'b1_101001100101_110_1_101001100101;
      patterns[54063] = 29'b1_101001100101_111_1_101001100101;
      patterns[54064] = 29'b1_101001100110_000_1_101001100110;
      patterns[54065] = 29'b1_101001100110_001_1_100110101001;
      patterns[54066] = 29'b1_101001100110_010_1_010011001101;
      patterns[54067] = 29'b1_101001100110_011_0_100110011011;
      patterns[54068] = 29'b1_101001100110_100_0_110100110011;
      patterns[54069] = 29'b1_101001100110_101_1_011010011001;
      patterns[54070] = 29'b1_101001100110_110_1_101001100110;
      patterns[54071] = 29'b1_101001100110_111_1_101001100110;
      patterns[54072] = 29'b1_101001100111_000_1_101001100111;
      patterns[54073] = 29'b1_101001100111_001_1_100111101001;
      patterns[54074] = 29'b1_101001100111_010_1_010011001111;
      patterns[54075] = 29'b1_101001100111_011_0_100110011111;
      patterns[54076] = 29'b1_101001100111_100_1_110100110011;
      patterns[54077] = 29'b1_101001100111_101_1_111010011001;
      patterns[54078] = 29'b1_101001100111_110_1_101001100111;
      patterns[54079] = 29'b1_101001100111_111_1_101001100111;
      patterns[54080] = 29'b1_101001101000_000_1_101001101000;
      patterns[54081] = 29'b1_101001101000_001_1_101000101001;
      patterns[54082] = 29'b1_101001101000_010_1_010011010001;
      patterns[54083] = 29'b1_101001101000_011_0_100110100011;
      patterns[54084] = 29'b1_101001101000_100_0_110100110100;
      patterns[54085] = 29'b1_101001101000_101_0_011010011010;
      patterns[54086] = 29'b1_101001101000_110_1_101001101000;
      patterns[54087] = 29'b1_101001101000_111_1_101001101000;
      patterns[54088] = 29'b1_101001101001_000_1_101001101001;
      patterns[54089] = 29'b1_101001101001_001_1_101001101001;
      patterns[54090] = 29'b1_101001101001_010_1_010011010011;
      patterns[54091] = 29'b1_101001101001_011_0_100110100111;
      patterns[54092] = 29'b1_101001101001_100_1_110100110100;
      patterns[54093] = 29'b1_101001101001_101_0_111010011010;
      patterns[54094] = 29'b1_101001101001_110_1_101001101001;
      patterns[54095] = 29'b1_101001101001_111_1_101001101001;
      patterns[54096] = 29'b1_101001101010_000_1_101001101010;
      patterns[54097] = 29'b1_101001101010_001_1_101010101001;
      patterns[54098] = 29'b1_101001101010_010_1_010011010101;
      patterns[54099] = 29'b1_101001101010_011_0_100110101011;
      patterns[54100] = 29'b1_101001101010_100_0_110100110101;
      patterns[54101] = 29'b1_101001101010_101_1_011010011010;
      patterns[54102] = 29'b1_101001101010_110_1_101001101010;
      patterns[54103] = 29'b1_101001101010_111_1_101001101010;
      patterns[54104] = 29'b1_101001101011_000_1_101001101011;
      patterns[54105] = 29'b1_101001101011_001_1_101011101001;
      patterns[54106] = 29'b1_101001101011_010_1_010011010111;
      patterns[54107] = 29'b1_101001101011_011_0_100110101111;
      patterns[54108] = 29'b1_101001101011_100_1_110100110101;
      patterns[54109] = 29'b1_101001101011_101_1_111010011010;
      patterns[54110] = 29'b1_101001101011_110_1_101001101011;
      patterns[54111] = 29'b1_101001101011_111_1_101001101011;
      patterns[54112] = 29'b1_101001101100_000_1_101001101100;
      patterns[54113] = 29'b1_101001101100_001_1_101100101001;
      patterns[54114] = 29'b1_101001101100_010_1_010011011001;
      patterns[54115] = 29'b1_101001101100_011_0_100110110011;
      patterns[54116] = 29'b1_101001101100_100_0_110100110110;
      patterns[54117] = 29'b1_101001101100_101_0_011010011011;
      patterns[54118] = 29'b1_101001101100_110_1_101001101100;
      patterns[54119] = 29'b1_101001101100_111_1_101001101100;
      patterns[54120] = 29'b1_101001101101_000_1_101001101101;
      patterns[54121] = 29'b1_101001101101_001_1_101101101001;
      patterns[54122] = 29'b1_101001101101_010_1_010011011011;
      patterns[54123] = 29'b1_101001101101_011_0_100110110111;
      patterns[54124] = 29'b1_101001101101_100_1_110100110110;
      patterns[54125] = 29'b1_101001101101_101_0_111010011011;
      patterns[54126] = 29'b1_101001101101_110_1_101001101101;
      patterns[54127] = 29'b1_101001101101_111_1_101001101101;
      patterns[54128] = 29'b1_101001101110_000_1_101001101110;
      patterns[54129] = 29'b1_101001101110_001_1_101110101001;
      patterns[54130] = 29'b1_101001101110_010_1_010011011101;
      patterns[54131] = 29'b1_101001101110_011_0_100110111011;
      patterns[54132] = 29'b1_101001101110_100_0_110100110111;
      patterns[54133] = 29'b1_101001101110_101_1_011010011011;
      patterns[54134] = 29'b1_101001101110_110_1_101001101110;
      patterns[54135] = 29'b1_101001101110_111_1_101001101110;
      patterns[54136] = 29'b1_101001101111_000_1_101001101111;
      patterns[54137] = 29'b1_101001101111_001_1_101111101001;
      patterns[54138] = 29'b1_101001101111_010_1_010011011111;
      patterns[54139] = 29'b1_101001101111_011_0_100110111111;
      patterns[54140] = 29'b1_101001101111_100_1_110100110111;
      patterns[54141] = 29'b1_101001101111_101_1_111010011011;
      patterns[54142] = 29'b1_101001101111_110_1_101001101111;
      patterns[54143] = 29'b1_101001101111_111_1_101001101111;
      patterns[54144] = 29'b1_101001110000_000_1_101001110000;
      patterns[54145] = 29'b1_101001110000_001_1_110000101001;
      patterns[54146] = 29'b1_101001110000_010_1_010011100001;
      patterns[54147] = 29'b1_101001110000_011_0_100111000011;
      patterns[54148] = 29'b1_101001110000_100_0_110100111000;
      patterns[54149] = 29'b1_101001110000_101_0_011010011100;
      patterns[54150] = 29'b1_101001110000_110_1_101001110000;
      patterns[54151] = 29'b1_101001110000_111_1_101001110000;
      patterns[54152] = 29'b1_101001110001_000_1_101001110001;
      patterns[54153] = 29'b1_101001110001_001_1_110001101001;
      patterns[54154] = 29'b1_101001110001_010_1_010011100011;
      patterns[54155] = 29'b1_101001110001_011_0_100111000111;
      patterns[54156] = 29'b1_101001110001_100_1_110100111000;
      patterns[54157] = 29'b1_101001110001_101_0_111010011100;
      patterns[54158] = 29'b1_101001110001_110_1_101001110001;
      patterns[54159] = 29'b1_101001110001_111_1_101001110001;
      patterns[54160] = 29'b1_101001110010_000_1_101001110010;
      patterns[54161] = 29'b1_101001110010_001_1_110010101001;
      patterns[54162] = 29'b1_101001110010_010_1_010011100101;
      patterns[54163] = 29'b1_101001110010_011_0_100111001011;
      patterns[54164] = 29'b1_101001110010_100_0_110100111001;
      patterns[54165] = 29'b1_101001110010_101_1_011010011100;
      patterns[54166] = 29'b1_101001110010_110_1_101001110010;
      patterns[54167] = 29'b1_101001110010_111_1_101001110010;
      patterns[54168] = 29'b1_101001110011_000_1_101001110011;
      patterns[54169] = 29'b1_101001110011_001_1_110011101001;
      patterns[54170] = 29'b1_101001110011_010_1_010011100111;
      patterns[54171] = 29'b1_101001110011_011_0_100111001111;
      patterns[54172] = 29'b1_101001110011_100_1_110100111001;
      patterns[54173] = 29'b1_101001110011_101_1_111010011100;
      patterns[54174] = 29'b1_101001110011_110_1_101001110011;
      patterns[54175] = 29'b1_101001110011_111_1_101001110011;
      patterns[54176] = 29'b1_101001110100_000_1_101001110100;
      patterns[54177] = 29'b1_101001110100_001_1_110100101001;
      patterns[54178] = 29'b1_101001110100_010_1_010011101001;
      patterns[54179] = 29'b1_101001110100_011_0_100111010011;
      patterns[54180] = 29'b1_101001110100_100_0_110100111010;
      patterns[54181] = 29'b1_101001110100_101_0_011010011101;
      patterns[54182] = 29'b1_101001110100_110_1_101001110100;
      patterns[54183] = 29'b1_101001110100_111_1_101001110100;
      patterns[54184] = 29'b1_101001110101_000_1_101001110101;
      patterns[54185] = 29'b1_101001110101_001_1_110101101001;
      patterns[54186] = 29'b1_101001110101_010_1_010011101011;
      patterns[54187] = 29'b1_101001110101_011_0_100111010111;
      patterns[54188] = 29'b1_101001110101_100_1_110100111010;
      patterns[54189] = 29'b1_101001110101_101_0_111010011101;
      patterns[54190] = 29'b1_101001110101_110_1_101001110101;
      patterns[54191] = 29'b1_101001110101_111_1_101001110101;
      patterns[54192] = 29'b1_101001110110_000_1_101001110110;
      patterns[54193] = 29'b1_101001110110_001_1_110110101001;
      patterns[54194] = 29'b1_101001110110_010_1_010011101101;
      patterns[54195] = 29'b1_101001110110_011_0_100111011011;
      patterns[54196] = 29'b1_101001110110_100_0_110100111011;
      patterns[54197] = 29'b1_101001110110_101_1_011010011101;
      patterns[54198] = 29'b1_101001110110_110_1_101001110110;
      patterns[54199] = 29'b1_101001110110_111_1_101001110110;
      patterns[54200] = 29'b1_101001110111_000_1_101001110111;
      patterns[54201] = 29'b1_101001110111_001_1_110111101001;
      patterns[54202] = 29'b1_101001110111_010_1_010011101111;
      patterns[54203] = 29'b1_101001110111_011_0_100111011111;
      patterns[54204] = 29'b1_101001110111_100_1_110100111011;
      patterns[54205] = 29'b1_101001110111_101_1_111010011101;
      patterns[54206] = 29'b1_101001110111_110_1_101001110111;
      patterns[54207] = 29'b1_101001110111_111_1_101001110111;
      patterns[54208] = 29'b1_101001111000_000_1_101001111000;
      patterns[54209] = 29'b1_101001111000_001_1_111000101001;
      patterns[54210] = 29'b1_101001111000_010_1_010011110001;
      patterns[54211] = 29'b1_101001111000_011_0_100111100011;
      patterns[54212] = 29'b1_101001111000_100_0_110100111100;
      patterns[54213] = 29'b1_101001111000_101_0_011010011110;
      patterns[54214] = 29'b1_101001111000_110_1_101001111000;
      patterns[54215] = 29'b1_101001111000_111_1_101001111000;
      patterns[54216] = 29'b1_101001111001_000_1_101001111001;
      patterns[54217] = 29'b1_101001111001_001_1_111001101001;
      patterns[54218] = 29'b1_101001111001_010_1_010011110011;
      patterns[54219] = 29'b1_101001111001_011_0_100111100111;
      patterns[54220] = 29'b1_101001111001_100_1_110100111100;
      patterns[54221] = 29'b1_101001111001_101_0_111010011110;
      patterns[54222] = 29'b1_101001111001_110_1_101001111001;
      patterns[54223] = 29'b1_101001111001_111_1_101001111001;
      patterns[54224] = 29'b1_101001111010_000_1_101001111010;
      patterns[54225] = 29'b1_101001111010_001_1_111010101001;
      patterns[54226] = 29'b1_101001111010_010_1_010011110101;
      patterns[54227] = 29'b1_101001111010_011_0_100111101011;
      patterns[54228] = 29'b1_101001111010_100_0_110100111101;
      patterns[54229] = 29'b1_101001111010_101_1_011010011110;
      patterns[54230] = 29'b1_101001111010_110_1_101001111010;
      patterns[54231] = 29'b1_101001111010_111_1_101001111010;
      patterns[54232] = 29'b1_101001111011_000_1_101001111011;
      patterns[54233] = 29'b1_101001111011_001_1_111011101001;
      patterns[54234] = 29'b1_101001111011_010_1_010011110111;
      patterns[54235] = 29'b1_101001111011_011_0_100111101111;
      patterns[54236] = 29'b1_101001111011_100_1_110100111101;
      patterns[54237] = 29'b1_101001111011_101_1_111010011110;
      patterns[54238] = 29'b1_101001111011_110_1_101001111011;
      patterns[54239] = 29'b1_101001111011_111_1_101001111011;
      patterns[54240] = 29'b1_101001111100_000_1_101001111100;
      patterns[54241] = 29'b1_101001111100_001_1_111100101001;
      patterns[54242] = 29'b1_101001111100_010_1_010011111001;
      patterns[54243] = 29'b1_101001111100_011_0_100111110011;
      patterns[54244] = 29'b1_101001111100_100_0_110100111110;
      patterns[54245] = 29'b1_101001111100_101_0_011010011111;
      patterns[54246] = 29'b1_101001111100_110_1_101001111100;
      patterns[54247] = 29'b1_101001111100_111_1_101001111100;
      patterns[54248] = 29'b1_101001111101_000_1_101001111101;
      patterns[54249] = 29'b1_101001111101_001_1_111101101001;
      patterns[54250] = 29'b1_101001111101_010_1_010011111011;
      patterns[54251] = 29'b1_101001111101_011_0_100111110111;
      patterns[54252] = 29'b1_101001111101_100_1_110100111110;
      patterns[54253] = 29'b1_101001111101_101_0_111010011111;
      patterns[54254] = 29'b1_101001111101_110_1_101001111101;
      patterns[54255] = 29'b1_101001111101_111_1_101001111101;
      patterns[54256] = 29'b1_101001111110_000_1_101001111110;
      patterns[54257] = 29'b1_101001111110_001_1_111110101001;
      patterns[54258] = 29'b1_101001111110_010_1_010011111101;
      patterns[54259] = 29'b1_101001111110_011_0_100111111011;
      patterns[54260] = 29'b1_101001111110_100_0_110100111111;
      patterns[54261] = 29'b1_101001111110_101_1_011010011111;
      patterns[54262] = 29'b1_101001111110_110_1_101001111110;
      patterns[54263] = 29'b1_101001111110_111_1_101001111110;
      patterns[54264] = 29'b1_101001111111_000_1_101001111111;
      patterns[54265] = 29'b1_101001111111_001_1_111111101001;
      patterns[54266] = 29'b1_101001111111_010_1_010011111111;
      patterns[54267] = 29'b1_101001111111_011_0_100111111111;
      patterns[54268] = 29'b1_101001111111_100_1_110100111111;
      patterns[54269] = 29'b1_101001111111_101_1_111010011111;
      patterns[54270] = 29'b1_101001111111_110_1_101001111111;
      patterns[54271] = 29'b1_101001111111_111_1_101001111111;
      patterns[54272] = 29'b1_101010000000_000_1_101010000000;
      patterns[54273] = 29'b1_101010000000_001_1_000000101010;
      patterns[54274] = 29'b1_101010000000_010_1_010100000001;
      patterns[54275] = 29'b1_101010000000_011_0_101000000011;
      patterns[54276] = 29'b1_101010000000_100_0_110101000000;
      patterns[54277] = 29'b1_101010000000_101_0_011010100000;
      patterns[54278] = 29'b1_101010000000_110_1_101010000000;
      patterns[54279] = 29'b1_101010000000_111_1_101010000000;
      patterns[54280] = 29'b1_101010000001_000_1_101010000001;
      patterns[54281] = 29'b1_101010000001_001_1_000001101010;
      patterns[54282] = 29'b1_101010000001_010_1_010100000011;
      patterns[54283] = 29'b1_101010000001_011_0_101000000111;
      patterns[54284] = 29'b1_101010000001_100_1_110101000000;
      patterns[54285] = 29'b1_101010000001_101_0_111010100000;
      patterns[54286] = 29'b1_101010000001_110_1_101010000001;
      patterns[54287] = 29'b1_101010000001_111_1_101010000001;
      patterns[54288] = 29'b1_101010000010_000_1_101010000010;
      patterns[54289] = 29'b1_101010000010_001_1_000010101010;
      patterns[54290] = 29'b1_101010000010_010_1_010100000101;
      patterns[54291] = 29'b1_101010000010_011_0_101000001011;
      patterns[54292] = 29'b1_101010000010_100_0_110101000001;
      patterns[54293] = 29'b1_101010000010_101_1_011010100000;
      patterns[54294] = 29'b1_101010000010_110_1_101010000010;
      patterns[54295] = 29'b1_101010000010_111_1_101010000010;
      patterns[54296] = 29'b1_101010000011_000_1_101010000011;
      patterns[54297] = 29'b1_101010000011_001_1_000011101010;
      patterns[54298] = 29'b1_101010000011_010_1_010100000111;
      patterns[54299] = 29'b1_101010000011_011_0_101000001111;
      patterns[54300] = 29'b1_101010000011_100_1_110101000001;
      patterns[54301] = 29'b1_101010000011_101_1_111010100000;
      patterns[54302] = 29'b1_101010000011_110_1_101010000011;
      patterns[54303] = 29'b1_101010000011_111_1_101010000011;
      patterns[54304] = 29'b1_101010000100_000_1_101010000100;
      patterns[54305] = 29'b1_101010000100_001_1_000100101010;
      patterns[54306] = 29'b1_101010000100_010_1_010100001001;
      patterns[54307] = 29'b1_101010000100_011_0_101000010011;
      patterns[54308] = 29'b1_101010000100_100_0_110101000010;
      patterns[54309] = 29'b1_101010000100_101_0_011010100001;
      patterns[54310] = 29'b1_101010000100_110_1_101010000100;
      patterns[54311] = 29'b1_101010000100_111_1_101010000100;
      patterns[54312] = 29'b1_101010000101_000_1_101010000101;
      patterns[54313] = 29'b1_101010000101_001_1_000101101010;
      patterns[54314] = 29'b1_101010000101_010_1_010100001011;
      patterns[54315] = 29'b1_101010000101_011_0_101000010111;
      patterns[54316] = 29'b1_101010000101_100_1_110101000010;
      patterns[54317] = 29'b1_101010000101_101_0_111010100001;
      patterns[54318] = 29'b1_101010000101_110_1_101010000101;
      patterns[54319] = 29'b1_101010000101_111_1_101010000101;
      patterns[54320] = 29'b1_101010000110_000_1_101010000110;
      patterns[54321] = 29'b1_101010000110_001_1_000110101010;
      patterns[54322] = 29'b1_101010000110_010_1_010100001101;
      patterns[54323] = 29'b1_101010000110_011_0_101000011011;
      patterns[54324] = 29'b1_101010000110_100_0_110101000011;
      patterns[54325] = 29'b1_101010000110_101_1_011010100001;
      patterns[54326] = 29'b1_101010000110_110_1_101010000110;
      patterns[54327] = 29'b1_101010000110_111_1_101010000110;
      patterns[54328] = 29'b1_101010000111_000_1_101010000111;
      patterns[54329] = 29'b1_101010000111_001_1_000111101010;
      patterns[54330] = 29'b1_101010000111_010_1_010100001111;
      patterns[54331] = 29'b1_101010000111_011_0_101000011111;
      patterns[54332] = 29'b1_101010000111_100_1_110101000011;
      patterns[54333] = 29'b1_101010000111_101_1_111010100001;
      patterns[54334] = 29'b1_101010000111_110_1_101010000111;
      patterns[54335] = 29'b1_101010000111_111_1_101010000111;
      patterns[54336] = 29'b1_101010001000_000_1_101010001000;
      patterns[54337] = 29'b1_101010001000_001_1_001000101010;
      patterns[54338] = 29'b1_101010001000_010_1_010100010001;
      patterns[54339] = 29'b1_101010001000_011_0_101000100011;
      patterns[54340] = 29'b1_101010001000_100_0_110101000100;
      patterns[54341] = 29'b1_101010001000_101_0_011010100010;
      patterns[54342] = 29'b1_101010001000_110_1_101010001000;
      patterns[54343] = 29'b1_101010001000_111_1_101010001000;
      patterns[54344] = 29'b1_101010001001_000_1_101010001001;
      patterns[54345] = 29'b1_101010001001_001_1_001001101010;
      patterns[54346] = 29'b1_101010001001_010_1_010100010011;
      patterns[54347] = 29'b1_101010001001_011_0_101000100111;
      patterns[54348] = 29'b1_101010001001_100_1_110101000100;
      patterns[54349] = 29'b1_101010001001_101_0_111010100010;
      patterns[54350] = 29'b1_101010001001_110_1_101010001001;
      patterns[54351] = 29'b1_101010001001_111_1_101010001001;
      patterns[54352] = 29'b1_101010001010_000_1_101010001010;
      patterns[54353] = 29'b1_101010001010_001_1_001010101010;
      patterns[54354] = 29'b1_101010001010_010_1_010100010101;
      patterns[54355] = 29'b1_101010001010_011_0_101000101011;
      patterns[54356] = 29'b1_101010001010_100_0_110101000101;
      patterns[54357] = 29'b1_101010001010_101_1_011010100010;
      patterns[54358] = 29'b1_101010001010_110_1_101010001010;
      patterns[54359] = 29'b1_101010001010_111_1_101010001010;
      patterns[54360] = 29'b1_101010001011_000_1_101010001011;
      patterns[54361] = 29'b1_101010001011_001_1_001011101010;
      patterns[54362] = 29'b1_101010001011_010_1_010100010111;
      patterns[54363] = 29'b1_101010001011_011_0_101000101111;
      patterns[54364] = 29'b1_101010001011_100_1_110101000101;
      patterns[54365] = 29'b1_101010001011_101_1_111010100010;
      patterns[54366] = 29'b1_101010001011_110_1_101010001011;
      patterns[54367] = 29'b1_101010001011_111_1_101010001011;
      patterns[54368] = 29'b1_101010001100_000_1_101010001100;
      patterns[54369] = 29'b1_101010001100_001_1_001100101010;
      patterns[54370] = 29'b1_101010001100_010_1_010100011001;
      patterns[54371] = 29'b1_101010001100_011_0_101000110011;
      patterns[54372] = 29'b1_101010001100_100_0_110101000110;
      patterns[54373] = 29'b1_101010001100_101_0_011010100011;
      patterns[54374] = 29'b1_101010001100_110_1_101010001100;
      patterns[54375] = 29'b1_101010001100_111_1_101010001100;
      patterns[54376] = 29'b1_101010001101_000_1_101010001101;
      patterns[54377] = 29'b1_101010001101_001_1_001101101010;
      patterns[54378] = 29'b1_101010001101_010_1_010100011011;
      patterns[54379] = 29'b1_101010001101_011_0_101000110111;
      patterns[54380] = 29'b1_101010001101_100_1_110101000110;
      patterns[54381] = 29'b1_101010001101_101_0_111010100011;
      patterns[54382] = 29'b1_101010001101_110_1_101010001101;
      patterns[54383] = 29'b1_101010001101_111_1_101010001101;
      patterns[54384] = 29'b1_101010001110_000_1_101010001110;
      patterns[54385] = 29'b1_101010001110_001_1_001110101010;
      patterns[54386] = 29'b1_101010001110_010_1_010100011101;
      patterns[54387] = 29'b1_101010001110_011_0_101000111011;
      patterns[54388] = 29'b1_101010001110_100_0_110101000111;
      patterns[54389] = 29'b1_101010001110_101_1_011010100011;
      patterns[54390] = 29'b1_101010001110_110_1_101010001110;
      patterns[54391] = 29'b1_101010001110_111_1_101010001110;
      patterns[54392] = 29'b1_101010001111_000_1_101010001111;
      patterns[54393] = 29'b1_101010001111_001_1_001111101010;
      patterns[54394] = 29'b1_101010001111_010_1_010100011111;
      patterns[54395] = 29'b1_101010001111_011_0_101000111111;
      patterns[54396] = 29'b1_101010001111_100_1_110101000111;
      patterns[54397] = 29'b1_101010001111_101_1_111010100011;
      patterns[54398] = 29'b1_101010001111_110_1_101010001111;
      patterns[54399] = 29'b1_101010001111_111_1_101010001111;
      patterns[54400] = 29'b1_101010010000_000_1_101010010000;
      patterns[54401] = 29'b1_101010010000_001_1_010000101010;
      patterns[54402] = 29'b1_101010010000_010_1_010100100001;
      patterns[54403] = 29'b1_101010010000_011_0_101001000011;
      patterns[54404] = 29'b1_101010010000_100_0_110101001000;
      patterns[54405] = 29'b1_101010010000_101_0_011010100100;
      patterns[54406] = 29'b1_101010010000_110_1_101010010000;
      patterns[54407] = 29'b1_101010010000_111_1_101010010000;
      patterns[54408] = 29'b1_101010010001_000_1_101010010001;
      patterns[54409] = 29'b1_101010010001_001_1_010001101010;
      patterns[54410] = 29'b1_101010010001_010_1_010100100011;
      patterns[54411] = 29'b1_101010010001_011_0_101001000111;
      patterns[54412] = 29'b1_101010010001_100_1_110101001000;
      patterns[54413] = 29'b1_101010010001_101_0_111010100100;
      patterns[54414] = 29'b1_101010010001_110_1_101010010001;
      patterns[54415] = 29'b1_101010010001_111_1_101010010001;
      patterns[54416] = 29'b1_101010010010_000_1_101010010010;
      patterns[54417] = 29'b1_101010010010_001_1_010010101010;
      patterns[54418] = 29'b1_101010010010_010_1_010100100101;
      patterns[54419] = 29'b1_101010010010_011_0_101001001011;
      patterns[54420] = 29'b1_101010010010_100_0_110101001001;
      patterns[54421] = 29'b1_101010010010_101_1_011010100100;
      patterns[54422] = 29'b1_101010010010_110_1_101010010010;
      patterns[54423] = 29'b1_101010010010_111_1_101010010010;
      patterns[54424] = 29'b1_101010010011_000_1_101010010011;
      patterns[54425] = 29'b1_101010010011_001_1_010011101010;
      patterns[54426] = 29'b1_101010010011_010_1_010100100111;
      patterns[54427] = 29'b1_101010010011_011_0_101001001111;
      patterns[54428] = 29'b1_101010010011_100_1_110101001001;
      patterns[54429] = 29'b1_101010010011_101_1_111010100100;
      patterns[54430] = 29'b1_101010010011_110_1_101010010011;
      patterns[54431] = 29'b1_101010010011_111_1_101010010011;
      patterns[54432] = 29'b1_101010010100_000_1_101010010100;
      patterns[54433] = 29'b1_101010010100_001_1_010100101010;
      patterns[54434] = 29'b1_101010010100_010_1_010100101001;
      patterns[54435] = 29'b1_101010010100_011_0_101001010011;
      patterns[54436] = 29'b1_101010010100_100_0_110101001010;
      patterns[54437] = 29'b1_101010010100_101_0_011010100101;
      patterns[54438] = 29'b1_101010010100_110_1_101010010100;
      patterns[54439] = 29'b1_101010010100_111_1_101010010100;
      patterns[54440] = 29'b1_101010010101_000_1_101010010101;
      patterns[54441] = 29'b1_101010010101_001_1_010101101010;
      patterns[54442] = 29'b1_101010010101_010_1_010100101011;
      patterns[54443] = 29'b1_101010010101_011_0_101001010111;
      patterns[54444] = 29'b1_101010010101_100_1_110101001010;
      patterns[54445] = 29'b1_101010010101_101_0_111010100101;
      patterns[54446] = 29'b1_101010010101_110_1_101010010101;
      patterns[54447] = 29'b1_101010010101_111_1_101010010101;
      patterns[54448] = 29'b1_101010010110_000_1_101010010110;
      patterns[54449] = 29'b1_101010010110_001_1_010110101010;
      patterns[54450] = 29'b1_101010010110_010_1_010100101101;
      patterns[54451] = 29'b1_101010010110_011_0_101001011011;
      patterns[54452] = 29'b1_101010010110_100_0_110101001011;
      patterns[54453] = 29'b1_101010010110_101_1_011010100101;
      patterns[54454] = 29'b1_101010010110_110_1_101010010110;
      patterns[54455] = 29'b1_101010010110_111_1_101010010110;
      patterns[54456] = 29'b1_101010010111_000_1_101010010111;
      patterns[54457] = 29'b1_101010010111_001_1_010111101010;
      patterns[54458] = 29'b1_101010010111_010_1_010100101111;
      patterns[54459] = 29'b1_101010010111_011_0_101001011111;
      patterns[54460] = 29'b1_101010010111_100_1_110101001011;
      patterns[54461] = 29'b1_101010010111_101_1_111010100101;
      patterns[54462] = 29'b1_101010010111_110_1_101010010111;
      patterns[54463] = 29'b1_101010010111_111_1_101010010111;
      patterns[54464] = 29'b1_101010011000_000_1_101010011000;
      patterns[54465] = 29'b1_101010011000_001_1_011000101010;
      patterns[54466] = 29'b1_101010011000_010_1_010100110001;
      patterns[54467] = 29'b1_101010011000_011_0_101001100011;
      patterns[54468] = 29'b1_101010011000_100_0_110101001100;
      patterns[54469] = 29'b1_101010011000_101_0_011010100110;
      patterns[54470] = 29'b1_101010011000_110_1_101010011000;
      patterns[54471] = 29'b1_101010011000_111_1_101010011000;
      patterns[54472] = 29'b1_101010011001_000_1_101010011001;
      patterns[54473] = 29'b1_101010011001_001_1_011001101010;
      patterns[54474] = 29'b1_101010011001_010_1_010100110011;
      patterns[54475] = 29'b1_101010011001_011_0_101001100111;
      patterns[54476] = 29'b1_101010011001_100_1_110101001100;
      patterns[54477] = 29'b1_101010011001_101_0_111010100110;
      patterns[54478] = 29'b1_101010011001_110_1_101010011001;
      patterns[54479] = 29'b1_101010011001_111_1_101010011001;
      patterns[54480] = 29'b1_101010011010_000_1_101010011010;
      patterns[54481] = 29'b1_101010011010_001_1_011010101010;
      patterns[54482] = 29'b1_101010011010_010_1_010100110101;
      patterns[54483] = 29'b1_101010011010_011_0_101001101011;
      patterns[54484] = 29'b1_101010011010_100_0_110101001101;
      patterns[54485] = 29'b1_101010011010_101_1_011010100110;
      patterns[54486] = 29'b1_101010011010_110_1_101010011010;
      patterns[54487] = 29'b1_101010011010_111_1_101010011010;
      patterns[54488] = 29'b1_101010011011_000_1_101010011011;
      patterns[54489] = 29'b1_101010011011_001_1_011011101010;
      patterns[54490] = 29'b1_101010011011_010_1_010100110111;
      patterns[54491] = 29'b1_101010011011_011_0_101001101111;
      patterns[54492] = 29'b1_101010011011_100_1_110101001101;
      patterns[54493] = 29'b1_101010011011_101_1_111010100110;
      patterns[54494] = 29'b1_101010011011_110_1_101010011011;
      patterns[54495] = 29'b1_101010011011_111_1_101010011011;
      patterns[54496] = 29'b1_101010011100_000_1_101010011100;
      patterns[54497] = 29'b1_101010011100_001_1_011100101010;
      patterns[54498] = 29'b1_101010011100_010_1_010100111001;
      patterns[54499] = 29'b1_101010011100_011_0_101001110011;
      patterns[54500] = 29'b1_101010011100_100_0_110101001110;
      patterns[54501] = 29'b1_101010011100_101_0_011010100111;
      patterns[54502] = 29'b1_101010011100_110_1_101010011100;
      patterns[54503] = 29'b1_101010011100_111_1_101010011100;
      patterns[54504] = 29'b1_101010011101_000_1_101010011101;
      patterns[54505] = 29'b1_101010011101_001_1_011101101010;
      patterns[54506] = 29'b1_101010011101_010_1_010100111011;
      patterns[54507] = 29'b1_101010011101_011_0_101001110111;
      patterns[54508] = 29'b1_101010011101_100_1_110101001110;
      patterns[54509] = 29'b1_101010011101_101_0_111010100111;
      patterns[54510] = 29'b1_101010011101_110_1_101010011101;
      patterns[54511] = 29'b1_101010011101_111_1_101010011101;
      patterns[54512] = 29'b1_101010011110_000_1_101010011110;
      patterns[54513] = 29'b1_101010011110_001_1_011110101010;
      patterns[54514] = 29'b1_101010011110_010_1_010100111101;
      patterns[54515] = 29'b1_101010011110_011_0_101001111011;
      patterns[54516] = 29'b1_101010011110_100_0_110101001111;
      patterns[54517] = 29'b1_101010011110_101_1_011010100111;
      patterns[54518] = 29'b1_101010011110_110_1_101010011110;
      patterns[54519] = 29'b1_101010011110_111_1_101010011110;
      patterns[54520] = 29'b1_101010011111_000_1_101010011111;
      patterns[54521] = 29'b1_101010011111_001_1_011111101010;
      patterns[54522] = 29'b1_101010011111_010_1_010100111111;
      patterns[54523] = 29'b1_101010011111_011_0_101001111111;
      patterns[54524] = 29'b1_101010011111_100_1_110101001111;
      patterns[54525] = 29'b1_101010011111_101_1_111010100111;
      patterns[54526] = 29'b1_101010011111_110_1_101010011111;
      patterns[54527] = 29'b1_101010011111_111_1_101010011111;
      patterns[54528] = 29'b1_101010100000_000_1_101010100000;
      patterns[54529] = 29'b1_101010100000_001_1_100000101010;
      patterns[54530] = 29'b1_101010100000_010_1_010101000001;
      patterns[54531] = 29'b1_101010100000_011_0_101010000011;
      patterns[54532] = 29'b1_101010100000_100_0_110101010000;
      patterns[54533] = 29'b1_101010100000_101_0_011010101000;
      patterns[54534] = 29'b1_101010100000_110_1_101010100000;
      patterns[54535] = 29'b1_101010100000_111_1_101010100000;
      patterns[54536] = 29'b1_101010100001_000_1_101010100001;
      patterns[54537] = 29'b1_101010100001_001_1_100001101010;
      patterns[54538] = 29'b1_101010100001_010_1_010101000011;
      patterns[54539] = 29'b1_101010100001_011_0_101010000111;
      patterns[54540] = 29'b1_101010100001_100_1_110101010000;
      patterns[54541] = 29'b1_101010100001_101_0_111010101000;
      patterns[54542] = 29'b1_101010100001_110_1_101010100001;
      patterns[54543] = 29'b1_101010100001_111_1_101010100001;
      patterns[54544] = 29'b1_101010100010_000_1_101010100010;
      patterns[54545] = 29'b1_101010100010_001_1_100010101010;
      patterns[54546] = 29'b1_101010100010_010_1_010101000101;
      patterns[54547] = 29'b1_101010100010_011_0_101010001011;
      patterns[54548] = 29'b1_101010100010_100_0_110101010001;
      patterns[54549] = 29'b1_101010100010_101_1_011010101000;
      patterns[54550] = 29'b1_101010100010_110_1_101010100010;
      patterns[54551] = 29'b1_101010100010_111_1_101010100010;
      patterns[54552] = 29'b1_101010100011_000_1_101010100011;
      patterns[54553] = 29'b1_101010100011_001_1_100011101010;
      patterns[54554] = 29'b1_101010100011_010_1_010101000111;
      patterns[54555] = 29'b1_101010100011_011_0_101010001111;
      patterns[54556] = 29'b1_101010100011_100_1_110101010001;
      patterns[54557] = 29'b1_101010100011_101_1_111010101000;
      patterns[54558] = 29'b1_101010100011_110_1_101010100011;
      patterns[54559] = 29'b1_101010100011_111_1_101010100011;
      patterns[54560] = 29'b1_101010100100_000_1_101010100100;
      patterns[54561] = 29'b1_101010100100_001_1_100100101010;
      patterns[54562] = 29'b1_101010100100_010_1_010101001001;
      patterns[54563] = 29'b1_101010100100_011_0_101010010011;
      patterns[54564] = 29'b1_101010100100_100_0_110101010010;
      patterns[54565] = 29'b1_101010100100_101_0_011010101001;
      patterns[54566] = 29'b1_101010100100_110_1_101010100100;
      patterns[54567] = 29'b1_101010100100_111_1_101010100100;
      patterns[54568] = 29'b1_101010100101_000_1_101010100101;
      patterns[54569] = 29'b1_101010100101_001_1_100101101010;
      patterns[54570] = 29'b1_101010100101_010_1_010101001011;
      patterns[54571] = 29'b1_101010100101_011_0_101010010111;
      patterns[54572] = 29'b1_101010100101_100_1_110101010010;
      patterns[54573] = 29'b1_101010100101_101_0_111010101001;
      patterns[54574] = 29'b1_101010100101_110_1_101010100101;
      patterns[54575] = 29'b1_101010100101_111_1_101010100101;
      patterns[54576] = 29'b1_101010100110_000_1_101010100110;
      patterns[54577] = 29'b1_101010100110_001_1_100110101010;
      patterns[54578] = 29'b1_101010100110_010_1_010101001101;
      patterns[54579] = 29'b1_101010100110_011_0_101010011011;
      patterns[54580] = 29'b1_101010100110_100_0_110101010011;
      patterns[54581] = 29'b1_101010100110_101_1_011010101001;
      patterns[54582] = 29'b1_101010100110_110_1_101010100110;
      patterns[54583] = 29'b1_101010100110_111_1_101010100110;
      patterns[54584] = 29'b1_101010100111_000_1_101010100111;
      patterns[54585] = 29'b1_101010100111_001_1_100111101010;
      patterns[54586] = 29'b1_101010100111_010_1_010101001111;
      patterns[54587] = 29'b1_101010100111_011_0_101010011111;
      patterns[54588] = 29'b1_101010100111_100_1_110101010011;
      patterns[54589] = 29'b1_101010100111_101_1_111010101001;
      patterns[54590] = 29'b1_101010100111_110_1_101010100111;
      patterns[54591] = 29'b1_101010100111_111_1_101010100111;
      patterns[54592] = 29'b1_101010101000_000_1_101010101000;
      patterns[54593] = 29'b1_101010101000_001_1_101000101010;
      patterns[54594] = 29'b1_101010101000_010_1_010101010001;
      patterns[54595] = 29'b1_101010101000_011_0_101010100011;
      patterns[54596] = 29'b1_101010101000_100_0_110101010100;
      patterns[54597] = 29'b1_101010101000_101_0_011010101010;
      patterns[54598] = 29'b1_101010101000_110_1_101010101000;
      patterns[54599] = 29'b1_101010101000_111_1_101010101000;
      patterns[54600] = 29'b1_101010101001_000_1_101010101001;
      patterns[54601] = 29'b1_101010101001_001_1_101001101010;
      patterns[54602] = 29'b1_101010101001_010_1_010101010011;
      patterns[54603] = 29'b1_101010101001_011_0_101010100111;
      patterns[54604] = 29'b1_101010101001_100_1_110101010100;
      patterns[54605] = 29'b1_101010101001_101_0_111010101010;
      patterns[54606] = 29'b1_101010101001_110_1_101010101001;
      patterns[54607] = 29'b1_101010101001_111_1_101010101001;
      patterns[54608] = 29'b1_101010101010_000_1_101010101010;
      patterns[54609] = 29'b1_101010101010_001_1_101010101010;
      patterns[54610] = 29'b1_101010101010_010_1_010101010101;
      patterns[54611] = 29'b1_101010101010_011_0_101010101011;
      patterns[54612] = 29'b1_101010101010_100_0_110101010101;
      patterns[54613] = 29'b1_101010101010_101_1_011010101010;
      patterns[54614] = 29'b1_101010101010_110_1_101010101010;
      patterns[54615] = 29'b1_101010101010_111_1_101010101010;
      patterns[54616] = 29'b1_101010101011_000_1_101010101011;
      patterns[54617] = 29'b1_101010101011_001_1_101011101010;
      patterns[54618] = 29'b1_101010101011_010_1_010101010111;
      patterns[54619] = 29'b1_101010101011_011_0_101010101111;
      patterns[54620] = 29'b1_101010101011_100_1_110101010101;
      patterns[54621] = 29'b1_101010101011_101_1_111010101010;
      patterns[54622] = 29'b1_101010101011_110_1_101010101011;
      patterns[54623] = 29'b1_101010101011_111_1_101010101011;
      patterns[54624] = 29'b1_101010101100_000_1_101010101100;
      patterns[54625] = 29'b1_101010101100_001_1_101100101010;
      patterns[54626] = 29'b1_101010101100_010_1_010101011001;
      patterns[54627] = 29'b1_101010101100_011_0_101010110011;
      patterns[54628] = 29'b1_101010101100_100_0_110101010110;
      patterns[54629] = 29'b1_101010101100_101_0_011010101011;
      patterns[54630] = 29'b1_101010101100_110_1_101010101100;
      patterns[54631] = 29'b1_101010101100_111_1_101010101100;
      patterns[54632] = 29'b1_101010101101_000_1_101010101101;
      patterns[54633] = 29'b1_101010101101_001_1_101101101010;
      patterns[54634] = 29'b1_101010101101_010_1_010101011011;
      patterns[54635] = 29'b1_101010101101_011_0_101010110111;
      patterns[54636] = 29'b1_101010101101_100_1_110101010110;
      patterns[54637] = 29'b1_101010101101_101_0_111010101011;
      patterns[54638] = 29'b1_101010101101_110_1_101010101101;
      patterns[54639] = 29'b1_101010101101_111_1_101010101101;
      patterns[54640] = 29'b1_101010101110_000_1_101010101110;
      patterns[54641] = 29'b1_101010101110_001_1_101110101010;
      patterns[54642] = 29'b1_101010101110_010_1_010101011101;
      patterns[54643] = 29'b1_101010101110_011_0_101010111011;
      patterns[54644] = 29'b1_101010101110_100_0_110101010111;
      patterns[54645] = 29'b1_101010101110_101_1_011010101011;
      patterns[54646] = 29'b1_101010101110_110_1_101010101110;
      patterns[54647] = 29'b1_101010101110_111_1_101010101110;
      patterns[54648] = 29'b1_101010101111_000_1_101010101111;
      patterns[54649] = 29'b1_101010101111_001_1_101111101010;
      patterns[54650] = 29'b1_101010101111_010_1_010101011111;
      patterns[54651] = 29'b1_101010101111_011_0_101010111111;
      patterns[54652] = 29'b1_101010101111_100_1_110101010111;
      patterns[54653] = 29'b1_101010101111_101_1_111010101011;
      patterns[54654] = 29'b1_101010101111_110_1_101010101111;
      patterns[54655] = 29'b1_101010101111_111_1_101010101111;
      patterns[54656] = 29'b1_101010110000_000_1_101010110000;
      patterns[54657] = 29'b1_101010110000_001_1_110000101010;
      patterns[54658] = 29'b1_101010110000_010_1_010101100001;
      patterns[54659] = 29'b1_101010110000_011_0_101011000011;
      patterns[54660] = 29'b1_101010110000_100_0_110101011000;
      patterns[54661] = 29'b1_101010110000_101_0_011010101100;
      patterns[54662] = 29'b1_101010110000_110_1_101010110000;
      patterns[54663] = 29'b1_101010110000_111_1_101010110000;
      patterns[54664] = 29'b1_101010110001_000_1_101010110001;
      patterns[54665] = 29'b1_101010110001_001_1_110001101010;
      patterns[54666] = 29'b1_101010110001_010_1_010101100011;
      patterns[54667] = 29'b1_101010110001_011_0_101011000111;
      patterns[54668] = 29'b1_101010110001_100_1_110101011000;
      patterns[54669] = 29'b1_101010110001_101_0_111010101100;
      patterns[54670] = 29'b1_101010110001_110_1_101010110001;
      patterns[54671] = 29'b1_101010110001_111_1_101010110001;
      patterns[54672] = 29'b1_101010110010_000_1_101010110010;
      patterns[54673] = 29'b1_101010110010_001_1_110010101010;
      patterns[54674] = 29'b1_101010110010_010_1_010101100101;
      patterns[54675] = 29'b1_101010110010_011_0_101011001011;
      patterns[54676] = 29'b1_101010110010_100_0_110101011001;
      patterns[54677] = 29'b1_101010110010_101_1_011010101100;
      patterns[54678] = 29'b1_101010110010_110_1_101010110010;
      patterns[54679] = 29'b1_101010110010_111_1_101010110010;
      patterns[54680] = 29'b1_101010110011_000_1_101010110011;
      patterns[54681] = 29'b1_101010110011_001_1_110011101010;
      patterns[54682] = 29'b1_101010110011_010_1_010101100111;
      patterns[54683] = 29'b1_101010110011_011_0_101011001111;
      patterns[54684] = 29'b1_101010110011_100_1_110101011001;
      patterns[54685] = 29'b1_101010110011_101_1_111010101100;
      patterns[54686] = 29'b1_101010110011_110_1_101010110011;
      patterns[54687] = 29'b1_101010110011_111_1_101010110011;
      patterns[54688] = 29'b1_101010110100_000_1_101010110100;
      patterns[54689] = 29'b1_101010110100_001_1_110100101010;
      patterns[54690] = 29'b1_101010110100_010_1_010101101001;
      patterns[54691] = 29'b1_101010110100_011_0_101011010011;
      patterns[54692] = 29'b1_101010110100_100_0_110101011010;
      patterns[54693] = 29'b1_101010110100_101_0_011010101101;
      patterns[54694] = 29'b1_101010110100_110_1_101010110100;
      patterns[54695] = 29'b1_101010110100_111_1_101010110100;
      patterns[54696] = 29'b1_101010110101_000_1_101010110101;
      patterns[54697] = 29'b1_101010110101_001_1_110101101010;
      patterns[54698] = 29'b1_101010110101_010_1_010101101011;
      patterns[54699] = 29'b1_101010110101_011_0_101011010111;
      patterns[54700] = 29'b1_101010110101_100_1_110101011010;
      patterns[54701] = 29'b1_101010110101_101_0_111010101101;
      patterns[54702] = 29'b1_101010110101_110_1_101010110101;
      patterns[54703] = 29'b1_101010110101_111_1_101010110101;
      patterns[54704] = 29'b1_101010110110_000_1_101010110110;
      patterns[54705] = 29'b1_101010110110_001_1_110110101010;
      patterns[54706] = 29'b1_101010110110_010_1_010101101101;
      patterns[54707] = 29'b1_101010110110_011_0_101011011011;
      patterns[54708] = 29'b1_101010110110_100_0_110101011011;
      patterns[54709] = 29'b1_101010110110_101_1_011010101101;
      patterns[54710] = 29'b1_101010110110_110_1_101010110110;
      patterns[54711] = 29'b1_101010110110_111_1_101010110110;
      patterns[54712] = 29'b1_101010110111_000_1_101010110111;
      patterns[54713] = 29'b1_101010110111_001_1_110111101010;
      patterns[54714] = 29'b1_101010110111_010_1_010101101111;
      patterns[54715] = 29'b1_101010110111_011_0_101011011111;
      patterns[54716] = 29'b1_101010110111_100_1_110101011011;
      patterns[54717] = 29'b1_101010110111_101_1_111010101101;
      patterns[54718] = 29'b1_101010110111_110_1_101010110111;
      patterns[54719] = 29'b1_101010110111_111_1_101010110111;
      patterns[54720] = 29'b1_101010111000_000_1_101010111000;
      patterns[54721] = 29'b1_101010111000_001_1_111000101010;
      patterns[54722] = 29'b1_101010111000_010_1_010101110001;
      patterns[54723] = 29'b1_101010111000_011_0_101011100011;
      patterns[54724] = 29'b1_101010111000_100_0_110101011100;
      patterns[54725] = 29'b1_101010111000_101_0_011010101110;
      patterns[54726] = 29'b1_101010111000_110_1_101010111000;
      patterns[54727] = 29'b1_101010111000_111_1_101010111000;
      patterns[54728] = 29'b1_101010111001_000_1_101010111001;
      patterns[54729] = 29'b1_101010111001_001_1_111001101010;
      patterns[54730] = 29'b1_101010111001_010_1_010101110011;
      patterns[54731] = 29'b1_101010111001_011_0_101011100111;
      patterns[54732] = 29'b1_101010111001_100_1_110101011100;
      patterns[54733] = 29'b1_101010111001_101_0_111010101110;
      patterns[54734] = 29'b1_101010111001_110_1_101010111001;
      patterns[54735] = 29'b1_101010111001_111_1_101010111001;
      patterns[54736] = 29'b1_101010111010_000_1_101010111010;
      patterns[54737] = 29'b1_101010111010_001_1_111010101010;
      patterns[54738] = 29'b1_101010111010_010_1_010101110101;
      patterns[54739] = 29'b1_101010111010_011_0_101011101011;
      patterns[54740] = 29'b1_101010111010_100_0_110101011101;
      patterns[54741] = 29'b1_101010111010_101_1_011010101110;
      patterns[54742] = 29'b1_101010111010_110_1_101010111010;
      patterns[54743] = 29'b1_101010111010_111_1_101010111010;
      patterns[54744] = 29'b1_101010111011_000_1_101010111011;
      patterns[54745] = 29'b1_101010111011_001_1_111011101010;
      patterns[54746] = 29'b1_101010111011_010_1_010101110111;
      patterns[54747] = 29'b1_101010111011_011_0_101011101111;
      patterns[54748] = 29'b1_101010111011_100_1_110101011101;
      patterns[54749] = 29'b1_101010111011_101_1_111010101110;
      patterns[54750] = 29'b1_101010111011_110_1_101010111011;
      patterns[54751] = 29'b1_101010111011_111_1_101010111011;
      patterns[54752] = 29'b1_101010111100_000_1_101010111100;
      patterns[54753] = 29'b1_101010111100_001_1_111100101010;
      patterns[54754] = 29'b1_101010111100_010_1_010101111001;
      patterns[54755] = 29'b1_101010111100_011_0_101011110011;
      patterns[54756] = 29'b1_101010111100_100_0_110101011110;
      patterns[54757] = 29'b1_101010111100_101_0_011010101111;
      patterns[54758] = 29'b1_101010111100_110_1_101010111100;
      patterns[54759] = 29'b1_101010111100_111_1_101010111100;
      patterns[54760] = 29'b1_101010111101_000_1_101010111101;
      patterns[54761] = 29'b1_101010111101_001_1_111101101010;
      patterns[54762] = 29'b1_101010111101_010_1_010101111011;
      patterns[54763] = 29'b1_101010111101_011_0_101011110111;
      patterns[54764] = 29'b1_101010111101_100_1_110101011110;
      patterns[54765] = 29'b1_101010111101_101_0_111010101111;
      patterns[54766] = 29'b1_101010111101_110_1_101010111101;
      patterns[54767] = 29'b1_101010111101_111_1_101010111101;
      patterns[54768] = 29'b1_101010111110_000_1_101010111110;
      patterns[54769] = 29'b1_101010111110_001_1_111110101010;
      patterns[54770] = 29'b1_101010111110_010_1_010101111101;
      patterns[54771] = 29'b1_101010111110_011_0_101011111011;
      patterns[54772] = 29'b1_101010111110_100_0_110101011111;
      patterns[54773] = 29'b1_101010111110_101_1_011010101111;
      patterns[54774] = 29'b1_101010111110_110_1_101010111110;
      patterns[54775] = 29'b1_101010111110_111_1_101010111110;
      patterns[54776] = 29'b1_101010111111_000_1_101010111111;
      patterns[54777] = 29'b1_101010111111_001_1_111111101010;
      patterns[54778] = 29'b1_101010111111_010_1_010101111111;
      patterns[54779] = 29'b1_101010111111_011_0_101011111111;
      patterns[54780] = 29'b1_101010111111_100_1_110101011111;
      patterns[54781] = 29'b1_101010111111_101_1_111010101111;
      patterns[54782] = 29'b1_101010111111_110_1_101010111111;
      patterns[54783] = 29'b1_101010111111_111_1_101010111111;
      patterns[54784] = 29'b1_101011000000_000_1_101011000000;
      patterns[54785] = 29'b1_101011000000_001_1_000000101011;
      patterns[54786] = 29'b1_101011000000_010_1_010110000001;
      patterns[54787] = 29'b1_101011000000_011_0_101100000011;
      patterns[54788] = 29'b1_101011000000_100_0_110101100000;
      patterns[54789] = 29'b1_101011000000_101_0_011010110000;
      patterns[54790] = 29'b1_101011000000_110_1_101011000000;
      patterns[54791] = 29'b1_101011000000_111_1_101011000000;
      patterns[54792] = 29'b1_101011000001_000_1_101011000001;
      patterns[54793] = 29'b1_101011000001_001_1_000001101011;
      patterns[54794] = 29'b1_101011000001_010_1_010110000011;
      patterns[54795] = 29'b1_101011000001_011_0_101100000111;
      patterns[54796] = 29'b1_101011000001_100_1_110101100000;
      patterns[54797] = 29'b1_101011000001_101_0_111010110000;
      patterns[54798] = 29'b1_101011000001_110_1_101011000001;
      patterns[54799] = 29'b1_101011000001_111_1_101011000001;
      patterns[54800] = 29'b1_101011000010_000_1_101011000010;
      patterns[54801] = 29'b1_101011000010_001_1_000010101011;
      patterns[54802] = 29'b1_101011000010_010_1_010110000101;
      patterns[54803] = 29'b1_101011000010_011_0_101100001011;
      patterns[54804] = 29'b1_101011000010_100_0_110101100001;
      patterns[54805] = 29'b1_101011000010_101_1_011010110000;
      patterns[54806] = 29'b1_101011000010_110_1_101011000010;
      patterns[54807] = 29'b1_101011000010_111_1_101011000010;
      patterns[54808] = 29'b1_101011000011_000_1_101011000011;
      patterns[54809] = 29'b1_101011000011_001_1_000011101011;
      patterns[54810] = 29'b1_101011000011_010_1_010110000111;
      patterns[54811] = 29'b1_101011000011_011_0_101100001111;
      patterns[54812] = 29'b1_101011000011_100_1_110101100001;
      patterns[54813] = 29'b1_101011000011_101_1_111010110000;
      patterns[54814] = 29'b1_101011000011_110_1_101011000011;
      patterns[54815] = 29'b1_101011000011_111_1_101011000011;
      patterns[54816] = 29'b1_101011000100_000_1_101011000100;
      patterns[54817] = 29'b1_101011000100_001_1_000100101011;
      patterns[54818] = 29'b1_101011000100_010_1_010110001001;
      patterns[54819] = 29'b1_101011000100_011_0_101100010011;
      patterns[54820] = 29'b1_101011000100_100_0_110101100010;
      patterns[54821] = 29'b1_101011000100_101_0_011010110001;
      patterns[54822] = 29'b1_101011000100_110_1_101011000100;
      patterns[54823] = 29'b1_101011000100_111_1_101011000100;
      patterns[54824] = 29'b1_101011000101_000_1_101011000101;
      patterns[54825] = 29'b1_101011000101_001_1_000101101011;
      patterns[54826] = 29'b1_101011000101_010_1_010110001011;
      patterns[54827] = 29'b1_101011000101_011_0_101100010111;
      patterns[54828] = 29'b1_101011000101_100_1_110101100010;
      patterns[54829] = 29'b1_101011000101_101_0_111010110001;
      patterns[54830] = 29'b1_101011000101_110_1_101011000101;
      patterns[54831] = 29'b1_101011000101_111_1_101011000101;
      patterns[54832] = 29'b1_101011000110_000_1_101011000110;
      patterns[54833] = 29'b1_101011000110_001_1_000110101011;
      patterns[54834] = 29'b1_101011000110_010_1_010110001101;
      patterns[54835] = 29'b1_101011000110_011_0_101100011011;
      patterns[54836] = 29'b1_101011000110_100_0_110101100011;
      patterns[54837] = 29'b1_101011000110_101_1_011010110001;
      patterns[54838] = 29'b1_101011000110_110_1_101011000110;
      patterns[54839] = 29'b1_101011000110_111_1_101011000110;
      patterns[54840] = 29'b1_101011000111_000_1_101011000111;
      patterns[54841] = 29'b1_101011000111_001_1_000111101011;
      patterns[54842] = 29'b1_101011000111_010_1_010110001111;
      patterns[54843] = 29'b1_101011000111_011_0_101100011111;
      patterns[54844] = 29'b1_101011000111_100_1_110101100011;
      patterns[54845] = 29'b1_101011000111_101_1_111010110001;
      patterns[54846] = 29'b1_101011000111_110_1_101011000111;
      patterns[54847] = 29'b1_101011000111_111_1_101011000111;
      patterns[54848] = 29'b1_101011001000_000_1_101011001000;
      patterns[54849] = 29'b1_101011001000_001_1_001000101011;
      patterns[54850] = 29'b1_101011001000_010_1_010110010001;
      patterns[54851] = 29'b1_101011001000_011_0_101100100011;
      patterns[54852] = 29'b1_101011001000_100_0_110101100100;
      patterns[54853] = 29'b1_101011001000_101_0_011010110010;
      patterns[54854] = 29'b1_101011001000_110_1_101011001000;
      patterns[54855] = 29'b1_101011001000_111_1_101011001000;
      patterns[54856] = 29'b1_101011001001_000_1_101011001001;
      patterns[54857] = 29'b1_101011001001_001_1_001001101011;
      patterns[54858] = 29'b1_101011001001_010_1_010110010011;
      patterns[54859] = 29'b1_101011001001_011_0_101100100111;
      patterns[54860] = 29'b1_101011001001_100_1_110101100100;
      patterns[54861] = 29'b1_101011001001_101_0_111010110010;
      patterns[54862] = 29'b1_101011001001_110_1_101011001001;
      patterns[54863] = 29'b1_101011001001_111_1_101011001001;
      patterns[54864] = 29'b1_101011001010_000_1_101011001010;
      patterns[54865] = 29'b1_101011001010_001_1_001010101011;
      patterns[54866] = 29'b1_101011001010_010_1_010110010101;
      patterns[54867] = 29'b1_101011001010_011_0_101100101011;
      patterns[54868] = 29'b1_101011001010_100_0_110101100101;
      patterns[54869] = 29'b1_101011001010_101_1_011010110010;
      patterns[54870] = 29'b1_101011001010_110_1_101011001010;
      patterns[54871] = 29'b1_101011001010_111_1_101011001010;
      patterns[54872] = 29'b1_101011001011_000_1_101011001011;
      patterns[54873] = 29'b1_101011001011_001_1_001011101011;
      patterns[54874] = 29'b1_101011001011_010_1_010110010111;
      patterns[54875] = 29'b1_101011001011_011_0_101100101111;
      patterns[54876] = 29'b1_101011001011_100_1_110101100101;
      patterns[54877] = 29'b1_101011001011_101_1_111010110010;
      patterns[54878] = 29'b1_101011001011_110_1_101011001011;
      patterns[54879] = 29'b1_101011001011_111_1_101011001011;
      patterns[54880] = 29'b1_101011001100_000_1_101011001100;
      patterns[54881] = 29'b1_101011001100_001_1_001100101011;
      patterns[54882] = 29'b1_101011001100_010_1_010110011001;
      patterns[54883] = 29'b1_101011001100_011_0_101100110011;
      patterns[54884] = 29'b1_101011001100_100_0_110101100110;
      patterns[54885] = 29'b1_101011001100_101_0_011010110011;
      patterns[54886] = 29'b1_101011001100_110_1_101011001100;
      patterns[54887] = 29'b1_101011001100_111_1_101011001100;
      patterns[54888] = 29'b1_101011001101_000_1_101011001101;
      patterns[54889] = 29'b1_101011001101_001_1_001101101011;
      patterns[54890] = 29'b1_101011001101_010_1_010110011011;
      patterns[54891] = 29'b1_101011001101_011_0_101100110111;
      patterns[54892] = 29'b1_101011001101_100_1_110101100110;
      patterns[54893] = 29'b1_101011001101_101_0_111010110011;
      patterns[54894] = 29'b1_101011001101_110_1_101011001101;
      patterns[54895] = 29'b1_101011001101_111_1_101011001101;
      patterns[54896] = 29'b1_101011001110_000_1_101011001110;
      patterns[54897] = 29'b1_101011001110_001_1_001110101011;
      patterns[54898] = 29'b1_101011001110_010_1_010110011101;
      patterns[54899] = 29'b1_101011001110_011_0_101100111011;
      patterns[54900] = 29'b1_101011001110_100_0_110101100111;
      patterns[54901] = 29'b1_101011001110_101_1_011010110011;
      patterns[54902] = 29'b1_101011001110_110_1_101011001110;
      patterns[54903] = 29'b1_101011001110_111_1_101011001110;
      patterns[54904] = 29'b1_101011001111_000_1_101011001111;
      patterns[54905] = 29'b1_101011001111_001_1_001111101011;
      patterns[54906] = 29'b1_101011001111_010_1_010110011111;
      patterns[54907] = 29'b1_101011001111_011_0_101100111111;
      patterns[54908] = 29'b1_101011001111_100_1_110101100111;
      patterns[54909] = 29'b1_101011001111_101_1_111010110011;
      patterns[54910] = 29'b1_101011001111_110_1_101011001111;
      patterns[54911] = 29'b1_101011001111_111_1_101011001111;
      patterns[54912] = 29'b1_101011010000_000_1_101011010000;
      patterns[54913] = 29'b1_101011010000_001_1_010000101011;
      patterns[54914] = 29'b1_101011010000_010_1_010110100001;
      patterns[54915] = 29'b1_101011010000_011_0_101101000011;
      patterns[54916] = 29'b1_101011010000_100_0_110101101000;
      patterns[54917] = 29'b1_101011010000_101_0_011010110100;
      patterns[54918] = 29'b1_101011010000_110_1_101011010000;
      patterns[54919] = 29'b1_101011010000_111_1_101011010000;
      patterns[54920] = 29'b1_101011010001_000_1_101011010001;
      patterns[54921] = 29'b1_101011010001_001_1_010001101011;
      patterns[54922] = 29'b1_101011010001_010_1_010110100011;
      patterns[54923] = 29'b1_101011010001_011_0_101101000111;
      patterns[54924] = 29'b1_101011010001_100_1_110101101000;
      patterns[54925] = 29'b1_101011010001_101_0_111010110100;
      patterns[54926] = 29'b1_101011010001_110_1_101011010001;
      patterns[54927] = 29'b1_101011010001_111_1_101011010001;
      patterns[54928] = 29'b1_101011010010_000_1_101011010010;
      patterns[54929] = 29'b1_101011010010_001_1_010010101011;
      patterns[54930] = 29'b1_101011010010_010_1_010110100101;
      patterns[54931] = 29'b1_101011010010_011_0_101101001011;
      patterns[54932] = 29'b1_101011010010_100_0_110101101001;
      patterns[54933] = 29'b1_101011010010_101_1_011010110100;
      patterns[54934] = 29'b1_101011010010_110_1_101011010010;
      patterns[54935] = 29'b1_101011010010_111_1_101011010010;
      patterns[54936] = 29'b1_101011010011_000_1_101011010011;
      patterns[54937] = 29'b1_101011010011_001_1_010011101011;
      patterns[54938] = 29'b1_101011010011_010_1_010110100111;
      patterns[54939] = 29'b1_101011010011_011_0_101101001111;
      patterns[54940] = 29'b1_101011010011_100_1_110101101001;
      patterns[54941] = 29'b1_101011010011_101_1_111010110100;
      patterns[54942] = 29'b1_101011010011_110_1_101011010011;
      patterns[54943] = 29'b1_101011010011_111_1_101011010011;
      patterns[54944] = 29'b1_101011010100_000_1_101011010100;
      patterns[54945] = 29'b1_101011010100_001_1_010100101011;
      patterns[54946] = 29'b1_101011010100_010_1_010110101001;
      patterns[54947] = 29'b1_101011010100_011_0_101101010011;
      patterns[54948] = 29'b1_101011010100_100_0_110101101010;
      patterns[54949] = 29'b1_101011010100_101_0_011010110101;
      patterns[54950] = 29'b1_101011010100_110_1_101011010100;
      patterns[54951] = 29'b1_101011010100_111_1_101011010100;
      patterns[54952] = 29'b1_101011010101_000_1_101011010101;
      patterns[54953] = 29'b1_101011010101_001_1_010101101011;
      patterns[54954] = 29'b1_101011010101_010_1_010110101011;
      patterns[54955] = 29'b1_101011010101_011_0_101101010111;
      patterns[54956] = 29'b1_101011010101_100_1_110101101010;
      patterns[54957] = 29'b1_101011010101_101_0_111010110101;
      patterns[54958] = 29'b1_101011010101_110_1_101011010101;
      patterns[54959] = 29'b1_101011010101_111_1_101011010101;
      patterns[54960] = 29'b1_101011010110_000_1_101011010110;
      patterns[54961] = 29'b1_101011010110_001_1_010110101011;
      patterns[54962] = 29'b1_101011010110_010_1_010110101101;
      patterns[54963] = 29'b1_101011010110_011_0_101101011011;
      patterns[54964] = 29'b1_101011010110_100_0_110101101011;
      patterns[54965] = 29'b1_101011010110_101_1_011010110101;
      patterns[54966] = 29'b1_101011010110_110_1_101011010110;
      patterns[54967] = 29'b1_101011010110_111_1_101011010110;
      patterns[54968] = 29'b1_101011010111_000_1_101011010111;
      patterns[54969] = 29'b1_101011010111_001_1_010111101011;
      patterns[54970] = 29'b1_101011010111_010_1_010110101111;
      patterns[54971] = 29'b1_101011010111_011_0_101101011111;
      patterns[54972] = 29'b1_101011010111_100_1_110101101011;
      patterns[54973] = 29'b1_101011010111_101_1_111010110101;
      patterns[54974] = 29'b1_101011010111_110_1_101011010111;
      patterns[54975] = 29'b1_101011010111_111_1_101011010111;
      patterns[54976] = 29'b1_101011011000_000_1_101011011000;
      patterns[54977] = 29'b1_101011011000_001_1_011000101011;
      patterns[54978] = 29'b1_101011011000_010_1_010110110001;
      patterns[54979] = 29'b1_101011011000_011_0_101101100011;
      patterns[54980] = 29'b1_101011011000_100_0_110101101100;
      patterns[54981] = 29'b1_101011011000_101_0_011010110110;
      patterns[54982] = 29'b1_101011011000_110_1_101011011000;
      patterns[54983] = 29'b1_101011011000_111_1_101011011000;
      patterns[54984] = 29'b1_101011011001_000_1_101011011001;
      patterns[54985] = 29'b1_101011011001_001_1_011001101011;
      patterns[54986] = 29'b1_101011011001_010_1_010110110011;
      patterns[54987] = 29'b1_101011011001_011_0_101101100111;
      patterns[54988] = 29'b1_101011011001_100_1_110101101100;
      patterns[54989] = 29'b1_101011011001_101_0_111010110110;
      patterns[54990] = 29'b1_101011011001_110_1_101011011001;
      patterns[54991] = 29'b1_101011011001_111_1_101011011001;
      patterns[54992] = 29'b1_101011011010_000_1_101011011010;
      patterns[54993] = 29'b1_101011011010_001_1_011010101011;
      patterns[54994] = 29'b1_101011011010_010_1_010110110101;
      patterns[54995] = 29'b1_101011011010_011_0_101101101011;
      patterns[54996] = 29'b1_101011011010_100_0_110101101101;
      patterns[54997] = 29'b1_101011011010_101_1_011010110110;
      patterns[54998] = 29'b1_101011011010_110_1_101011011010;
      patterns[54999] = 29'b1_101011011010_111_1_101011011010;
      patterns[55000] = 29'b1_101011011011_000_1_101011011011;
      patterns[55001] = 29'b1_101011011011_001_1_011011101011;
      patterns[55002] = 29'b1_101011011011_010_1_010110110111;
      patterns[55003] = 29'b1_101011011011_011_0_101101101111;
      patterns[55004] = 29'b1_101011011011_100_1_110101101101;
      patterns[55005] = 29'b1_101011011011_101_1_111010110110;
      patterns[55006] = 29'b1_101011011011_110_1_101011011011;
      patterns[55007] = 29'b1_101011011011_111_1_101011011011;
      patterns[55008] = 29'b1_101011011100_000_1_101011011100;
      patterns[55009] = 29'b1_101011011100_001_1_011100101011;
      patterns[55010] = 29'b1_101011011100_010_1_010110111001;
      patterns[55011] = 29'b1_101011011100_011_0_101101110011;
      patterns[55012] = 29'b1_101011011100_100_0_110101101110;
      patterns[55013] = 29'b1_101011011100_101_0_011010110111;
      patterns[55014] = 29'b1_101011011100_110_1_101011011100;
      patterns[55015] = 29'b1_101011011100_111_1_101011011100;
      patterns[55016] = 29'b1_101011011101_000_1_101011011101;
      patterns[55017] = 29'b1_101011011101_001_1_011101101011;
      patterns[55018] = 29'b1_101011011101_010_1_010110111011;
      patterns[55019] = 29'b1_101011011101_011_0_101101110111;
      patterns[55020] = 29'b1_101011011101_100_1_110101101110;
      patterns[55021] = 29'b1_101011011101_101_0_111010110111;
      patterns[55022] = 29'b1_101011011101_110_1_101011011101;
      patterns[55023] = 29'b1_101011011101_111_1_101011011101;
      patterns[55024] = 29'b1_101011011110_000_1_101011011110;
      patterns[55025] = 29'b1_101011011110_001_1_011110101011;
      patterns[55026] = 29'b1_101011011110_010_1_010110111101;
      patterns[55027] = 29'b1_101011011110_011_0_101101111011;
      patterns[55028] = 29'b1_101011011110_100_0_110101101111;
      patterns[55029] = 29'b1_101011011110_101_1_011010110111;
      patterns[55030] = 29'b1_101011011110_110_1_101011011110;
      patterns[55031] = 29'b1_101011011110_111_1_101011011110;
      patterns[55032] = 29'b1_101011011111_000_1_101011011111;
      patterns[55033] = 29'b1_101011011111_001_1_011111101011;
      patterns[55034] = 29'b1_101011011111_010_1_010110111111;
      patterns[55035] = 29'b1_101011011111_011_0_101101111111;
      patterns[55036] = 29'b1_101011011111_100_1_110101101111;
      patterns[55037] = 29'b1_101011011111_101_1_111010110111;
      patterns[55038] = 29'b1_101011011111_110_1_101011011111;
      patterns[55039] = 29'b1_101011011111_111_1_101011011111;
      patterns[55040] = 29'b1_101011100000_000_1_101011100000;
      patterns[55041] = 29'b1_101011100000_001_1_100000101011;
      patterns[55042] = 29'b1_101011100000_010_1_010111000001;
      patterns[55043] = 29'b1_101011100000_011_0_101110000011;
      patterns[55044] = 29'b1_101011100000_100_0_110101110000;
      patterns[55045] = 29'b1_101011100000_101_0_011010111000;
      patterns[55046] = 29'b1_101011100000_110_1_101011100000;
      patterns[55047] = 29'b1_101011100000_111_1_101011100000;
      patterns[55048] = 29'b1_101011100001_000_1_101011100001;
      patterns[55049] = 29'b1_101011100001_001_1_100001101011;
      patterns[55050] = 29'b1_101011100001_010_1_010111000011;
      patterns[55051] = 29'b1_101011100001_011_0_101110000111;
      patterns[55052] = 29'b1_101011100001_100_1_110101110000;
      patterns[55053] = 29'b1_101011100001_101_0_111010111000;
      patterns[55054] = 29'b1_101011100001_110_1_101011100001;
      patterns[55055] = 29'b1_101011100001_111_1_101011100001;
      patterns[55056] = 29'b1_101011100010_000_1_101011100010;
      patterns[55057] = 29'b1_101011100010_001_1_100010101011;
      patterns[55058] = 29'b1_101011100010_010_1_010111000101;
      patterns[55059] = 29'b1_101011100010_011_0_101110001011;
      patterns[55060] = 29'b1_101011100010_100_0_110101110001;
      patterns[55061] = 29'b1_101011100010_101_1_011010111000;
      patterns[55062] = 29'b1_101011100010_110_1_101011100010;
      patterns[55063] = 29'b1_101011100010_111_1_101011100010;
      patterns[55064] = 29'b1_101011100011_000_1_101011100011;
      patterns[55065] = 29'b1_101011100011_001_1_100011101011;
      patterns[55066] = 29'b1_101011100011_010_1_010111000111;
      patterns[55067] = 29'b1_101011100011_011_0_101110001111;
      patterns[55068] = 29'b1_101011100011_100_1_110101110001;
      patterns[55069] = 29'b1_101011100011_101_1_111010111000;
      patterns[55070] = 29'b1_101011100011_110_1_101011100011;
      patterns[55071] = 29'b1_101011100011_111_1_101011100011;
      patterns[55072] = 29'b1_101011100100_000_1_101011100100;
      patterns[55073] = 29'b1_101011100100_001_1_100100101011;
      patterns[55074] = 29'b1_101011100100_010_1_010111001001;
      patterns[55075] = 29'b1_101011100100_011_0_101110010011;
      patterns[55076] = 29'b1_101011100100_100_0_110101110010;
      patterns[55077] = 29'b1_101011100100_101_0_011010111001;
      patterns[55078] = 29'b1_101011100100_110_1_101011100100;
      patterns[55079] = 29'b1_101011100100_111_1_101011100100;
      patterns[55080] = 29'b1_101011100101_000_1_101011100101;
      patterns[55081] = 29'b1_101011100101_001_1_100101101011;
      patterns[55082] = 29'b1_101011100101_010_1_010111001011;
      patterns[55083] = 29'b1_101011100101_011_0_101110010111;
      patterns[55084] = 29'b1_101011100101_100_1_110101110010;
      patterns[55085] = 29'b1_101011100101_101_0_111010111001;
      patterns[55086] = 29'b1_101011100101_110_1_101011100101;
      patterns[55087] = 29'b1_101011100101_111_1_101011100101;
      patterns[55088] = 29'b1_101011100110_000_1_101011100110;
      patterns[55089] = 29'b1_101011100110_001_1_100110101011;
      patterns[55090] = 29'b1_101011100110_010_1_010111001101;
      patterns[55091] = 29'b1_101011100110_011_0_101110011011;
      patterns[55092] = 29'b1_101011100110_100_0_110101110011;
      patterns[55093] = 29'b1_101011100110_101_1_011010111001;
      patterns[55094] = 29'b1_101011100110_110_1_101011100110;
      patterns[55095] = 29'b1_101011100110_111_1_101011100110;
      patterns[55096] = 29'b1_101011100111_000_1_101011100111;
      patterns[55097] = 29'b1_101011100111_001_1_100111101011;
      patterns[55098] = 29'b1_101011100111_010_1_010111001111;
      patterns[55099] = 29'b1_101011100111_011_0_101110011111;
      patterns[55100] = 29'b1_101011100111_100_1_110101110011;
      patterns[55101] = 29'b1_101011100111_101_1_111010111001;
      patterns[55102] = 29'b1_101011100111_110_1_101011100111;
      patterns[55103] = 29'b1_101011100111_111_1_101011100111;
      patterns[55104] = 29'b1_101011101000_000_1_101011101000;
      patterns[55105] = 29'b1_101011101000_001_1_101000101011;
      patterns[55106] = 29'b1_101011101000_010_1_010111010001;
      patterns[55107] = 29'b1_101011101000_011_0_101110100011;
      patterns[55108] = 29'b1_101011101000_100_0_110101110100;
      patterns[55109] = 29'b1_101011101000_101_0_011010111010;
      patterns[55110] = 29'b1_101011101000_110_1_101011101000;
      patterns[55111] = 29'b1_101011101000_111_1_101011101000;
      patterns[55112] = 29'b1_101011101001_000_1_101011101001;
      patterns[55113] = 29'b1_101011101001_001_1_101001101011;
      patterns[55114] = 29'b1_101011101001_010_1_010111010011;
      patterns[55115] = 29'b1_101011101001_011_0_101110100111;
      patterns[55116] = 29'b1_101011101001_100_1_110101110100;
      patterns[55117] = 29'b1_101011101001_101_0_111010111010;
      patterns[55118] = 29'b1_101011101001_110_1_101011101001;
      patterns[55119] = 29'b1_101011101001_111_1_101011101001;
      patterns[55120] = 29'b1_101011101010_000_1_101011101010;
      patterns[55121] = 29'b1_101011101010_001_1_101010101011;
      patterns[55122] = 29'b1_101011101010_010_1_010111010101;
      patterns[55123] = 29'b1_101011101010_011_0_101110101011;
      patterns[55124] = 29'b1_101011101010_100_0_110101110101;
      patterns[55125] = 29'b1_101011101010_101_1_011010111010;
      patterns[55126] = 29'b1_101011101010_110_1_101011101010;
      patterns[55127] = 29'b1_101011101010_111_1_101011101010;
      patterns[55128] = 29'b1_101011101011_000_1_101011101011;
      patterns[55129] = 29'b1_101011101011_001_1_101011101011;
      patterns[55130] = 29'b1_101011101011_010_1_010111010111;
      patterns[55131] = 29'b1_101011101011_011_0_101110101111;
      patterns[55132] = 29'b1_101011101011_100_1_110101110101;
      patterns[55133] = 29'b1_101011101011_101_1_111010111010;
      patterns[55134] = 29'b1_101011101011_110_1_101011101011;
      patterns[55135] = 29'b1_101011101011_111_1_101011101011;
      patterns[55136] = 29'b1_101011101100_000_1_101011101100;
      patterns[55137] = 29'b1_101011101100_001_1_101100101011;
      patterns[55138] = 29'b1_101011101100_010_1_010111011001;
      patterns[55139] = 29'b1_101011101100_011_0_101110110011;
      patterns[55140] = 29'b1_101011101100_100_0_110101110110;
      patterns[55141] = 29'b1_101011101100_101_0_011010111011;
      patterns[55142] = 29'b1_101011101100_110_1_101011101100;
      patterns[55143] = 29'b1_101011101100_111_1_101011101100;
      patterns[55144] = 29'b1_101011101101_000_1_101011101101;
      patterns[55145] = 29'b1_101011101101_001_1_101101101011;
      patterns[55146] = 29'b1_101011101101_010_1_010111011011;
      patterns[55147] = 29'b1_101011101101_011_0_101110110111;
      patterns[55148] = 29'b1_101011101101_100_1_110101110110;
      patterns[55149] = 29'b1_101011101101_101_0_111010111011;
      patterns[55150] = 29'b1_101011101101_110_1_101011101101;
      patterns[55151] = 29'b1_101011101101_111_1_101011101101;
      patterns[55152] = 29'b1_101011101110_000_1_101011101110;
      patterns[55153] = 29'b1_101011101110_001_1_101110101011;
      patterns[55154] = 29'b1_101011101110_010_1_010111011101;
      patterns[55155] = 29'b1_101011101110_011_0_101110111011;
      patterns[55156] = 29'b1_101011101110_100_0_110101110111;
      patterns[55157] = 29'b1_101011101110_101_1_011010111011;
      patterns[55158] = 29'b1_101011101110_110_1_101011101110;
      patterns[55159] = 29'b1_101011101110_111_1_101011101110;
      patterns[55160] = 29'b1_101011101111_000_1_101011101111;
      patterns[55161] = 29'b1_101011101111_001_1_101111101011;
      patterns[55162] = 29'b1_101011101111_010_1_010111011111;
      patterns[55163] = 29'b1_101011101111_011_0_101110111111;
      patterns[55164] = 29'b1_101011101111_100_1_110101110111;
      patterns[55165] = 29'b1_101011101111_101_1_111010111011;
      patterns[55166] = 29'b1_101011101111_110_1_101011101111;
      patterns[55167] = 29'b1_101011101111_111_1_101011101111;
      patterns[55168] = 29'b1_101011110000_000_1_101011110000;
      patterns[55169] = 29'b1_101011110000_001_1_110000101011;
      patterns[55170] = 29'b1_101011110000_010_1_010111100001;
      patterns[55171] = 29'b1_101011110000_011_0_101111000011;
      patterns[55172] = 29'b1_101011110000_100_0_110101111000;
      patterns[55173] = 29'b1_101011110000_101_0_011010111100;
      patterns[55174] = 29'b1_101011110000_110_1_101011110000;
      patterns[55175] = 29'b1_101011110000_111_1_101011110000;
      patterns[55176] = 29'b1_101011110001_000_1_101011110001;
      patterns[55177] = 29'b1_101011110001_001_1_110001101011;
      patterns[55178] = 29'b1_101011110001_010_1_010111100011;
      patterns[55179] = 29'b1_101011110001_011_0_101111000111;
      patterns[55180] = 29'b1_101011110001_100_1_110101111000;
      patterns[55181] = 29'b1_101011110001_101_0_111010111100;
      patterns[55182] = 29'b1_101011110001_110_1_101011110001;
      patterns[55183] = 29'b1_101011110001_111_1_101011110001;
      patterns[55184] = 29'b1_101011110010_000_1_101011110010;
      patterns[55185] = 29'b1_101011110010_001_1_110010101011;
      patterns[55186] = 29'b1_101011110010_010_1_010111100101;
      patterns[55187] = 29'b1_101011110010_011_0_101111001011;
      patterns[55188] = 29'b1_101011110010_100_0_110101111001;
      patterns[55189] = 29'b1_101011110010_101_1_011010111100;
      patterns[55190] = 29'b1_101011110010_110_1_101011110010;
      patterns[55191] = 29'b1_101011110010_111_1_101011110010;
      patterns[55192] = 29'b1_101011110011_000_1_101011110011;
      patterns[55193] = 29'b1_101011110011_001_1_110011101011;
      patterns[55194] = 29'b1_101011110011_010_1_010111100111;
      patterns[55195] = 29'b1_101011110011_011_0_101111001111;
      patterns[55196] = 29'b1_101011110011_100_1_110101111001;
      patterns[55197] = 29'b1_101011110011_101_1_111010111100;
      patterns[55198] = 29'b1_101011110011_110_1_101011110011;
      patterns[55199] = 29'b1_101011110011_111_1_101011110011;
      patterns[55200] = 29'b1_101011110100_000_1_101011110100;
      patterns[55201] = 29'b1_101011110100_001_1_110100101011;
      patterns[55202] = 29'b1_101011110100_010_1_010111101001;
      patterns[55203] = 29'b1_101011110100_011_0_101111010011;
      patterns[55204] = 29'b1_101011110100_100_0_110101111010;
      patterns[55205] = 29'b1_101011110100_101_0_011010111101;
      patterns[55206] = 29'b1_101011110100_110_1_101011110100;
      patterns[55207] = 29'b1_101011110100_111_1_101011110100;
      patterns[55208] = 29'b1_101011110101_000_1_101011110101;
      patterns[55209] = 29'b1_101011110101_001_1_110101101011;
      patterns[55210] = 29'b1_101011110101_010_1_010111101011;
      patterns[55211] = 29'b1_101011110101_011_0_101111010111;
      patterns[55212] = 29'b1_101011110101_100_1_110101111010;
      patterns[55213] = 29'b1_101011110101_101_0_111010111101;
      patterns[55214] = 29'b1_101011110101_110_1_101011110101;
      patterns[55215] = 29'b1_101011110101_111_1_101011110101;
      patterns[55216] = 29'b1_101011110110_000_1_101011110110;
      patterns[55217] = 29'b1_101011110110_001_1_110110101011;
      patterns[55218] = 29'b1_101011110110_010_1_010111101101;
      patterns[55219] = 29'b1_101011110110_011_0_101111011011;
      patterns[55220] = 29'b1_101011110110_100_0_110101111011;
      patterns[55221] = 29'b1_101011110110_101_1_011010111101;
      patterns[55222] = 29'b1_101011110110_110_1_101011110110;
      patterns[55223] = 29'b1_101011110110_111_1_101011110110;
      patterns[55224] = 29'b1_101011110111_000_1_101011110111;
      patterns[55225] = 29'b1_101011110111_001_1_110111101011;
      patterns[55226] = 29'b1_101011110111_010_1_010111101111;
      patterns[55227] = 29'b1_101011110111_011_0_101111011111;
      patterns[55228] = 29'b1_101011110111_100_1_110101111011;
      patterns[55229] = 29'b1_101011110111_101_1_111010111101;
      patterns[55230] = 29'b1_101011110111_110_1_101011110111;
      patterns[55231] = 29'b1_101011110111_111_1_101011110111;
      patterns[55232] = 29'b1_101011111000_000_1_101011111000;
      patterns[55233] = 29'b1_101011111000_001_1_111000101011;
      patterns[55234] = 29'b1_101011111000_010_1_010111110001;
      patterns[55235] = 29'b1_101011111000_011_0_101111100011;
      patterns[55236] = 29'b1_101011111000_100_0_110101111100;
      patterns[55237] = 29'b1_101011111000_101_0_011010111110;
      patterns[55238] = 29'b1_101011111000_110_1_101011111000;
      patterns[55239] = 29'b1_101011111000_111_1_101011111000;
      patterns[55240] = 29'b1_101011111001_000_1_101011111001;
      patterns[55241] = 29'b1_101011111001_001_1_111001101011;
      patterns[55242] = 29'b1_101011111001_010_1_010111110011;
      patterns[55243] = 29'b1_101011111001_011_0_101111100111;
      patterns[55244] = 29'b1_101011111001_100_1_110101111100;
      patterns[55245] = 29'b1_101011111001_101_0_111010111110;
      patterns[55246] = 29'b1_101011111001_110_1_101011111001;
      patterns[55247] = 29'b1_101011111001_111_1_101011111001;
      patterns[55248] = 29'b1_101011111010_000_1_101011111010;
      patterns[55249] = 29'b1_101011111010_001_1_111010101011;
      patterns[55250] = 29'b1_101011111010_010_1_010111110101;
      patterns[55251] = 29'b1_101011111010_011_0_101111101011;
      patterns[55252] = 29'b1_101011111010_100_0_110101111101;
      patterns[55253] = 29'b1_101011111010_101_1_011010111110;
      patterns[55254] = 29'b1_101011111010_110_1_101011111010;
      patterns[55255] = 29'b1_101011111010_111_1_101011111010;
      patterns[55256] = 29'b1_101011111011_000_1_101011111011;
      patterns[55257] = 29'b1_101011111011_001_1_111011101011;
      patterns[55258] = 29'b1_101011111011_010_1_010111110111;
      patterns[55259] = 29'b1_101011111011_011_0_101111101111;
      patterns[55260] = 29'b1_101011111011_100_1_110101111101;
      patterns[55261] = 29'b1_101011111011_101_1_111010111110;
      patterns[55262] = 29'b1_101011111011_110_1_101011111011;
      patterns[55263] = 29'b1_101011111011_111_1_101011111011;
      patterns[55264] = 29'b1_101011111100_000_1_101011111100;
      patterns[55265] = 29'b1_101011111100_001_1_111100101011;
      patterns[55266] = 29'b1_101011111100_010_1_010111111001;
      patterns[55267] = 29'b1_101011111100_011_0_101111110011;
      patterns[55268] = 29'b1_101011111100_100_0_110101111110;
      patterns[55269] = 29'b1_101011111100_101_0_011010111111;
      patterns[55270] = 29'b1_101011111100_110_1_101011111100;
      patterns[55271] = 29'b1_101011111100_111_1_101011111100;
      patterns[55272] = 29'b1_101011111101_000_1_101011111101;
      patterns[55273] = 29'b1_101011111101_001_1_111101101011;
      patterns[55274] = 29'b1_101011111101_010_1_010111111011;
      patterns[55275] = 29'b1_101011111101_011_0_101111110111;
      patterns[55276] = 29'b1_101011111101_100_1_110101111110;
      patterns[55277] = 29'b1_101011111101_101_0_111010111111;
      patterns[55278] = 29'b1_101011111101_110_1_101011111101;
      patterns[55279] = 29'b1_101011111101_111_1_101011111101;
      patterns[55280] = 29'b1_101011111110_000_1_101011111110;
      patterns[55281] = 29'b1_101011111110_001_1_111110101011;
      patterns[55282] = 29'b1_101011111110_010_1_010111111101;
      patterns[55283] = 29'b1_101011111110_011_0_101111111011;
      patterns[55284] = 29'b1_101011111110_100_0_110101111111;
      patterns[55285] = 29'b1_101011111110_101_1_011010111111;
      patterns[55286] = 29'b1_101011111110_110_1_101011111110;
      patterns[55287] = 29'b1_101011111110_111_1_101011111110;
      patterns[55288] = 29'b1_101011111111_000_1_101011111111;
      patterns[55289] = 29'b1_101011111111_001_1_111111101011;
      patterns[55290] = 29'b1_101011111111_010_1_010111111111;
      patterns[55291] = 29'b1_101011111111_011_0_101111111111;
      patterns[55292] = 29'b1_101011111111_100_1_110101111111;
      patterns[55293] = 29'b1_101011111111_101_1_111010111111;
      patterns[55294] = 29'b1_101011111111_110_1_101011111111;
      patterns[55295] = 29'b1_101011111111_111_1_101011111111;
      patterns[55296] = 29'b1_101100000000_000_1_101100000000;
      patterns[55297] = 29'b1_101100000000_001_1_000000101100;
      patterns[55298] = 29'b1_101100000000_010_1_011000000001;
      patterns[55299] = 29'b1_101100000000_011_0_110000000011;
      patterns[55300] = 29'b1_101100000000_100_0_110110000000;
      patterns[55301] = 29'b1_101100000000_101_0_011011000000;
      patterns[55302] = 29'b1_101100000000_110_1_101100000000;
      patterns[55303] = 29'b1_101100000000_111_1_101100000000;
      patterns[55304] = 29'b1_101100000001_000_1_101100000001;
      patterns[55305] = 29'b1_101100000001_001_1_000001101100;
      patterns[55306] = 29'b1_101100000001_010_1_011000000011;
      patterns[55307] = 29'b1_101100000001_011_0_110000000111;
      patterns[55308] = 29'b1_101100000001_100_1_110110000000;
      patterns[55309] = 29'b1_101100000001_101_0_111011000000;
      patterns[55310] = 29'b1_101100000001_110_1_101100000001;
      patterns[55311] = 29'b1_101100000001_111_1_101100000001;
      patterns[55312] = 29'b1_101100000010_000_1_101100000010;
      patterns[55313] = 29'b1_101100000010_001_1_000010101100;
      patterns[55314] = 29'b1_101100000010_010_1_011000000101;
      patterns[55315] = 29'b1_101100000010_011_0_110000001011;
      patterns[55316] = 29'b1_101100000010_100_0_110110000001;
      patterns[55317] = 29'b1_101100000010_101_1_011011000000;
      patterns[55318] = 29'b1_101100000010_110_1_101100000010;
      patterns[55319] = 29'b1_101100000010_111_1_101100000010;
      patterns[55320] = 29'b1_101100000011_000_1_101100000011;
      patterns[55321] = 29'b1_101100000011_001_1_000011101100;
      patterns[55322] = 29'b1_101100000011_010_1_011000000111;
      patterns[55323] = 29'b1_101100000011_011_0_110000001111;
      patterns[55324] = 29'b1_101100000011_100_1_110110000001;
      patterns[55325] = 29'b1_101100000011_101_1_111011000000;
      patterns[55326] = 29'b1_101100000011_110_1_101100000011;
      patterns[55327] = 29'b1_101100000011_111_1_101100000011;
      patterns[55328] = 29'b1_101100000100_000_1_101100000100;
      patterns[55329] = 29'b1_101100000100_001_1_000100101100;
      patterns[55330] = 29'b1_101100000100_010_1_011000001001;
      patterns[55331] = 29'b1_101100000100_011_0_110000010011;
      patterns[55332] = 29'b1_101100000100_100_0_110110000010;
      patterns[55333] = 29'b1_101100000100_101_0_011011000001;
      patterns[55334] = 29'b1_101100000100_110_1_101100000100;
      patterns[55335] = 29'b1_101100000100_111_1_101100000100;
      patterns[55336] = 29'b1_101100000101_000_1_101100000101;
      patterns[55337] = 29'b1_101100000101_001_1_000101101100;
      patterns[55338] = 29'b1_101100000101_010_1_011000001011;
      patterns[55339] = 29'b1_101100000101_011_0_110000010111;
      patterns[55340] = 29'b1_101100000101_100_1_110110000010;
      patterns[55341] = 29'b1_101100000101_101_0_111011000001;
      patterns[55342] = 29'b1_101100000101_110_1_101100000101;
      patterns[55343] = 29'b1_101100000101_111_1_101100000101;
      patterns[55344] = 29'b1_101100000110_000_1_101100000110;
      patterns[55345] = 29'b1_101100000110_001_1_000110101100;
      patterns[55346] = 29'b1_101100000110_010_1_011000001101;
      patterns[55347] = 29'b1_101100000110_011_0_110000011011;
      patterns[55348] = 29'b1_101100000110_100_0_110110000011;
      patterns[55349] = 29'b1_101100000110_101_1_011011000001;
      patterns[55350] = 29'b1_101100000110_110_1_101100000110;
      patterns[55351] = 29'b1_101100000110_111_1_101100000110;
      patterns[55352] = 29'b1_101100000111_000_1_101100000111;
      patterns[55353] = 29'b1_101100000111_001_1_000111101100;
      patterns[55354] = 29'b1_101100000111_010_1_011000001111;
      patterns[55355] = 29'b1_101100000111_011_0_110000011111;
      patterns[55356] = 29'b1_101100000111_100_1_110110000011;
      patterns[55357] = 29'b1_101100000111_101_1_111011000001;
      patterns[55358] = 29'b1_101100000111_110_1_101100000111;
      patterns[55359] = 29'b1_101100000111_111_1_101100000111;
      patterns[55360] = 29'b1_101100001000_000_1_101100001000;
      patterns[55361] = 29'b1_101100001000_001_1_001000101100;
      patterns[55362] = 29'b1_101100001000_010_1_011000010001;
      patterns[55363] = 29'b1_101100001000_011_0_110000100011;
      patterns[55364] = 29'b1_101100001000_100_0_110110000100;
      patterns[55365] = 29'b1_101100001000_101_0_011011000010;
      patterns[55366] = 29'b1_101100001000_110_1_101100001000;
      patterns[55367] = 29'b1_101100001000_111_1_101100001000;
      patterns[55368] = 29'b1_101100001001_000_1_101100001001;
      patterns[55369] = 29'b1_101100001001_001_1_001001101100;
      patterns[55370] = 29'b1_101100001001_010_1_011000010011;
      patterns[55371] = 29'b1_101100001001_011_0_110000100111;
      patterns[55372] = 29'b1_101100001001_100_1_110110000100;
      patterns[55373] = 29'b1_101100001001_101_0_111011000010;
      patterns[55374] = 29'b1_101100001001_110_1_101100001001;
      patterns[55375] = 29'b1_101100001001_111_1_101100001001;
      patterns[55376] = 29'b1_101100001010_000_1_101100001010;
      patterns[55377] = 29'b1_101100001010_001_1_001010101100;
      patterns[55378] = 29'b1_101100001010_010_1_011000010101;
      patterns[55379] = 29'b1_101100001010_011_0_110000101011;
      patterns[55380] = 29'b1_101100001010_100_0_110110000101;
      patterns[55381] = 29'b1_101100001010_101_1_011011000010;
      patterns[55382] = 29'b1_101100001010_110_1_101100001010;
      patterns[55383] = 29'b1_101100001010_111_1_101100001010;
      patterns[55384] = 29'b1_101100001011_000_1_101100001011;
      patterns[55385] = 29'b1_101100001011_001_1_001011101100;
      patterns[55386] = 29'b1_101100001011_010_1_011000010111;
      patterns[55387] = 29'b1_101100001011_011_0_110000101111;
      patterns[55388] = 29'b1_101100001011_100_1_110110000101;
      patterns[55389] = 29'b1_101100001011_101_1_111011000010;
      patterns[55390] = 29'b1_101100001011_110_1_101100001011;
      patterns[55391] = 29'b1_101100001011_111_1_101100001011;
      patterns[55392] = 29'b1_101100001100_000_1_101100001100;
      patterns[55393] = 29'b1_101100001100_001_1_001100101100;
      patterns[55394] = 29'b1_101100001100_010_1_011000011001;
      patterns[55395] = 29'b1_101100001100_011_0_110000110011;
      patterns[55396] = 29'b1_101100001100_100_0_110110000110;
      patterns[55397] = 29'b1_101100001100_101_0_011011000011;
      patterns[55398] = 29'b1_101100001100_110_1_101100001100;
      patterns[55399] = 29'b1_101100001100_111_1_101100001100;
      patterns[55400] = 29'b1_101100001101_000_1_101100001101;
      patterns[55401] = 29'b1_101100001101_001_1_001101101100;
      patterns[55402] = 29'b1_101100001101_010_1_011000011011;
      patterns[55403] = 29'b1_101100001101_011_0_110000110111;
      patterns[55404] = 29'b1_101100001101_100_1_110110000110;
      patterns[55405] = 29'b1_101100001101_101_0_111011000011;
      patterns[55406] = 29'b1_101100001101_110_1_101100001101;
      patterns[55407] = 29'b1_101100001101_111_1_101100001101;
      patterns[55408] = 29'b1_101100001110_000_1_101100001110;
      patterns[55409] = 29'b1_101100001110_001_1_001110101100;
      patterns[55410] = 29'b1_101100001110_010_1_011000011101;
      patterns[55411] = 29'b1_101100001110_011_0_110000111011;
      patterns[55412] = 29'b1_101100001110_100_0_110110000111;
      patterns[55413] = 29'b1_101100001110_101_1_011011000011;
      patterns[55414] = 29'b1_101100001110_110_1_101100001110;
      patterns[55415] = 29'b1_101100001110_111_1_101100001110;
      patterns[55416] = 29'b1_101100001111_000_1_101100001111;
      patterns[55417] = 29'b1_101100001111_001_1_001111101100;
      patterns[55418] = 29'b1_101100001111_010_1_011000011111;
      patterns[55419] = 29'b1_101100001111_011_0_110000111111;
      patterns[55420] = 29'b1_101100001111_100_1_110110000111;
      patterns[55421] = 29'b1_101100001111_101_1_111011000011;
      patterns[55422] = 29'b1_101100001111_110_1_101100001111;
      patterns[55423] = 29'b1_101100001111_111_1_101100001111;
      patterns[55424] = 29'b1_101100010000_000_1_101100010000;
      patterns[55425] = 29'b1_101100010000_001_1_010000101100;
      patterns[55426] = 29'b1_101100010000_010_1_011000100001;
      patterns[55427] = 29'b1_101100010000_011_0_110001000011;
      patterns[55428] = 29'b1_101100010000_100_0_110110001000;
      patterns[55429] = 29'b1_101100010000_101_0_011011000100;
      patterns[55430] = 29'b1_101100010000_110_1_101100010000;
      patterns[55431] = 29'b1_101100010000_111_1_101100010000;
      patterns[55432] = 29'b1_101100010001_000_1_101100010001;
      patterns[55433] = 29'b1_101100010001_001_1_010001101100;
      patterns[55434] = 29'b1_101100010001_010_1_011000100011;
      patterns[55435] = 29'b1_101100010001_011_0_110001000111;
      patterns[55436] = 29'b1_101100010001_100_1_110110001000;
      patterns[55437] = 29'b1_101100010001_101_0_111011000100;
      patterns[55438] = 29'b1_101100010001_110_1_101100010001;
      patterns[55439] = 29'b1_101100010001_111_1_101100010001;
      patterns[55440] = 29'b1_101100010010_000_1_101100010010;
      patterns[55441] = 29'b1_101100010010_001_1_010010101100;
      patterns[55442] = 29'b1_101100010010_010_1_011000100101;
      patterns[55443] = 29'b1_101100010010_011_0_110001001011;
      patterns[55444] = 29'b1_101100010010_100_0_110110001001;
      patterns[55445] = 29'b1_101100010010_101_1_011011000100;
      patterns[55446] = 29'b1_101100010010_110_1_101100010010;
      patterns[55447] = 29'b1_101100010010_111_1_101100010010;
      patterns[55448] = 29'b1_101100010011_000_1_101100010011;
      patterns[55449] = 29'b1_101100010011_001_1_010011101100;
      patterns[55450] = 29'b1_101100010011_010_1_011000100111;
      patterns[55451] = 29'b1_101100010011_011_0_110001001111;
      patterns[55452] = 29'b1_101100010011_100_1_110110001001;
      patterns[55453] = 29'b1_101100010011_101_1_111011000100;
      patterns[55454] = 29'b1_101100010011_110_1_101100010011;
      patterns[55455] = 29'b1_101100010011_111_1_101100010011;
      patterns[55456] = 29'b1_101100010100_000_1_101100010100;
      patterns[55457] = 29'b1_101100010100_001_1_010100101100;
      patterns[55458] = 29'b1_101100010100_010_1_011000101001;
      patterns[55459] = 29'b1_101100010100_011_0_110001010011;
      patterns[55460] = 29'b1_101100010100_100_0_110110001010;
      patterns[55461] = 29'b1_101100010100_101_0_011011000101;
      patterns[55462] = 29'b1_101100010100_110_1_101100010100;
      patterns[55463] = 29'b1_101100010100_111_1_101100010100;
      patterns[55464] = 29'b1_101100010101_000_1_101100010101;
      patterns[55465] = 29'b1_101100010101_001_1_010101101100;
      patterns[55466] = 29'b1_101100010101_010_1_011000101011;
      patterns[55467] = 29'b1_101100010101_011_0_110001010111;
      patterns[55468] = 29'b1_101100010101_100_1_110110001010;
      patterns[55469] = 29'b1_101100010101_101_0_111011000101;
      patterns[55470] = 29'b1_101100010101_110_1_101100010101;
      patterns[55471] = 29'b1_101100010101_111_1_101100010101;
      patterns[55472] = 29'b1_101100010110_000_1_101100010110;
      patterns[55473] = 29'b1_101100010110_001_1_010110101100;
      patterns[55474] = 29'b1_101100010110_010_1_011000101101;
      patterns[55475] = 29'b1_101100010110_011_0_110001011011;
      patterns[55476] = 29'b1_101100010110_100_0_110110001011;
      patterns[55477] = 29'b1_101100010110_101_1_011011000101;
      patterns[55478] = 29'b1_101100010110_110_1_101100010110;
      patterns[55479] = 29'b1_101100010110_111_1_101100010110;
      patterns[55480] = 29'b1_101100010111_000_1_101100010111;
      patterns[55481] = 29'b1_101100010111_001_1_010111101100;
      patterns[55482] = 29'b1_101100010111_010_1_011000101111;
      patterns[55483] = 29'b1_101100010111_011_0_110001011111;
      patterns[55484] = 29'b1_101100010111_100_1_110110001011;
      patterns[55485] = 29'b1_101100010111_101_1_111011000101;
      patterns[55486] = 29'b1_101100010111_110_1_101100010111;
      patterns[55487] = 29'b1_101100010111_111_1_101100010111;
      patterns[55488] = 29'b1_101100011000_000_1_101100011000;
      patterns[55489] = 29'b1_101100011000_001_1_011000101100;
      patterns[55490] = 29'b1_101100011000_010_1_011000110001;
      patterns[55491] = 29'b1_101100011000_011_0_110001100011;
      patterns[55492] = 29'b1_101100011000_100_0_110110001100;
      patterns[55493] = 29'b1_101100011000_101_0_011011000110;
      patterns[55494] = 29'b1_101100011000_110_1_101100011000;
      patterns[55495] = 29'b1_101100011000_111_1_101100011000;
      patterns[55496] = 29'b1_101100011001_000_1_101100011001;
      patterns[55497] = 29'b1_101100011001_001_1_011001101100;
      patterns[55498] = 29'b1_101100011001_010_1_011000110011;
      patterns[55499] = 29'b1_101100011001_011_0_110001100111;
      patterns[55500] = 29'b1_101100011001_100_1_110110001100;
      patterns[55501] = 29'b1_101100011001_101_0_111011000110;
      patterns[55502] = 29'b1_101100011001_110_1_101100011001;
      patterns[55503] = 29'b1_101100011001_111_1_101100011001;
      patterns[55504] = 29'b1_101100011010_000_1_101100011010;
      patterns[55505] = 29'b1_101100011010_001_1_011010101100;
      patterns[55506] = 29'b1_101100011010_010_1_011000110101;
      patterns[55507] = 29'b1_101100011010_011_0_110001101011;
      patterns[55508] = 29'b1_101100011010_100_0_110110001101;
      patterns[55509] = 29'b1_101100011010_101_1_011011000110;
      patterns[55510] = 29'b1_101100011010_110_1_101100011010;
      patterns[55511] = 29'b1_101100011010_111_1_101100011010;
      patterns[55512] = 29'b1_101100011011_000_1_101100011011;
      patterns[55513] = 29'b1_101100011011_001_1_011011101100;
      patterns[55514] = 29'b1_101100011011_010_1_011000110111;
      patterns[55515] = 29'b1_101100011011_011_0_110001101111;
      patterns[55516] = 29'b1_101100011011_100_1_110110001101;
      patterns[55517] = 29'b1_101100011011_101_1_111011000110;
      patterns[55518] = 29'b1_101100011011_110_1_101100011011;
      patterns[55519] = 29'b1_101100011011_111_1_101100011011;
      patterns[55520] = 29'b1_101100011100_000_1_101100011100;
      patterns[55521] = 29'b1_101100011100_001_1_011100101100;
      patterns[55522] = 29'b1_101100011100_010_1_011000111001;
      patterns[55523] = 29'b1_101100011100_011_0_110001110011;
      patterns[55524] = 29'b1_101100011100_100_0_110110001110;
      patterns[55525] = 29'b1_101100011100_101_0_011011000111;
      patterns[55526] = 29'b1_101100011100_110_1_101100011100;
      patterns[55527] = 29'b1_101100011100_111_1_101100011100;
      patterns[55528] = 29'b1_101100011101_000_1_101100011101;
      patterns[55529] = 29'b1_101100011101_001_1_011101101100;
      patterns[55530] = 29'b1_101100011101_010_1_011000111011;
      patterns[55531] = 29'b1_101100011101_011_0_110001110111;
      patterns[55532] = 29'b1_101100011101_100_1_110110001110;
      patterns[55533] = 29'b1_101100011101_101_0_111011000111;
      patterns[55534] = 29'b1_101100011101_110_1_101100011101;
      patterns[55535] = 29'b1_101100011101_111_1_101100011101;
      patterns[55536] = 29'b1_101100011110_000_1_101100011110;
      patterns[55537] = 29'b1_101100011110_001_1_011110101100;
      patterns[55538] = 29'b1_101100011110_010_1_011000111101;
      patterns[55539] = 29'b1_101100011110_011_0_110001111011;
      patterns[55540] = 29'b1_101100011110_100_0_110110001111;
      patterns[55541] = 29'b1_101100011110_101_1_011011000111;
      patterns[55542] = 29'b1_101100011110_110_1_101100011110;
      patterns[55543] = 29'b1_101100011110_111_1_101100011110;
      patterns[55544] = 29'b1_101100011111_000_1_101100011111;
      patterns[55545] = 29'b1_101100011111_001_1_011111101100;
      patterns[55546] = 29'b1_101100011111_010_1_011000111111;
      patterns[55547] = 29'b1_101100011111_011_0_110001111111;
      patterns[55548] = 29'b1_101100011111_100_1_110110001111;
      patterns[55549] = 29'b1_101100011111_101_1_111011000111;
      patterns[55550] = 29'b1_101100011111_110_1_101100011111;
      patterns[55551] = 29'b1_101100011111_111_1_101100011111;
      patterns[55552] = 29'b1_101100100000_000_1_101100100000;
      patterns[55553] = 29'b1_101100100000_001_1_100000101100;
      patterns[55554] = 29'b1_101100100000_010_1_011001000001;
      patterns[55555] = 29'b1_101100100000_011_0_110010000011;
      patterns[55556] = 29'b1_101100100000_100_0_110110010000;
      patterns[55557] = 29'b1_101100100000_101_0_011011001000;
      patterns[55558] = 29'b1_101100100000_110_1_101100100000;
      patterns[55559] = 29'b1_101100100000_111_1_101100100000;
      patterns[55560] = 29'b1_101100100001_000_1_101100100001;
      patterns[55561] = 29'b1_101100100001_001_1_100001101100;
      patterns[55562] = 29'b1_101100100001_010_1_011001000011;
      patterns[55563] = 29'b1_101100100001_011_0_110010000111;
      patterns[55564] = 29'b1_101100100001_100_1_110110010000;
      patterns[55565] = 29'b1_101100100001_101_0_111011001000;
      patterns[55566] = 29'b1_101100100001_110_1_101100100001;
      patterns[55567] = 29'b1_101100100001_111_1_101100100001;
      patterns[55568] = 29'b1_101100100010_000_1_101100100010;
      patterns[55569] = 29'b1_101100100010_001_1_100010101100;
      patterns[55570] = 29'b1_101100100010_010_1_011001000101;
      patterns[55571] = 29'b1_101100100010_011_0_110010001011;
      patterns[55572] = 29'b1_101100100010_100_0_110110010001;
      patterns[55573] = 29'b1_101100100010_101_1_011011001000;
      patterns[55574] = 29'b1_101100100010_110_1_101100100010;
      patterns[55575] = 29'b1_101100100010_111_1_101100100010;
      patterns[55576] = 29'b1_101100100011_000_1_101100100011;
      patterns[55577] = 29'b1_101100100011_001_1_100011101100;
      patterns[55578] = 29'b1_101100100011_010_1_011001000111;
      patterns[55579] = 29'b1_101100100011_011_0_110010001111;
      patterns[55580] = 29'b1_101100100011_100_1_110110010001;
      patterns[55581] = 29'b1_101100100011_101_1_111011001000;
      patterns[55582] = 29'b1_101100100011_110_1_101100100011;
      patterns[55583] = 29'b1_101100100011_111_1_101100100011;
      patterns[55584] = 29'b1_101100100100_000_1_101100100100;
      patterns[55585] = 29'b1_101100100100_001_1_100100101100;
      patterns[55586] = 29'b1_101100100100_010_1_011001001001;
      patterns[55587] = 29'b1_101100100100_011_0_110010010011;
      patterns[55588] = 29'b1_101100100100_100_0_110110010010;
      patterns[55589] = 29'b1_101100100100_101_0_011011001001;
      patterns[55590] = 29'b1_101100100100_110_1_101100100100;
      patterns[55591] = 29'b1_101100100100_111_1_101100100100;
      patterns[55592] = 29'b1_101100100101_000_1_101100100101;
      patterns[55593] = 29'b1_101100100101_001_1_100101101100;
      patterns[55594] = 29'b1_101100100101_010_1_011001001011;
      patterns[55595] = 29'b1_101100100101_011_0_110010010111;
      patterns[55596] = 29'b1_101100100101_100_1_110110010010;
      patterns[55597] = 29'b1_101100100101_101_0_111011001001;
      patterns[55598] = 29'b1_101100100101_110_1_101100100101;
      patterns[55599] = 29'b1_101100100101_111_1_101100100101;
      patterns[55600] = 29'b1_101100100110_000_1_101100100110;
      patterns[55601] = 29'b1_101100100110_001_1_100110101100;
      patterns[55602] = 29'b1_101100100110_010_1_011001001101;
      patterns[55603] = 29'b1_101100100110_011_0_110010011011;
      patterns[55604] = 29'b1_101100100110_100_0_110110010011;
      patterns[55605] = 29'b1_101100100110_101_1_011011001001;
      patterns[55606] = 29'b1_101100100110_110_1_101100100110;
      patterns[55607] = 29'b1_101100100110_111_1_101100100110;
      patterns[55608] = 29'b1_101100100111_000_1_101100100111;
      patterns[55609] = 29'b1_101100100111_001_1_100111101100;
      patterns[55610] = 29'b1_101100100111_010_1_011001001111;
      patterns[55611] = 29'b1_101100100111_011_0_110010011111;
      patterns[55612] = 29'b1_101100100111_100_1_110110010011;
      patterns[55613] = 29'b1_101100100111_101_1_111011001001;
      patterns[55614] = 29'b1_101100100111_110_1_101100100111;
      patterns[55615] = 29'b1_101100100111_111_1_101100100111;
      patterns[55616] = 29'b1_101100101000_000_1_101100101000;
      patterns[55617] = 29'b1_101100101000_001_1_101000101100;
      patterns[55618] = 29'b1_101100101000_010_1_011001010001;
      patterns[55619] = 29'b1_101100101000_011_0_110010100011;
      patterns[55620] = 29'b1_101100101000_100_0_110110010100;
      patterns[55621] = 29'b1_101100101000_101_0_011011001010;
      patterns[55622] = 29'b1_101100101000_110_1_101100101000;
      patterns[55623] = 29'b1_101100101000_111_1_101100101000;
      patterns[55624] = 29'b1_101100101001_000_1_101100101001;
      patterns[55625] = 29'b1_101100101001_001_1_101001101100;
      patterns[55626] = 29'b1_101100101001_010_1_011001010011;
      patterns[55627] = 29'b1_101100101001_011_0_110010100111;
      patterns[55628] = 29'b1_101100101001_100_1_110110010100;
      patterns[55629] = 29'b1_101100101001_101_0_111011001010;
      patterns[55630] = 29'b1_101100101001_110_1_101100101001;
      patterns[55631] = 29'b1_101100101001_111_1_101100101001;
      patterns[55632] = 29'b1_101100101010_000_1_101100101010;
      patterns[55633] = 29'b1_101100101010_001_1_101010101100;
      patterns[55634] = 29'b1_101100101010_010_1_011001010101;
      patterns[55635] = 29'b1_101100101010_011_0_110010101011;
      patterns[55636] = 29'b1_101100101010_100_0_110110010101;
      patterns[55637] = 29'b1_101100101010_101_1_011011001010;
      patterns[55638] = 29'b1_101100101010_110_1_101100101010;
      patterns[55639] = 29'b1_101100101010_111_1_101100101010;
      patterns[55640] = 29'b1_101100101011_000_1_101100101011;
      patterns[55641] = 29'b1_101100101011_001_1_101011101100;
      patterns[55642] = 29'b1_101100101011_010_1_011001010111;
      patterns[55643] = 29'b1_101100101011_011_0_110010101111;
      patterns[55644] = 29'b1_101100101011_100_1_110110010101;
      patterns[55645] = 29'b1_101100101011_101_1_111011001010;
      patterns[55646] = 29'b1_101100101011_110_1_101100101011;
      patterns[55647] = 29'b1_101100101011_111_1_101100101011;
      patterns[55648] = 29'b1_101100101100_000_1_101100101100;
      patterns[55649] = 29'b1_101100101100_001_1_101100101100;
      patterns[55650] = 29'b1_101100101100_010_1_011001011001;
      patterns[55651] = 29'b1_101100101100_011_0_110010110011;
      patterns[55652] = 29'b1_101100101100_100_0_110110010110;
      patterns[55653] = 29'b1_101100101100_101_0_011011001011;
      patterns[55654] = 29'b1_101100101100_110_1_101100101100;
      patterns[55655] = 29'b1_101100101100_111_1_101100101100;
      patterns[55656] = 29'b1_101100101101_000_1_101100101101;
      patterns[55657] = 29'b1_101100101101_001_1_101101101100;
      patterns[55658] = 29'b1_101100101101_010_1_011001011011;
      patterns[55659] = 29'b1_101100101101_011_0_110010110111;
      patterns[55660] = 29'b1_101100101101_100_1_110110010110;
      patterns[55661] = 29'b1_101100101101_101_0_111011001011;
      patterns[55662] = 29'b1_101100101101_110_1_101100101101;
      patterns[55663] = 29'b1_101100101101_111_1_101100101101;
      patterns[55664] = 29'b1_101100101110_000_1_101100101110;
      patterns[55665] = 29'b1_101100101110_001_1_101110101100;
      patterns[55666] = 29'b1_101100101110_010_1_011001011101;
      patterns[55667] = 29'b1_101100101110_011_0_110010111011;
      patterns[55668] = 29'b1_101100101110_100_0_110110010111;
      patterns[55669] = 29'b1_101100101110_101_1_011011001011;
      patterns[55670] = 29'b1_101100101110_110_1_101100101110;
      patterns[55671] = 29'b1_101100101110_111_1_101100101110;
      patterns[55672] = 29'b1_101100101111_000_1_101100101111;
      patterns[55673] = 29'b1_101100101111_001_1_101111101100;
      patterns[55674] = 29'b1_101100101111_010_1_011001011111;
      patterns[55675] = 29'b1_101100101111_011_0_110010111111;
      patterns[55676] = 29'b1_101100101111_100_1_110110010111;
      patterns[55677] = 29'b1_101100101111_101_1_111011001011;
      patterns[55678] = 29'b1_101100101111_110_1_101100101111;
      patterns[55679] = 29'b1_101100101111_111_1_101100101111;
      patterns[55680] = 29'b1_101100110000_000_1_101100110000;
      patterns[55681] = 29'b1_101100110000_001_1_110000101100;
      patterns[55682] = 29'b1_101100110000_010_1_011001100001;
      patterns[55683] = 29'b1_101100110000_011_0_110011000011;
      patterns[55684] = 29'b1_101100110000_100_0_110110011000;
      patterns[55685] = 29'b1_101100110000_101_0_011011001100;
      patterns[55686] = 29'b1_101100110000_110_1_101100110000;
      patterns[55687] = 29'b1_101100110000_111_1_101100110000;
      patterns[55688] = 29'b1_101100110001_000_1_101100110001;
      patterns[55689] = 29'b1_101100110001_001_1_110001101100;
      patterns[55690] = 29'b1_101100110001_010_1_011001100011;
      patterns[55691] = 29'b1_101100110001_011_0_110011000111;
      patterns[55692] = 29'b1_101100110001_100_1_110110011000;
      patterns[55693] = 29'b1_101100110001_101_0_111011001100;
      patterns[55694] = 29'b1_101100110001_110_1_101100110001;
      patterns[55695] = 29'b1_101100110001_111_1_101100110001;
      patterns[55696] = 29'b1_101100110010_000_1_101100110010;
      patterns[55697] = 29'b1_101100110010_001_1_110010101100;
      patterns[55698] = 29'b1_101100110010_010_1_011001100101;
      patterns[55699] = 29'b1_101100110010_011_0_110011001011;
      patterns[55700] = 29'b1_101100110010_100_0_110110011001;
      patterns[55701] = 29'b1_101100110010_101_1_011011001100;
      patterns[55702] = 29'b1_101100110010_110_1_101100110010;
      patterns[55703] = 29'b1_101100110010_111_1_101100110010;
      patterns[55704] = 29'b1_101100110011_000_1_101100110011;
      patterns[55705] = 29'b1_101100110011_001_1_110011101100;
      patterns[55706] = 29'b1_101100110011_010_1_011001100111;
      patterns[55707] = 29'b1_101100110011_011_0_110011001111;
      patterns[55708] = 29'b1_101100110011_100_1_110110011001;
      patterns[55709] = 29'b1_101100110011_101_1_111011001100;
      patterns[55710] = 29'b1_101100110011_110_1_101100110011;
      patterns[55711] = 29'b1_101100110011_111_1_101100110011;
      patterns[55712] = 29'b1_101100110100_000_1_101100110100;
      patterns[55713] = 29'b1_101100110100_001_1_110100101100;
      patterns[55714] = 29'b1_101100110100_010_1_011001101001;
      patterns[55715] = 29'b1_101100110100_011_0_110011010011;
      patterns[55716] = 29'b1_101100110100_100_0_110110011010;
      patterns[55717] = 29'b1_101100110100_101_0_011011001101;
      patterns[55718] = 29'b1_101100110100_110_1_101100110100;
      patterns[55719] = 29'b1_101100110100_111_1_101100110100;
      patterns[55720] = 29'b1_101100110101_000_1_101100110101;
      patterns[55721] = 29'b1_101100110101_001_1_110101101100;
      patterns[55722] = 29'b1_101100110101_010_1_011001101011;
      patterns[55723] = 29'b1_101100110101_011_0_110011010111;
      patterns[55724] = 29'b1_101100110101_100_1_110110011010;
      patterns[55725] = 29'b1_101100110101_101_0_111011001101;
      patterns[55726] = 29'b1_101100110101_110_1_101100110101;
      patterns[55727] = 29'b1_101100110101_111_1_101100110101;
      patterns[55728] = 29'b1_101100110110_000_1_101100110110;
      patterns[55729] = 29'b1_101100110110_001_1_110110101100;
      patterns[55730] = 29'b1_101100110110_010_1_011001101101;
      patterns[55731] = 29'b1_101100110110_011_0_110011011011;
      patterns[55732] = 29'b1_101100110110_100_0_110110011011;
      patterns[55733] = 29'b1_101100110110_101_1_011011001101;
      patterns[55734] = 29'b1_101100110110_110_1_101100110110;
      patterns[55735] = 29'b1_101100110110_111_1_101100110110;
      patterns[55736] = 29'b1_101100110111_000_1_101100110111;
      patterns[55737] = 29'b1_101100110111_001_1_110111101100;
      patterns[55738] = 29'b1_101100110111_010_1_011001101111;
      patterns[55739] = 29'b1_101100110111_011_0_110011011111;
      patterns[55740] = 29'b1_101100110111_100_1_110110011011;
      patterns[55741] = 29'b1_101100110111_101_1_111011001101;
      patterns[55742] = 29'b1_101100110111_110_1_101100110111;
      patterns[55743] = 29'b1_101100110111_111_1_101100110111;
      patterns[55744] = 29'b1_101100111000_000_1_101100111000;
      patterns[55745] = 29'b1_101100111000_001_1_111000101100;
      patterns[55746] = 29'b1_101100111000_010_1_011001110001;
      patterns[55747] = 29'b1_101100111000_011_0_110011100011;
      patterns[55748] = 29'b1_101100111000_100_0_110110011100;
      patterns[55749] = 29'b1_101100111000_101_0_011011001110;
      patterns[55750] = 29'b1_101100111000_110_1_101100111000;
      patterns[55751] = 29'b1_101100111000_111_1_101100111000;
      patterns[55752] = 29'b1_101100111001_000_1_101100111001;
      patterns[55753] = 29'b1_101100111001_001_1_111001101100;
      patterns[55754] = 29'b1_101100111001_010_1_011001110011;
      patterns[55755] = 29'b1_101100111001_011_0_110011100111;
      patterns[55756] = 29'b1_101100111001_100_1_110110011100;
      patterns[55757] = 29'b1_101100111001_101_0_111011001110;
      patterns[55758] = 29'b1_101100111001_110_1_101100111001;
      patterns[55759] = 29'b1_101100111001_111_1_101100111001;
      patterns[55760] = 29'b1_101100111010_000_1_101100111010;
      patterns[55761] = 29'b1_101100111010_001_1_111010101100;
      patterns[55762] = 29'b1_101100111010_010_1_011001110101;
      patterns[55763] = 29'b1_101100111010_011_0_110011101011;
      patterns[55764] = 29'b1_101100111010_100_0_110110011101;
      patterns[55765] = 29'b1_101100111010_101_1_011011001110;
      patterns[55766] = 29'b1_101100111010_110_1_101100111010;
      patterns[55767] = 29'b1_101100111010_111_1_101100111010;
      patterns[55768] = 29'b1_101100111011_000_1_101100111011;
      patterns[55769] = 29'b1_101100111011_001_1_111011101100;
      patterns[55770] = 29'b1_101100111011_010_1_011001110111;
      patterns[55771] = 29'b1_101100111011_011_0_110011101111;
      patterns[55772] = 29'b1_101100111011_100_1_110110011101;
      patterns[55773] = 29'b1_101100111011_101_1_111011001110;
      patterns[55774] = 29'b1_101100111011_110_1_101100111011;
      patterns[55775] = 29'b1_101100111011_111_1_101100111011;
      patterns[55776] = 29'b1_101100111100_000_1_101100111100;
      patterns[55777] = 29'b1_101100111100_001_1_111100101100;
      patterns[55778] = 29'b1_101100111100_010_1_011001111001;
      patterns[55779] = 29'b1_101100111100_011_0_110011110011;
      patterns[55780] = 29'b1_101100111100_100_0_110110011110;
      patterns[55781] = 29'b1_101100111100_101_0_011011001111;
      patterns[55782] = 29'b1_101100111100_110_1_101100111100;
      patterns[55783] = 29'b1_101100111100_111_1_101100111100;
      patterns[55784] = 29'b1_101100111101_000_1_101100111101;
      patterns[55785] = 29'b1_101100111101_001_1_111101101100;
      patterns[55786] = 29'b1_101100111101_010_1_011001111011;
      patterns[55787] = 29'b1_101100111101_011_0_110011110111;
      patterns[55788] = 29'b1_101100111101_100_1_110110011110;
      patterns[55789] = 29'b1_101100111101_101_0_111011001111;
      patterns[55790] = 29'b1_101100111101_110_1_101100111101;
      patterns[55791] = 29'b1_101100111101_111_1_101100111101;
      patterns[55792] = 29'b1_101100111110_000_1_101100111110;
      patterns[55793] = 29'b1_101100111110_001_1_111110101100;
      patterns[55794] = 29'b1_101100111110_010_1_011001111101;
      patterns[55795] = 29'b1_101100111110_011_0_110011111011;
      patterns[55796] = 29'b1_101100111110_100_0_110110011111;
      patterns[55797] = 29'b1_101100111110_101_1_011011001111;
      patterns[55798] = 29'b1_101100111110_110_1_101100111110;
      patterns[55799] = 29'b1_101100111110_111_1_101100111110;
      patterns[55800] = 29'b1_101100111111_000_1_101100111111;
      patterns[55801] = 29'b1_101100111111_001_1_111111101100;
      patterns[55802] = 29'b1_101100111111_010_1_011001111111;
      patterns[55803] = 29'b1_101100111111_011_0_110011111111;
      patterns[55804] = 29'b1_101100111111_100_1_110110011111;
      patterns[55805] = 29'b1_101100111111_101_1_111011001111;
      patterns[55806] = 29'b1_101100111111_110_1_101100111111;
      patterns[55807] = 29'b1_101100111111_111_1_101100111111;
      patterns[55808] = 29'b1_101101000000_000_1_101101000000;
      patterns[55809] = 29'b1_101101000000_001_1_000000101101;
      patterns[55810] = 29'b1_101101000000_010_1_011010000001;
      patterns[55811] = 29'b1_101101000000_011_0_110100000011;
      patterns[55812] = 29'b1_101101000000_100_0_110110100000;
      patterns[55813] = 29'b1_101101000000_101_0_011011010000;
      patterns[55814] = 29'b1_101101000000_110_1_101101000000;
      patterns[55815] = 29'b1_101101000000_111_1_101101000000;
      patterns[55816] = 29'b1_101101000001_000_1_101101000001;
      patterns[55817] = 29'b1_101101000001_001_1_000001101101;
      patterns[55818] = 29'b1_101101000001_010_1_011010000011;
      patterns[55819] = 29'b1_101101000001_011_0_110100000111;
      patterns[55820] = 29'b1_101101000001_100_1_110110100000;
      patterns[55821] = 29'b1_101101000001_101_0_111011010000;
      patterns[55822] = 29'b1_101101000001_110_1_101101000001;
      patterns[55823] = 29'b1_101101000001_111_1_101101000001;
      patterns[55824] = 29'b1_101101000010_000_1_101101000010;
      patterns[55825] = 29'b1_101101000010_001_1_000010101101;
      patterns[55826] = 29'b1_101101000010_010_1_011010000101;
      patterns[55827] = 29'b1_101101000010_011_0_110100001011;
      patterns[55828] = 29'b1_101101000010_100_0_110110100001;
      patterns[55829] = 29'b1_101101000010_101_1_011011010000;
      patterns[55830] = 29'b1_101101000010_110_1_101101000010;
      patterns[55831] = 29'b1_101101000010_111_1_101101000010;
      patterns[55832] = 29'b1_101101000011_000_1_101101000011;
      patterns[55833] = 29'b1_101101000011_001_1_000011101101;
      patterns[55834] = 29'b1_101101000011_010_1_011010000111;
      patterns[55835] = 29'b1_101101000011_011_0_110100001111;
      patterns[55836] = 29'b1_101101000011_100_1_110110100001;
      patterns[55837] = 29'b1_101101000011_101_1_111011010000;
      patterns[55838] = 29'b1_101101000011_110_1_101101000011;
      patterns[55839] = 29'b1_101101000011_111_1_101101000011;
      patterns[55840] = 29'b1_101101000100_000_1_101101000100;
      patterns[55841] = 29'b1_101101000100_001_1_000100101101;
      patterns[55842] = 29'b1_101101000100_010_1_011010001001;
      patterns[55843] = 29'b1_101101000100_011_0_110100010011;
      patterns[55844] = 29'b1_101101000100_100_0_110110100010;
      patterns[55845] = 29'b1_101101000100_101_0_011011010001;
      patterns[55846] = 29'b1_101101000100_110_1_101101000100;
      patterns[55847] = 29'b1_101101000100_111_1_101101000100;
      patterns[55848] = 29'b1_101101000101_000_1_101101000101;
      patterns[55849] = 29'b1_101101000101_001_1_000101101101;
      patterns[55850] = 29'b1_101101000101_010_1_011010001011;
      patterns[55851] = 29'b1_101101000101_011_0_110100010111;
      patterns[55852] = 29'b1_101101000101_100_1_110110100010;
      patterns[55853] = 29'b1_101101000101_101_0_111011010001;
      patterns[55854] = 29'b1_101101000101_110_1_101101000101;
      patterns[55855] = 29'b1_101101000101_111_1_101101000101;
      patterns[55856] = 29'b1_101101000110_000_1_101101000110;
      patterns[55857] = 29'b1_101101000110_001_1_000110101101;
      patterns[55858] = 29'b1_101101000110_010_1_011010001101;
      patterns[55859] = 29'b1_101101000110_011_0_110100011011;
      patterns[55860] = 29'b1_101101000110_100_0_110110100011;
      patterns[55861] = 29'b1_101101000110_101_1_011011010001;
      patterns[55862] = 29'b1_101101000110_110_1_101101000110;
      patterns[55863] = 29'b1_101101000110_111_1_101101000110;
      patterns[55864] = 29'b1_101101000111_000_1_101101000111;
      patterns[55865] = 29'b1_101101000111_001_1_000111101101;
      patterns[55866] = 29'b1_101101000111_010_1_011010001111;
      patterns[55867] = 29'b1_101101000111_011_0_110100011111;
      patterns[55868] = 29'b1_101101000111_100_1_110110100011;
      patterns[55869] = 29'b1_101101000111_101_1_111011010001;
      patterns[55870] = 29'b1_101101000111_110_1_101101000111;
      patterns[55871] = 29'b1_101101000111_111_1_101101000111;
      patterns[55872] = 29'b1_101101001000_000_1_101101001000;
      patterns[55873] = 29'b1_101101001000_001_1_001000101101;
      patterns[55874] = 29'b1_101101001000_010_1_011010010001;
      patterns[55875] = 29'b1_101101001000_011_0_110100100011;
      patterns[55876] = 29'b1_101101001000_100_0_110110100100;
      patterns[55877] = 29'b1_101101001000_101_0_011011010010;
      patterns[55878] = 29'b1_101101001000_110_1_101101001000;
      patterns[55879] = 29'b1_101101001000_111_1_101101001000;
      patterns[55880] = 29'b1_101101001001_000_1_101101001001;
      patterns[55881] = 29'b1_101101001001_001_1_001001101101;
      patterns[55882] = 29'b1_101101001001_010_1_011010010011;
      patterns[55883] = 29'b1_101101001001_011_0_110100100111;
      patterns[55884] = 29'b1_101101001001_100_1_110110100100;
      patterns[55885] = 29'b1_101101001001_101_0_111011010010;
      patterns[55886] = 29'b1_101101001001_110_1_101101001001;
      patterns[55887] = 29'b1_101101001001_111_1_101101001001;
      patterns[55888] = 29'b1_101101001010_000_1_101101001010;
      patterns[55889] = 29'b1_101101001010_001_1_001010101101;
      patterns[55890] = 29'b1_101101001010_010_1_011010010101;
      patterns[55891] = 29'b1_101101001010_011_0_110100101011;
      patterns[55892] = 29'b1_101101001010_100_0_110110100101;
      patterns[55893] = 29'b1_101101001010_101_1_011011010010;
      patterns[55894] = 29'b1_101101001010_110_1_101101001010;
      patterns[55895] = 29'b1_101101001010_111_1_101101001010;
      patterns[55896] = 29'b1_101101001011_000_1_101101001011;
      patterns[55897] = 29'b1_101101001011_001_1_001011101101;
      patterns[55898] = 29'b1_101101001011_010_1_011010010111;
      patterns[55899] = 29'b1_101101001011_011_0_110100101111;
      patterns[55900] = 29'b1_101101001011_100_1_110110100101;
      patterns[55901] = 29'b1_101101001011_101_1_111011010010;
      patterns[55902] = 29'b1_101101001011_110_1_101101001011;
      patterns[55903] = 29'b1_101101001011_111_1_101101001011;
      patterns[55904] = 29'b1_101101001100_000_1_101101001100;
      patterns[55905] = 29'b1_101101001100_001_1_001100101101;
      patterns[55906] = 29'b1_101101001100_010_1_011010011001;
      patterns[55907] = 29'b1_101101001100_011_0_110100110011;
      patterns[55908] = 29'b1_101101001100_100_0_110110100110;
      patterns[55909] = 29'b1_101101001100_101_0_011011010011;
      patterns[55910] = 29'b1_101101001100_110_1_101101001100;
      patterns[55911] = 29'b1_101101001100_111_1_101101001100;
      patterns[55912] = 29'b1_101101001101_000_1_101101001101;
      patterns[55913] = 29'b1_101101001101_001_1_001101101101;
      patterns[55914] = 29'b1_101101001101_010_1_011010011011;
      patterns[55915] = 29'b1_101101001101_011_0_110100110111;
      patterns[55916] = 29'b1_101101001101_100_1_110110100110;
      patterns[55917] = 29'b1_101101001101_101_0_111011010011;
      patterns[55918] = 29'b1_101101001101_110_1_101101001101;
      patterns[55919] = 29'b1_101101001101_111_1_101101001101;
      patterns[55920] = 29'b1_101101001110_000_1_101101001110;
      patterns[55921] = 29'b1_101101001110_001_1_001110101101;
      patterns[55922] = 29'b1_101101001110_010_1_011010011101;
      patterns[55923] = 29'b1_101101001110_011_0_110100111011;
      patterns[55924] = 29'b1_101101001110_100_0_110110100111;
      patterns[55925] = 29'b1_101101001110_101_1_011011010011;
      patterns[55926] = 29'b1_101101001110_110_1_101101001110;
      patterns[55927] = 29'b1_101101001110_111_1_101101001110;
      patterns[55928] = 29'b1_101101001111_000_1_101101001111;
      patterns[55929] = 29'b1_101101001111_001_1_001111101101;
      patterns[55930] = 29'b1_101101001111_010_1_011010011111;
      patterns[55931] = 29'b1_101101001111_011_0_110100111111;
      patterns[55932] = 29'b1_101101001111_100_1_110110100111;
      patterns[55933] = 29'b1_101101001111_101_1_111011010011;
      patterns[55934] = 29'b1_101101001111_110_1_101101001111;
      patterns[55935] = 29'b1_101101001111_111_1_101101001111;
      patterns[55936] = 29'b1_101101010000_000_1_101101010000;
      patterns[55937] = 29'b1_101101010000_001_1_010000101101;
      patterns[55938] = 29'b1_101101010000_010_1_011010100001;
      patterns[55939] = 29'b1_101101010000_011_0_110101000011;
      patterns[55940] = 29'b1_101101010000_100_0_110110101000;
      patterns[55941] = 29'b1_101101010000_101_0_011011010100;
      patterns[55942] = 29'b1_101101010000_110_1_101101010000;
      patterns[55943] = 29'b1_101101010000_111_1_101101010000;
      patterns[55944] = 29'b1_101101010001_000_1_101101010001;
      patterns[55945] = 29'b1_101101010001_001_1_010001101101;
      patterns[55946] = 29'b1_101101010001_010_1_011010100011;
      patterns[55947] = 29'b1_101101010001_011_0_110101000111;
      patterns[55948] = 29'b1_101101010001_100_1_110110101000;
      patterns[55949] = 29'b1_101101010001_101_0_111011010100;
      patterns[55950] = 29'b1_101101010001_110_1_101101010001;
      patterns[55951] = 29'b1_101101010001_111_1_101101010001;
      patterns[55952] = 29'b1_101101010010_000_1_101101010010;
      patterns[55953] = 29'b1_101101010010_001_1_010010101101;
      patterns[55954] = 29'b1_101101010010_010_1_011010100101;
      patterns[55955] = 29'b1_101101010010_011_0_110101001011;
      patterns[55956] = 29'b1_101101010010_100_0_110110101001;
      patterns[55957] = 29'b1_101101010010_101_1_011011010100;
      patterns[55958] = 29'b1_101101010010_110_1_101101010010;
      patterns[55959] = 29'b1_101101010010_111_1_101101010010;
      patterns[55960] = 29'b1_101101010011_000_1_101101010011;
      patterns[55961] = 29'b1_101101010011_001_1_010011101101;
      patterns[55962] = 29'b1_101101010011_010_1_011010100111;
      patterns[55963] = 29'b1_101101010011_011_0_110101001111;
      patterns[55964] = 29'b1_101101010011_100_1_110110101001;
      patterns[55965] = 29'b1_101101010011_101_1_111011010100;
      patterns[55966] = 29'b1_101101010011_110_1_101101010011;
      patterns[55967] = 29'b1_101101010011_111_1_101101010011;
      patterns[55968] = 29'b1_101101010100_000_1_101101010100;
      patterns[55969] = 29'b1_101101010100_001_1_010100101101;
      patterns[55970] = 29'b1_101101010100_010_1_011010101001;
      patterns[55971] = 29'b1_101101010100_011_0_110101010011;
      patterns[55972] = 29'b1_101101010100_100_0_110110101010;
      patterns[55973] = 29'b1_101101010100_101_0_011011010101;
      patterns[55974] = 29'b1_101101010100_110_1_101101010100;
      patterns[55975] = 29'b1_101101010100_111_1_101101010100;
      patterns[55976] = 29'b1_101101010101_000_1_101101010101;
      patterns[55977] = 29'b1_101101010101_001_1_010101101101;
      patterns[55978] = 29'b1_101101010101_010_1_011010101011;
      patterns[55979] = 29'b1_101101010101_011_0_110101010111;
      patterns[55980] = 29'b1_101101010101_100_1_110110101010;
      patterns[55981] = 29'b1_101101010101_101_0_111011010101;
      patterns[55982] = 29'b1_101101010101_110_1_101101010101;
      patterns[55983] = 29'b1_101101010101_111_1_101101010101;
      patterns[55984] = 29'b1_101101010110_000_1_101101010110;
      patterns[55985] = 29'b1_101101010110_001_1_010110101101;
      patterns[55986] = 29'b1_101101010110_010_1_011010101101;
      patterns[55987] = 29'b1_101101010110_011_0_110101011011;
      patterns[55988] = 29'b1_101101010110_100_0_110110101011;
      patterns[55989] = 29'b1_101101010110_101_1_011011010101;
      patterns[55990] = 29'b1_101101010110_110_1_101101010110;
      patterns[55991] = 29'b1_101101010110_111_1_101101010110;
      patterns[55992] = 29'b1_101101010111_000_1_101101010111;
      patterns[55993] = 29'b1_101101010111_001_1_010111101101;
      patterns[55994] = 29'b1_101101010111_010_1_011010101111;
      patterns[55995] = 29'b1_101101010111_011_0_110101011111;
      patterns[55996] = 29'b1_101101010111_100_1_110110101011;
      patterns[55997] = 29'b1_101101010111_101_1_111011010101;
      patterns[55998] = 29'b1_101101010111_110_1_101101010111;
      patterns[55999] = 29'b1_101101010111_111_1_101101010111;
      patterns[56000] = 29'b1_101101011000_000_1_101101011000;
      patterns[56001] = 29'b1_101101011000_001_1_011000101101;
      patterns[56002] = 29'b1_101101011000_010_1_011010110001;
      patterns[56003] = 29'b1_101101011000_011_0_110101100011;
      patterns[56004] = 29'b1_101101011000_100_0_110110101100;
      patterns[56005] = 29'b1_101101011000_101_0_011011010110;
      patterns[56006] = 29'b1_101101011000_110_1_101101011000;
      patterns[56007] = 29'b1_101101011000_111_1_101101011000;
      patterns[56008] = 29'b1_101101011001_000_1_101101011001;
      patterns[56009] = 29'b1_101101011001_001_1_011001101101;
      patterns[56010] = 29'b1_101101011001_010_1_011010110011;
      patterns[56011] = 29'b1_101101011001_011_0_110101100111;
      patterns[56012] = 29'b1_101101011001_100_1_110110101100;
      patterns[56013] = 29'b1_101101011001_101_0_111011010110;
      patterns[56014] = 29'b1_101101011001_110_1_101101011001;
      patterns[56015] = 29'b1_101101011001_111_1_101101011001;
      patterns[56016] = 29'b1_101101011010_000_1_101101011010;
      patterns[56017] = 29'b1_101101011010_001_1_011010101101;
      patterns[56018] = 29'b1_101101011010_010_1_011010110101;
      patterns[56019] = 29'b1_101101011010_011_0_110101101011;
      patterns[56020] = 29'b1_101101011010_100_0_110110101101;
      patterns[56021] = 29'b1_101101011010_101_1_011011010110;
      patterns[56022] = 29'b1_101101011010_110_1_101101011010;
      patterns[56023] = 29'b1_101101011010_111_1_101101011010;
      patterns[56024] = 29'b1_101101011011_000_1_101101011011;
      patterns[56025] = 29'b1_101101011011_001_1_011011101101;
      patterns[56026] = 29'b1_101101011011_010_1_011010110111;
      patterns[56027] = 29'b1_101101011011_011_0_110101101111;
      patterns[56028] = 29'b1_101101011011_100_1_110110101101;
      patterns[56029] = 29'b1_101101011011_101_1_111011010110;
      patterns[56030] = 29'b1_101101011011_110_1_101101011011;
      patterns[56031] = 29'b1_101101011011_111_1_101101011011;
      patterns[56032] = 29'b1_101101011100_000_1_101101011100;
      patterns[56033] = 29'b1_101101011100_001_1_011100101101;
      patterns[56034] = 29'b1_101101011100_010_1_011010111001;
      patterns[56035] = 29'b1_101101011100_011_0_110101110011;
      patterns[56036] = 29'b1_101101011100_100_0_110110101110;
      patterns[56037] = 29'b1_101101011100_101_0_011011010111;
      patterns[56038] = 29'b1_101101011100_110_1_101101011100;
      patterns[56039] = 29'b1_101101011100_111_1_101101011100;
      patterns[56040] = 29'b1_101101011101_000_1_101101011101;
      patterns[56041] = 29'b1_101101011101_001_1_011101101101;
      patterns[56042] = 29'b1_101101011101_010_1_011010111011;
      patterns[56043] = 29'b1_101101011101_011_0_110101110111;
      patterns[56044] = 29'b1_101101011101_100_1_110110101110;
      patterns[56045] = 29'b1_101101011101_101_0_111011010111;
      patterns[56046] = 29'b1_101101011101_110_1_101101011101;
      patterns[56047] = 29'b1_101101011101_111_1_101101011101;
      patterns[56048] = 29'b1_101101011110_000_1_101101011110;
      patterns[56049] = 29'b1_101101011110_001_1_011110101101;
      patterns[56050] = 29'b1_101101011110_010_1_011010111101;
      patterns[56051] = 29'b1_101101011110_011_0_110101111011;
      patterns[56052] = 29'b1_101101011110_100_0_110110101111;
      patterns[56053] = 29'b1_101101011110_101_1_011011010111;
      patterns[56054] = 29'b1_101101011110_110_1_101101011110;
      patterns[56055] = 29'b1_101101011110_111_1_101101011110;
      patterns[56056] = 29'b1_101101011111_000_1_101101011111;
      patterns[56057] = 29'b1_101101011111_001_1_011111101101;
      patterns[56058] = 29'b1_101101011111_010_1_011010111111;
      patterns[56059] = 29'b1_101101011111_011_0_110101111111;
      patterns[56060] = 29'b1_101101011111_100_1_110110101111;
      patterns[56061] = 29'b1_101101011111_101_1_111011010111;
      patterns[56062] = 29'b1_101101011111_110_1_101101011111;
      patterns[56063] = 29'b1_101101011111_111_1_101101011111;
      patterns[56064] = 29'b1_101101100000_000_1_101101100000;
      patterns[56065] = 29'b1_101101100000_001_1_100000101101;
      patterns[56066] = 29'b1_101101100000_010_1_011011000001;
      patterns[56067] = 29'b1_101101100000_011_0_110110000011;
      patterns[56068] = 29'b1_101101100000_100_0_110110110000;
      patterns[56069] = 29'b1_101101100000_101_0_011011011000;
      patterns[56070] = 29'b1_101101100000_110_1_101101100000;
      patterns[56071] = 29'b1_101101100000_111_1_101101100000;
      patterns[56072] = 29'b1_101101100001_000_1_101101100001;
      patterns[56073] = 29'b1_101101100001_001_1_100001101101;
      patterns[56074] = 29'b1_101101100001_010_1_011011000011;
      patterns[56075] = 29'b1_101101100001_011_0_110110000111;
      patterns[56076] = 29'b1_101101100001_100_1_110110110000;
      patterns[56077] = 29'b1_101101100001_101_0_111011011000;
      patterns[56078] = 29'b1_101101100001_110_1_101101100001;
      patterns[56079] = 29'b1_101101100001_111_1_101101100001;
      patterns[56080] = 29'b1_101101100010_000_1_101101100010;
      patterns[56081] = 29'b1_101101100010_001_1_100010101101;
      patterns[56082] = 29'b1_101101100010_010_1_011011000101;
      patterns[56083] = 29'b1_101101100010_011_0_110110001011;
      patterns[56084] = 29'b1_101101100010_100_0_110110110001;
      patterns[56085] = 29'b1_101101100010_101_1_011011011000;
      patterns[56086] = 29'b1_101101100010_110_1_101101100010;
      patterns[56087] = 29'b1_101101100010_111_1_101101100010;
      patterns[56088] = 29'b1_101101100011_000_1_101101100011;
      patterns[56089] = 29'b1_101101100011_001_1_100011101101;
      patterns[56090] = 29'b1_101101100011_010_1_011011000111;
      patterns[56091] = 29'b1_101101100011_011_0_110110001111;
      patterns[56092] = 29'b1_101101100011_100_1_110110110001;
      patterns[56093] = 29'b1_101101100011_101_1_111011011000;
      patterns[56094] = 29'b1_101101100011_110_1_101101100011;
      patterns[56095] = 29'b1_101101100011_111_1_101101100011;
      patterns[56096] = 29'b1_101101100100_000_1_101101100100;
      patterns[56097] = 29'b1_101101100100_001_1_100100101101;
      patterns[56098] = 29'b1_101101100100_010_1_011011001001;
      patterns[56099] = 29'b1_101101100100_011_0_110110010011;
      patterns[56100] = 29'b1_101101100100_100_0_110110110010;
      patterns[56101] = 29'b1_101101100100_101_0_011011011001;
      patterns[56102] = 29'b1_101101100100_110_1_101101100100;
      patterns[56103] = 29'b1_101101100100_111_1_101101100100;
      patterns[56104] = 29'b1_101101100101_000_1_101101100101;
      patterns[56105] = 29'b1_101101100101_001_1_100101101101;
      patterns[56106] = 29'b1_101101100101_010_1_011011001011;
      patterns[56107] = 29'b1_101101100101_011_0_110110010111;
      patterns[56108] = 29'b1_101101100101_100_1_110110110010;
      patterns[56109] = 29'b1_101101100101_101_0_111011011001;
      patterns[56110] = 29'b1_101101100101_110_1_101101100101;
      patterns[56111] = 29'b1_101101100101_111_1_101101100101;
      patterns[56112] = 29'b1_101101100110_000_1_101101100110;
      patterns[56113] = 29'b1_101101100110_001_1_100110101101;
      patterns[56114] = 29'b1_101101100110_010_1_011011001101;
      patterns[56115] = 29'b1_101101100110_011_0_110110011011;
      patterns[56116] = 29'b1_101101100110_100_0_110110110011;
      patterns[56117] = 29'b1_101101100110_101_1_011011011001;
      patterns[56118] = 29'b1_101101100110_110_1_101101100110;
      patterns[56119] = 29'b1_101101100110_111_1_101101100110;
      patterns[56120] = 29'b1_101101100111_000_1_101101100111;
      patterns[56121] = 29'b1_101101100111_001_1_100111101101;
      patterns[56122] = 29'b1_101101100111_010_1_011011001111;
      patterns[56123] = 29'b1_101101100111_011_0_110110011111;
      patterns[56124] = 29'b1_101101100111_100_1_110110110011;
      patterns[56125] = 29'b1_101101100111_101_1_111011011001;
      patterns[56126] = 29'b1_101101100111_110_1_101101100111;
      patterns[56127] = 29'b1_101101100111_111_1_101101100111;
      patterns[56128] = 29'b1_101101101000_000_1_101101101000;
      patterns[56129] = 29'b1_101101101000_001_1_101000101101;
      patterns[56130] = 29'b1_101101101000_010_1_011011010001;
      patterns[56131] = 29'b1_101101101000_011_0_110110100011;
      patterns[56132] = 29'b1_101101101000_100_0_110110110100;
      patterns[56133] = 29'b1_101101101000_101_0_011011011010;
      patterns[56134] = 29'b1_101101101000_110_1_101101101000;
      patterns[56135] = 29'b1_101101101000_111_1_101101101000;
      patterns[56136] = 29'b1_101101101001_000_1_101101101001;
      patterns[56137] = 29'b1_101101101001_001_1_101001101101;
      patterns[56138] = 29'b1_101101101001_010_1_011011010011;
      patterns[56139] = 29'b1_101101101001_011_0_110110100111;
      patterns[56140] = 29'b1_101101101001_100_1_110110110100;
      patterns[56141] = 29'b1_101101101001_101_0_111011011010;
      patterns[56142] = 29'b1_101101101001_110_1_101101101001;
      patterns[56143] = 29'b1_101101101001_111_1_101101101001;
      patterns[56144] = 29'b1_101101101010_000_1_101101101010;
      patterns[56145] = 29'b1_101101101010_001_1_101010101101;
      patterns[56146] = 29'b1_101101101010_010_1_011011010101;
      patterns[56147] = 29'b1_101101101010_011_0_110110101011;
      patterns[56148] = 29'b1_101101101010_100_0_110110110101;
      patterns[56149] = 29'b1_101101101010_101_1_011011011010;
      patterns[56150] = 29'b1_101101101010_110_1_101101101010;
      patterns[56151] = 29'b1_101101101010_111_1_101101101010;
      patterns[56152] = 29'b1_101101101011_000_1_101101101011;
      patterns[56153] = 29'b1_101101101011_001_1_101011101101;
      patterns[56154] = 29'b1_101101101011_010_1_011011010111;
      patterns[56155] = 29'b1_101101101011_011_0_110110101111;
      patterns[56156] = 29'b1_101101101011_100_1_110110110101;
      patterns[56157] = 29'b1_101101101011_101_1_111011011010;
      patterns[56158] = 29'b1_101101101011_110_1_101101101011;
      patterns[56159] = 29'b1_101101101011_111_1_101101101011;
      patterns[56160] = 29'b1_101101101100_000_1_101101101100;
      patterns[56161] = 29'b1_101101101100_001_1_101100101101;
      patterns[56162] = 29'b1_101101101100_010_1_011011011001;
      patterns[56163] = 29'b1_101101101100_011_0_110110110011;
      patterns[56164] = 29'b1_101101101100_100_0_110110110110;
      patterns[56165] = 29'b1_101101101100_101_0_011011011011;
      patterns[56166] = 29'b1_101101101100_110_1_101101101100;
      patterns[56167] = 29'b1_101101101100_111_1_101101101100;
      patterns[56168] = 29'b1_101101101101_000_1_101101101101;
      patterns[56169] = 29'b1_101101101101_001_1_101101101101;
      patterns[56170] = 29'b1_101101101101_010_1_011011011011;
      patterns[56171] = 29'b1_101101101101_011_0_110110110111;
      patterns[56172] = 29'b1_101101101101_100_1_110110110110;
      patterns[56173] = 29'b1_101101101101_101_0_111011011011;
      patterns[56174] = 29'b1_101101101101_110_1_101101101101;
      patterns[56175] = 29'b1_101101101101_111_1_101101101101;
      patterns[56176] = 29'b1_101101101110_000_1_101101101110;
      patterns[56177] = 29'b1_101101101110_001_1_101110101101;
      patterns[56178] = 29'b1_101101101110_010_1_011011011101;
      patterns[56179] = 29'b1_101101101110_011_0_110110111011;
      patterns[56180] = 29'b1_101101101110_100_0_110110110111;
      patterns[56181] = 29'b1_101101101110_101_1_011011011011;
      patterns[56182] = 29'b1_101101101110_110_1_101101101110;
      patterns[56183] = 29'b1_101101101110_111_1_101101101110;
      patterns[56184] = 29'b1_101101101111_000_1_101101101111;
      patterns[56185] = 29'b1_101101101111_001_1_101111101101;
      patterns[56186] = 29'b1_101101101111_010_1_011011011111;
      patterns[56187] = 29'b1_101101101111_011_0_110110111111;
      patterns[56188] = 29'b1_101101101111_100_1_110110110111;
      patterns[56189] = 29'b1_101101101111_101_1_111011011011;
      patterns[56190] = 29'b1_101101101111_110_1_101101101111;
      patterns[56191] = 29'b1_101101101111_111_1_101101101111;
      patterns[56192] = 29'b1_101101110000_000_1_101101110000;
      patterns[56193] = 29'b1_101101110000_001_1_110000101101;
      patterns[56194] = 29'b1_101101110000_010_1_011011100001;
      patterns[56195] = 29'b1_101101110000_011_0_110111000011;
      patterns[56196] = 29'b1_101101110000_100_0_110110111000;
      patterns[56197] = 29'b1_101101110000_101_0_011011011100;
      patterns[56198] = 29'b1_101101110000_110_1_101101110000;
      patterns[56199] = 29'b1_101101110000_111_1_101101110000;
      patterns[56200] = 29'b1_101101110001_000_1_101101110001;
      patterns[56201] = 29'b1_101101110001_001_1_110001101101;
      patterns[56202] = 29'b1_101101110001_010_1_011011100011;
      patterns[56203] = 29'b1_101101110001_011_0_110111000111;
      patterns[56204] = 29'b1_101101110001_100_1_110110111000;
      patterns[56205] = 29'b1_101101110001_101_0_111011011100;
      patterns[56206] = 29'b1_101101110001_110_1_101101110001;
      patterns[56207] = 29'b1_101101110001_111_1_101101110001;
      patterns[56208] = 29'b1_101101110010_000_1_101101110010;
      patterns[56209] = 29'b1_101101110010_001_1_110010101101;
      patterns[56210] = 29'b1_101101110010_010_1_011011100101;
      patterns[56211] = 29'b1_101101110010_011_0_110111001011;
      patterns[56212] = 29'b1_101101110010_100_0_110110111001;
      patterns[56213] = 29'b1_101101110010_101_1_011011011100;
      patterns[56214] = 29'b1_101101110010_110_1_101101110010;
      patterns[56215] = 29'b1_101101110010_111_1_101101110010;
      patterns[56216] = 29'b1_101101110011_000_1_101101110011;
      patterns[56217] = 29'b1_101101110011_001_1_110011101101;
      patterns[56218] = 29'b1_101101110011_010_1_011011100111;
      patterns[56219] = 29'b1_101101110011_011_0_110111001111;
      patterns[56220] = 29'b1_101101110011_100_1_110110111001;
      patterns[56221] = 29'b1_101101110011_101_1_111011011100;
      patterns[56222] = 29'b1_101101110011_110_1_101101110011;
      patterns[56223] = 29'b1_101101110011_111_1_101101110011;
      patterns[56224] = 29'b1_101101110100_000_1_101101110100;
      patterns[56225] = 29'b1_101101110100_001_1_110100101101;
      patterns[56226] = 29'b1_101101110100_010_1_011011101001;
      patterns[56227] = 29'b1_101101110100_011_0_110111010011;
      patterns[56228] = 29'b1_101101110100_100_0_110110111010;
      patterns[56229] = 29'b1_101101110100_101_0_011011011101;
      patterns[56230] = 29'b1_101101110100_110_1_101101110100;
      patterns[56231] = 29'b1_101101110100_111_1_101101110100;
      patterns[56232] = 29'b1_101101110101_000_1_101101110101;
      patterns[56233] = 29'b1_101101110101_001_1_110101101101;
      patterns[56234] = 29'b1_101101110101_010_1_011011101011;
      patterns[56235] = 29'b1_101101110101_011_0_110111010111;
      patterns[56236] = 29'b1_101101110101_100_1_110110111010;
      patterns[56237] = 29'b1_101101110101_101_0_111011011101;
      patterns[56238] = 29'b1_101101110101_110_1_101101110101;
      patterns[56239] = 29'b1_101101110101_111_1_101101110101;
      patterns[56240] = 29'b1_101101110110_000_1_101101110110;
      patterns[56241] = 29'b1_101101110110_001_1_110110101101;
      patterns[56242] = 29'b1_101101110110_010_1_011011101101;
      patterns[56243] = 29'b1_101101110110_011_0_110111011011;
      patterns[56244] = 29'b1_101101110110_100_0_110110111011;
      patterns[56245] = 29'b1_101101110110_101_1_011011011101;
      patterns[56246] = 29'b1_101101110110_110_1_101101110110;
      patterns[56247] = 29'b1_101101110110_111_1_101101110110;
      patterns[56248] = 29'b1_101101110111_000_1_101101110111;
      patterns[56249] = 29'b1_101101110111_001_1_110111101101;
      patterns[56250] = 29'b1_101101110111_010_1_011011101111;
      patterns[56251] = 29'b1_101101110111_011_0_110111011111;
      patterns[56252] = 29'b1_101101110111_100_1_110110111011;
      patterns[56253] = 29'b1_101101110111_101_1_111011011101;
      patterns[56254] = 29'b1_101101110111_110_1_101101110111;
      patterns[56255] = 29'b1_101101110111_111_1_101101110111;
      patterns[56256] = 29'b1_101101111000_000_1_101101111000;
      patterns[56257] = 29'b1_101101111000_001_1_111000101101;
      patterns[56258] = 29'b1_101101111000_010_1_011011110001;
      patterns[56259] = 29'b1_101101111000_011_0_110111100011;
      patterns[56260] = 29'b1_101101111000_100_0_110110111100;
      patterns[56261] = 29'b1_101101111000_101_0_011011011110;
      patterns[56262] = 29'b1_101101111000_110_1_101101111000;
      patterns[56263] = 29'b1_101101111000_111_1_101101111000;
      patterns[56264] = 29'b1_101101111001_000_1_101101111001;
      patterns[56265] = 29'b1_101101111001_001_1_111001101101;
      patterns[56266] = 29'b1_101101111001_010_1_011011110011;
      patterns[56267] = 29'b1_101101111001_011_0_110111100111;
      patterns[56268] = 29'b1_101101111001_100_1_110110111100;
      patterns[56269] = 29'b1_101101111001_101_0_111011011110;
      patterns[56270] = 29'b1_101101111001_110_1_101101111001;
      patterns[56271] = 29'b1_101101111001_111_1_101101111001;
      patterns[56272] = 29'b1_101101111010_000_1_101101111010;
      patterns[56273] = 29'b1_101101111010_001_1_111010101101;
      patterns[56274] = 29'b1_101101111010_010_1_011011110101;
      patterns[56275] = 29'b1_101101111010_011_0_110111101011;
      patterns[56276] = 29'b1_101101111010_100_0_110110111101;
      patterns[56277] = 29'b1_101101111010_101_1_011011011110;
      patterns[56278] = 29'b1_101101111010_110_1_101101111010;
      patterns[56279] = 29'b1_101101111010_111_1_101101111010;
      patterns[56280] = 29'b1_101101111011_000_1_101101111011;
      patterns[56281] = 29'b1_101101111011_001_1_111011101101;
      patterns[56282] = 29'b1_101101111011_010_1_011011110111;
      patterns[56283] = 29'b1_101101111011_011_0_110111101111;
      patterns[56284] = 29'b1_101101111011_100_1_110110111101;
      patterns[56285] = 29'b1_101101111011_101_1_111011011110;
      patterns[56286] = 29'b1_101101111011_110_1_101101111011;
      patterns[56287] = 29'b1_101101111011_111_1_101101111011;
      patterns[56288] = 29'b1_101101111100_000_1_101101111100;
      patterns[56289] = 29'b1_101101111100_001_1_111100101101;
      patterns[56290] = 29'b1_101101111100_010_1_011011111001;
      patterns[56291] = 29'b1_101101111100_011_0_110111110011;
      patterns[56292] = 29'b1_101101111100_100_0_110110111110;
      patterns[56293] = 29'b1_101101111100_101_0_011011011111;
      patterns[56294] = 29'b1_101101111100_110_1_101101111100;
      patterns[56295] = 29'b1_101101111100_111_1_101101111100;
      patterns[56296] = 29'b1_101101111101_000_1_101101111101;
      patterns[56297] = 29'b1_101101111101_001_1_111101101101;
      patterns[56298] = 29'b1_101101111101_010_1_011011111011;
      patterns[56299] = 29'b1_101101111101_011_0_110111110111;
      patterns[56300] = 29'b1_101101111101_100_1_110110111110;
      patterns[56301] = 29'b1_101101111101_101_0_111011011111;
      patterns[56302] = 29'b1_101101111101_110_1_101101111101;
      patterns[56303] = 29'b1_101101111101_111_1_101101111101;
      patterns[56304] = 29'b1_101101111110_000_1_101101111110;
      patterns[56305] = 29'b1_101101111110_001_1_111110101101;
      patterns[56306] = 29'b1_101101111110_010_1_011011111101;
      patterns[56307] = 29'b1_101101111110_011_0_110111111011;
      patterns[56308] = 29'b1_101101111110_100_0_110110111111;
      patterns[56309] = 29'b1_101101111110_101_1_011011011111;
      patterns[56310] = 29'b1_101101111110_110_1_101101111110;
      patterns[56311] = 29'b1_101101111110_111_1_101101111110;
      patterns[56312] = 29'b1_101101111111_000_1_101101111111;
      patterns[56313] = 29'b1_101101111111_001_1_111111101101;
      patterns[56314] = 29'b1_101101111111_010_1_011011111111;
      patterns[56315] = 29'b1_101101111111_011_0_110111111111;
      patterns[56316] = 29'b1_101101111111_100_1_110110111111;
      patterns[56317] = 29'b1_101101111111_101_1_111011011111;
      patterns[56318] = 29'b1_101101111111_110_1_101101111111;
      patterns[56319] = 29'b1_101101111111_111_1_101101111111;
      patterns[56320] = 29'b1_101110000000_000_1_101110000000;
      patterns[56321] = 29'b1_101110000000_001_1_000000101110;
      patterns[56322] = 29'b1_101110000000_010_1_011100000001;
      patterns[56323] = 29'b1_101110000000_011_0_111000000011;
      patterns[56324] = 29'b1_101110000000_100_0_110111000000;
      patterns[56325] = 29'b1_101110000000_101_0_011011100000;
      patterns[56326] = 29'b1_101110000000_110_1_101110000000;
      patterns[56327] = 29'b1_101110000000_111_1_101110000000;
      patterns[56328] = 29'b1_101110000001_000_1_101110000001;
      patterns[56329] = 29'b1_101110000001_001_1_000001101110;
      patterns[56330] = 29'b1_101110000001_010_1_011100000011;
      patterns[56331] = 29'b1_101110000001_011_0_111000000111;
      patterns[56332] = 29'b1_101110000001_100_1_110111000000;
      patterns[56333] = 29'b1_101110000001_101_0_111011100000;
      patterns[56334] = 29'b1_101110000001_110_1_101110000001;
      patterns[56335] = 29'b1_101110000001_111_1_101110000001;
      patterns[56336] = 29'b1_101110000010_000_1_101110000010;
      patterns[56337] = 29'b1_101110000010_001_1_000010101110;
      patterns[56338] = 29'b1_101110000010_010_1_011100000101;
      patterns[56339] = 29'b1_101110000010_011_0_111000001011;
      patterns[56340] = 29'b1_101110000010_100_0_110111000001;
      patterns[56341] = 29'b1_101110000010_101_1_011011100000;
      patterns[56342] = 29'b1_101110000010_110_1_101110000010;
      patterns[56343] = 29'b1_101110000010_111_1_101110000010;
      patterns[56344] = 29'b1_101110000011_000_1_101110000011;
      patterns[56345] = 29'b1_101110000011_001_1_000011101110;
      patterns[56346] = 29'b1_101110000011_010_1_011100000111;
      patterns[56347] = 29'b1_101110000011_011_0_111000001111;
      patterns[56348] = 29'b1_101110000011_100_1_110111000001;
      patterns[56349] = 29'b1_101110000011_101_1_111011100000;
      patterns[56350] = 29'b1_101110000011_110_1_101110000011;
      patterns[56351] = 29'b1_101110000011_111_1_101110000011;
      patterns[56352] = 29'b1_101110000100_000_1_101110000100;
      patterns[56353] = 29'b1_101110000100_001_1_000100101110;
      patterns[56354] = 29'b1_101110000100_010_1_011100001001;
      patterns[56355] = 29'b1_101110000100_011_0_111000010011;
      patterns[56356] = 29'b1_101110000100_100_0_110111000010;
      patterns[56357] = 29'b1_101110000100_101_0_011011100001;
      patterns[56358] = 29'b1_101110000100_110_1_101110000100;
      patterns[56359] = 29'b1_101110000100_111_1_101110000100;
      patterns[56360] = 29'b1_101110000101_000_1_101110000101;
      patterns[56361] = 29'b1_101110000101_001_1_000101101110;
      patterns[56362] = 29'b1_101110000101_010_1_011100001011;
      patterns[56363] = 29'b1_101110000101_011_0_111000010111;
      patterns[56364] = 29'b1_101110000101_100_1_110111000010;
      patterns[56365] = 29'b1_101110000101_101_0_111011100001;
      patterns[56366] = 29'b1_101110000101_110_1_101110000101;
      patterns[56367] = 29'b1_101110000101_111_1_101110000101;
      patterns[56368] = 29'b1_101110000110_000_1_101110000110;
      patterns[56369] = 29'b1_101110000110_001_1_000110101110;
      patterns[56370] = 29'b1_101110000110_010_1_011100001101;
      patterns[56371] = 29'b1_101110000110_011_0_111000011011;
      patterns[56372] = 29'b1_101110000110_100_0_110111000011;
      patterns[56373] = 29'b1_101110000110_101_1_011011100001;
      patterns[56374] = 29'b1_101110000110_110_1_101110000110;
      patterns[56375] = 29'b1_101110000110_111_1_101110000110;
      patterns[56376] = 29'b1_101110000111_000_1_101110000111;
      patterns[56377] = 29'b1_101110000111_001_1_000111101110;
      patterns[56378] = 29'b1_101110000111_010_1_011100001111;
      patterns[56379] = 29'b1_101110000111_011_0_111000011111;
      patterns[56380] = 29'b1_101110000111_100_1_110111000011;
      patterns[56381] = 29'b1_101110000111_101_1_111011100001;
      patterns[56382] = 29'b1_101110000111_110_1_101110000111;
      patterns[56383] = 29'b1_101110000111_111_1_101110000111;
      patterns[56384] = 29'b1_101110001000_000_1_101110001000;
      patterns[56385] = 29'b1_101110001000_001_1_001000101110;
      patterns[56386] = 29'b1_101110001000_010_1_011100010001;
      patterns[56387] = 29'b1_101110001000_011_0_111000100011;
      patterns[56388] = 29'b1_101110001000_100_0_110111000100;
      patterns[56389] = 29'b1_101110001000_101_0_011011100010;
      patterns[56390] = 29'b1_101110001000_110_1_101110001000;
      patterns[56391] = 29'b1_101110001000_111_1_101110001000;
      patterns[56392] = 29'b1_101110001001_000_1_101110001001;
      patterns[56393] = 29'b1_101110001001_001_1_001001101110;
      patterns[56394] = 29'b1_101110001001_010_1_011100010011;
      patterns[56395] = 29'b1_101110001001_011_0_111000100111;
      patterns[56396] = 29'b1_101110001001_100_1_110111000100;
      patterns[56397] = 29'b1_101110001001_101_0_111011100010;
      patterns[56398] = 29'b1_101110001001_110_1_101110001001;
      patterns[56399] = 29'b1_101110001001_111_1_101110001001;
      patterns[56400] = 29'b1_101110001010_000_1_101110001010;
      patterns[56401] = 29'b1_101110001010_001_1_001010101110;
      patterns[56402] = 29'b1_101110001010_010_1_011100010101;
      patterns[56403] = 29'b1_101110001010_011_0_111000101011;
      patterns[56404] = 29'b1_101110001010_100_0_110111000101;
      patterns[56405] = 29'b1_101110001010_101_1_011011100010;
      patterns[56406] = 29'b1_101110001010_110_1_101110001010;
      patterns[56407] = 29'b1_101110001010_111_1_101110001010;
      patterns[56408] = 29'b1_101110001011_000_1_101110001011;
      patterns[56409] = 29'b1_101110001011_001_1_001011101110;
      patterns[56410] = 29'b1_101110001011_010_1_011100010111;
      patterns[56411] = 29'b1_101110001011_011_0_111000101111;
      patterns[56412] = 29'b1_101110001011_100_1_110111000101;
      patterns[56413] = 29'b1_101110001011_101_1_111011100010;
      patterns[56414] = 29'b1_101110001011_110_1_101110001011;
      patterns[56415] = 29'b1_101110001011_111_1_101110001011;
      patterns[56416] = 29'b1_101110001100_000_1_101110001100;
      patterns[56417] = 29'b1_101110001100_001_1_001100101110;
      patterns[56418] = 29'b1_101110001100_010_1_011100011001;
      patterns[56419] = 29'b1_101110001100_011_0_111000110011;
      patterns[56420] = 29'b1_101110001100_100_0_110111000110;
      patterns[56421] = 29'b1_101110001100_101_0_011011100011;
      patterns[56422] = 29'b1_101110001100_110_1_101110001100;
      patterns[56423] = 29'b1_101110001100_111_1_101110001100;
      patterns[56424] = 29'b1_101110001101_000_1_101110001101;
      patterns[56425] = 29'b1_101110001101_001_1_001101101110;
      patterns[56426] = 29'b1_101110001101_010_1_011100011011;
      patterns[56427] = 29'b1_101110001101_011_0_111000110111;
      patterns[56428] = 29'b1_101110001101_100_1_110111000110;
      patterns[56429] = 29'b1_101110001101_101_0_111011100011;
      patterns[56430] = 29'b1_101110001101_110_1_101110001101;
      patterns[56431] = 29'b1_101110001101_111_1_101110001101;
      patterns[56432] = 29'b1_101110001110_000_1_101110001110;
      patterns[56433] = 29'b1_101110001110_001_1_001110101110;
      patterns[56434] = 29'b1_101110001110_010_1_011100011101;
      patterns[56435] = 29'b1_101110001110_011_0_111000111011;
      patterns[56436] = 29'b1_101110001110_100_0_110111000111;
      patterns[56437] = 29'b1_101110001110_101_1_011011100011;
      patterns[56438] = 29'b1_101110001110_110_1_101110001110;
      patterns[56439] = 29'b1_101110001110_111_1_101110001110;
      patterns[56440] = 29'b1_101110001111_000_1_101110001111;
      patterns[56441] = 29'b1_101110001111_001_1_001111101110;
      patterns[56442] = 29'b1_101110001111_010_1_011100011111;
      patterns[56443] = 29'b1_101110001111_011_0_111000111111;
      patterns[56444] = 29'b1_101110001111_100_1_110111000111;
      patterns[56445] = 29'b1_101110001111_101_1_111011100011;
      patterns[56446] = 29'b1_101110001111_110_1_101110001111;
      patterns[56447] = 29'b1_101110001111_111_1_101110001111;
      patterns[56448] = 29'b1_101110010000_000_1_101110010000;
      patterns[56449] = 29'b1_101110010000_001_1_010000101110;
      patterns[56450] = 29'b1_101110010000_010_1_011100100001;
      patterns[56451] = 29'b1_101110010000_011_0_111001000011;
      patterns[56452] = 29'b1_101110010000_100_0_110111001000;
      patterns[56453] = 29'b1_101110010000_101_0_011011100100;
      patterns[56454] = 29'b1_101110010000_110_1_101110010000;
      patterns[56455] = 29'b1_101110010000_111_1_101110010000;
      patterns[56456] = 29'b1_101110010001_000_1_101110010001;
      patterns[56457] = 29'b1_101110010001_001_1_010001101110;
      patterns[56458] = 29'b1_101110010001_010_1_011100100011;
      patterns[56459] = 29'b1_101110010001_011_0_111001000111;
      patterns[56460] = 29'b1_101110010001_100_1_110111001000;
      patterns[56461] = 29'b1_101110010001_101_0_111011100100;
      patterns[56462] = 29'b1_101110010001_110_1_101110010001;
      patterns[56463] = 29'b1_101110010001_111_1_101110010001;
      patterns[56464] = 29'b1_101110010010_000_1_101110010010;
      patterns[56465] = 29'b1_101110010010_001_1_010010101110;
      patterns[56466] = 29'b1_101110010010_010_1_011100100101;
      patterns[56467] = 29'b1_101110010010_011_0_111001001011;
      patterns[56468] = 29'b1_101110010010_100_0_110111001001;
      patterns[56469] = 29'b1_101110010010_101_1_011011100100;
      patterns[56470] = 29'b1_101110010010_110_1_101110010010;
      patterns[56471] = 29'b1_101110010010_111_1_101110010010;
      patterns[56472] = 29'b1_101110010011_000_1_101110010011;
      patterns[56473] = 29'b1_101110010011_001_1_010011101110;
      patterns[56474] = 29'b1_101110010011_010_1_011100100111;
      patterns[56475] = 29'b1_101110010011_011_0_111001001111;
      patterns[56476] = 29'b1_101110010011_100_1_110111001001;
      patterns[56477] = 29'b1_101110010011_101_1_111011100100;
      patterns[56478] = 29'b1_101110010011_110_1_101110010011;
      patterns[56479] = 29'b1_101110010011_111_1_101110010011;
      patterns[56480] = 29'b1_101110010100_000_1_101110010100;
      patterns[56481] = 29'b1_101110010100_001_1_010100101110;
      patterns[56482] = 29'b1_101110010100_010_1_011100101001;
      patterns[56483] = 29'b1_101110010100_011_0_111001010011;
      patterns[56484] = 29'b1_101110010100_100_0_110111001010;
      patterns[56485] = 29'b1_101110010100_101_0_011011100101;
      patterns[56486] = 29'b1_101110010100_110_1_101110010100;
      patterns[56487] = 29'b1_101110010100_111_1_101110010100;
      patterns[56488] = 29'b1_101110010101_000_1_101110010101;
      patterns[56489] = 29'b1_101110010101_001_1_010101101110;
      patterns[56490] = 29'b1_101110010101_010_1_011100101011;
      patterns[56491] = 29'b1_101110010101_011_0_111001010111;
      patterns[56492] = 29'b1_101110010101_100_1_110111001010;
      patterns[56493] = 29'b1_101110010101_101_0_111011100101;
      patterns[56494] = 29'b1_101110010101_110_1_101110010101;
      patterns[56495] = 29'b1_101110010101_111_1_101110010101;
      patterns[56496] = 29'b1_101110010110_000_1_101110010110;
      patterns[56497] = 29'b1_101110010110_001_1_010110101110;
      patterns[56498] = 29'b1_101110010110_010_1_011100101101;
      patterns[56499] = 29'b1_101110010110_011_0_111001011011;
      patterns[56500] = 29'b1_101110010110_100_0_110111001011;
      patterns[56501] = 29'b1_101110010110_101_1_011011100101;
      patterns[56502] = 29'b1_101110010110_110_1_101110010110;
      patterns[56503] = 29'b1_101110010110_111_1_101110010110;
      patterns[56504] = 29'b1_101110010111_000_1_101110010111;
      patterns[56505] = 29'b1_101110010111_001_1_010111101110;
      patterns[56506] = 29'b1_101110010111_010_1_011100101111;
      patterns[56507] = 29'b1_101110010111_011_0_111001011111;
      patterns[56508] = 29'b1_101110010111_100_1_110111001011;
      patterns[56509] = 29'b1_101110010111_101_1_111011100101;
      patterns[56510] = 29'b1_101110010111_110_1_101110010111;
      patterns[56511] = 29'b1_101110010111_111_1_101110010111;
      patterns[56512] = 29'b1_101110011000_000_1_101110011000;
      patterns[56513] = 29'b1_101110011000_001_1_011000101110;
      patterns[56514] = 29'b1_101110011000_010_1_011100110001;
      patterns[56515] = 29'b1_101110011000_011_0_111001100011;
      patterns[56516] = 29'b1_101110011000_100_0_110111001100;
      patterns[56517] = 29'b1_101110011000_101_0_011011100110;
      patterns[56518] = 29'b1_101110011000_110_1_101110011000;
      patterns[56519] = 29'b1_101110011000_111_1_101110011000;
      patterns[56520] = 29'b1_101110011001_000_1_101110011001;
      patterns[56521] = 29'b1_101110011001_001_1_011001101110;
      patterns[56522] = 29'b1_101110011001_010_1_011100110011;
      patterns[56523] = 29'b1_101110011001_011_0_111001100111;
      patterns[56524] = 29'b1_101110011001_100_1_110111001100;
      patterns[56525] = 29'b1_101110011001_101_0_111011100110;
      patterns[56526] = 29'b1_101110011001_110_1_101110011001;
      patterns[56527] = 29'b1_101110011001_111_1_101110011001;
      patterns[56528] = 29'b1_101110011010_000_1_101110011010;
      patterns[56529] = 29'b1_101110011010_001_1_011010101110;
      patterns[56530] = 29'b1_101110011010_010_1_011100110101;
      patterns[56531] = 29'b1_101110011010_011_0_111001101011;
      patterns[56532] = 29'b1_101110011010_100_0_110111001101;
      patterns[56533] = 29'b1_101110011010_101_1_011011100110;
      patterns[56534] = 29'b1_101110011010_110_1_101110011010;
      patterns[56535] = 29'b1_101110011010_111_1_101110011010;
      patterns[56536] = 29'b1_101110011011_000_1_101110011011;
      patterns[56537] = 29'b1_101110011011_001_1_011011101110;
      patterns[56538] = 29'b1_101110011011_010_1_011100110111;
      patterns[56539] = 29'b1_101110011011_011_0_111001101111;
      patterns[56540] = 29'b1_101110011011_100_1_110111001101;
      patterns[56541] = 29'b1_101110011011_101_1_111011100110;
      patterns[56542] = 29'b1_101110011011_110_1_101110011011;
      patterns[56543] = 29'b1_101110011011_111_1_101110011011;
      patterns[56544] = 29'b1_101110011100_000_1_101110011100;
      patterns[56545] = 29'b1_101110011100_001_1_011100101110;
      patterns[56546] = 29'b1_101110011100_010_1_011100111001;
      patterns[56547] = 29'b1_101110011100_011_0_111001110011;
      patterns[56548] = 29'b1_101110011100_100_0_110111001110;
      patterns[56549] = 29'b1_101110011100_101_0_011011100111;
      patterns[56550] = 29'b1_101110011100_110_1_101110011100;
      patterns[56551] = 29'b1_101110011100_111_1_101110011100;
      patterns[56552] = 29'b1_101110011101_000_1_101110011101;
      patterns[56553] = 29'b1_101110011101_001_1_011101101110;
      patterns[56554] = 29'b1_101110011101_010_1_011100111011;
      patterns[56555] = 29'b1_101110011101_011_0_111001110111;
      patterns[56556] = 29'b1_101110011101_100_1_110111001110;
      patterns[56557] = 29'b1_101110011101_101_0_111011100111;
      patterns[56558] = 29'b1_101110011101_110_1_101110011101;
      patterns[56559] = 29'b1_101110011101_111_1_101110011101;
      patterns[56560] = 29'b1_101110011110_000_1_101110011110;
      patterns[56561] = 29'b1_101110011110_001_1_011110101110;
      patterns[56562] = 29'b1_101110011110_010_1_011100111101;
      patterns[56563] = 29'b1_101110011110_011_0_111001111011;
      patterns[56564] = 29'b1_101110011110_100_0_110111001111;
      patterns[56565] = 29'b1_101110011110_101_1_011011100111;
      patterns[56566] = 29'b1_101110011110_110_1_101110011110;
      patterns[56567] = 29'b1_101110011110_111_1_101110011110;
      patterns[56568] = 29'b1_101110011111_000_1_101110011111;
      patterns[56569] = 29'b1_101110011111_001_1_011111101110;
      patterns[56570] = 29'b1_101110011111_010_1_011100111111;
      patterns[56571] = 29'b1_101110011111_011_0_111001111111;
      patterns[56572] = 29'b1_101110011111_100_1_110111001111;
      patterns[56573] = 29'b1_101110011111_101_1_111011100111;
      patterns[56574] = 29'b1_101110011111_110_1_101110011111;
      patterns[56575] = 29'b1_101110011111_111_1_101110011111;
      patterns[56576] = 29'b1_101110100000_000_1_101110100000;
      patterns[56577] = 29'b1_101110100000_001_1_100000101110;
      patterns[56578] = 29'b1_101110100000_010_1_011101000001;
      patterns[56579] = 29'b1_101110100000_011_0_111010000011;
      patterns[56580] = 29'b1_101110100000_100_0_110111010000;
      patterns[56581] = 29'b1_101110100000_101_0_011011101000;
      patterns[56582] = 29'b1_101110100000_110_1_101110100000;
      patterns[56583] = 29'b1_101110100000_111_1_101110100000;
      patterns[56584] = 29'b1_101110100001_000_1_101110100001;
      patterns[56585] = 29'b1_101110100001_001_1_100001101110;
      patterns[56586] = 29'b1_101110100001_010_1_011101000011;
      patterns[56587] = 29'b1_101110100001_011_0_111010000111;
      patterns[56588] = 29'b1_101110100001_100_1_110111010000;
      patterns[56589] = 29'b1_101110100001_101_0_111011101000;
      patterns[56590] = 29'b1_101110100001_110_1_101110100001;
      patterns[56591] = 29'b1_101110100001_111_1_101110100001;
      patterns[56592] = 29'b1_101110100010_000_1_101110100010;
      patterns[56593] = 29'b1_101110100010_001_1_100010101110;
      patterns[56594] = 29'b1_101110100010_010_1_011101000101;
      patterns[56595] = 29'b1_101110100010_011_0_111010001011;
      patterns[56596] = 29'b1_101110100010_100_0_110111010001;
      patterns[56597] = 29'b1_101110100010_101_1_011011101000;
      patterns[56598] = 29'b1_101110100010_110_1_101110100010;
      patterns[56599] = 29'b1_101110100010_111_1_101110100010;
      patterns[56600] = 29'b1_101110100011_000_1_101110100011;
      patterns[56601] = 29'b1_101110100011_001_1_100011101110;
      patterns[56602] = 29'b1_101110100011_010_1_011101000111;
      patterns[56603] = 29'b1_101110100011_011_0_111010001111;
      patterns[56604] = 29'b1_101110100011_100_1_110111010001;
      patterns[56605] = 29'b1_101110100011_101_1_111011101000;
      patterns[56606] = 29'b1_101110100011_110_1_101110100011;
      patterns[56607] = 29'b1_101110100011_111_1_101110100011;
      patterns[56608] = 29'b1_101110100100_000_1_101110100100;
      patterns[56609] = 29'b1_101110100100_001_1_100100101110;
      patterns[56610] = 29'b1_101110100100_010_1_011101001001;
      patterns[56611] = 29'b1_101110100100_011_0_111010010011;
      patterns[56612] = 29'b1_101110100100_100_0_110111010010;
      patterns[56613] = 29'b1_101110100100_101_0_011011101001;
      patterns[56614] = 29'b1_101110100100_110_1_101110100100;
      patterns[56615] = 29'b1_101110100100_111_1_101110100100;
      patterns[56616] = 29'b1_101110100101_000_1_101110100101;
      patterns[56617] = 29'b1_101110100101_001_1_100101101110;
      patterns[56618] = 29'b1_101110100101_010_1_011101001011;
      patterns[56619] = 29'b1_101110100101_011_0_111010010111;
      patterns[56620] = 29'b1_101110100101_100_1_110111010010;
      patterns[56621] = 29'b1_101110100101_101_0_111011101001;
      patterns[56622] = 29'b1_101110100101_110_1_101110100101;
      patterns[56623] = 29'b1_101110100101_111_1_101110100101;
      patterns[56624] = 29'b1_101110100110_000_1_101110100110;
      patterns[56625] = 29'b1_101110100110_001_1_100110101110;
      patterns[56626] = 29'b1_101110100110_010_1_011101001101;
      patterns[56627] = 29'b1_101110100110_011_0_111010011011;
      patterns[56628] = 29'b1_101110100110_100_0_110111010011;
      patterns[56629] = 29'b1_101110100110_101_1_011011101001;
      patterns[56630] = 29'b1_101110100110_110_1_101110100110;
      patterns[56631] = 29'b1_101110100110_111_1_101110100110;
      patterns[56632] = 29'b1_101110100111_000_1_101110100111;
      patterns[56633] = 29'b1_101110100111_001_1_100111101110;
      patterns[56634] = 29'b1_101110100111_010_1_011101001111;
      patterns[56635] = 29'b1_101110100111_011_0_111010011111;
      patterns[56636] = 29'b1_101110100111_100_1_110111010011;
      patterns[56637] = 29'b1_101110100111_101_1_111011101001;
      patterns[56638] = 29'b1_101110100111_110_1_101110100111;
      patterns[56639] = 29'b1_101110100111_111_1_101110100111;
      patterns[56640] = 29'b1_101110101000_000_1_101110101000;
      patterns[56641] = 29'b1_101110101000_001_1_101000101110;
      patterns[56642] = 29'b1_101110101000_010_1_011101010001;
      patterns[56643] = 29'b1_101110101000_011_0_111010100011;
      patterns[56644] = 29'b1_101110101000_100_0_110111010100;
      patterns[56645] = 29'b1_101110101000_101_0_011011101010;
      patterns[56646] = 29'b1_101110101000_110_1_101110101000;
      patterns[56647] = 29'b1_101110101000_111_1_101110101000;
      patterns[56648] = 29'b1_101110101001_000_1_101110101001;
      patterns[56649] = 29'b1_101110101001_001_1_101001101110;
      patterns[56650] = 29'b1_101110101001_010_1_011101010011;
      patterns[56651] = 29'b1_101110101001_011_0_111010100111;
      patterns[56652] = 29'b1_101110101001_100_1_110111010100;
      patterns[56653] = 29'b1_101110101001_101_0_111011101010;
      patterns[56654] = 29'b1_101110101001_110_1_101110101001;
      patterns[56655] = 29'b1_101110101001_111_1_101110101001;
      patterns[56656] = 29'b1_101110101010_000_1_101110101010;
      patterns[56657] = 29'b1_101110101010_001_1_101010101110;
      patterns[56658] = 29'b1_101110101010_010_1_011101010101;
      patterns[56659] = 29'b1_101110101010_011_0_111010101011;
      patterns[56660] = 29'b1_101110101010_100_0_110111010101;
      patterns[56661] = 29'b1_101110101010_101_1_011011101010;
      patterns[56662] = 29'b1_101110101010_110_1_101110101010;
      patterns[56663] = 29'b1_101110101010_111_1_101110101010;
      patterns[56664] = 29'b1_101110101011_000_1_101110101011;
      patterns[56665] = 29'b1_101110101011_001_1_101011101110;
      patterns[56666] = 29'b1_101110101011_010_1_011101010111;
      patterns[56667] = 29'b1_101110101011_011_0_111010101111;
      patterns[56668] = 29'b1_101110101011_100_1_110111010101;
      patterns[56669] = 29'b1_101110101011_101_1_111011101010;
      patterns[56670] = 29'b1_101110101011_110_1_101110101011;
      patterns[56671] = 29'b1_101110101011_111_1_101110101011;
      patterns[56672] = 29'b1_101110101100_000_1_101110101100;
      patterns[56673] = 29'b1_101110101100_001_1_101100101110;
      patterns[56674] = 29'b1_101110101100_010_1_011101011001;
      patterns[56675] = 29'b1_101110101100_011_0_111010110011;
      patterns[56676] = 29'b1_101110101100_100_0_110111010110;
      patterns[56677] = 29'b1_101110101100_101_0_011011101011;
      patterns[56678] = 29'b1_101110101100_110_1_101110101100;
      patterns[56679] = 29'b1_101110101100_111_1_101110101100;
      patterns[56680] = 29'b1_101110101101_000_1_101110101101;
      patterns[56681] = 29'b1_101110101101_001_1_101101101110;
      patterns[56682] = 29'b1_101110101101_010_1_011101011011;
      patterns[56683] = 29'b1_101110101101_011_0_111010110111;
      patterns[56684] = 29'b1_101110101101_100_1_110111010110;
      patterns[56685] = 29'b1_101110101101_101_0_111011101011;
      patterns[56686] = 29'b1_101110101101_110_1_101110101101;
      patterns[56687] = 29'b1_101110101101_111_1_101110101101;
      patterns[56688] = 29'b1_101110101110_000_1_101110101110;
      patterns[56689] = 29'b1_101110101110_001_1_101110101110;
      patterns[56690] = 29'b1_101110101110_010_1_011101011101;
      patterns[56691] = 29'b1_101110101110_011_0_111010111011;
      patterns[56692] = 29'b1_101110101110_100_0_110111010111;
      patterns[56693] = 29'b1_101110101110_101_1_011011101011;
      patterns[56694] = 29'b1_101110101110_110_1_101110101110;
      patterns[56695] = 29'b1_101110101110_111_1_101110101110;
      patterns[56696] = 29'b1_101110101111_000_1_101110101111;
      patterns[56697] = 29'b1_101110101111_001_1_101111101110;
      patterns[56698] = 29'b1_101110101111_010_1_011101011111;
      patterns[56699] = 29'b1_101110101111_011_0_111010111111;
      patterns[56700] = 29'b1_101110101111_100_1_110111010111;
      patterns[56701] = 29'b1_101110101111_101_1_111011101011;
      patterns[56702] = 29'b1_101110101111_110_1_101110101111;
      patterns[56703] = 29'b1_101110101111_111_1_101110101111;
      patterns[56704] = 29'b1_101110110000_000_1_101110110000;
      patterns[56705] = 29'b1_101110110000_001_1_110000101110;
      patterns[56706] = 29'b1_101110110000_010_1_011101100001;
      patterns[56707] = 29'b1_101110110000_011_0_111011000011;
      patterns[56708] = 29'b1_101110110000_100_0_110111011000;
      patterns[56709] = 29'b1_101110110000_101_0_011011101100;
      patterns[56710] = 29'b1_101110110000_110_1_101110110000;
      patterns[56711] = 29'b1_101110110000_111_1_101110110000;
      patterns[56712] = 29'b1_101110110001_000_1_101110110001;
      patterns[56713] = 29'b1_101110110001_001_1_110001101110;
      patterns[56714] = 29'b1_101110110001_010_1_011101100011;
      patterns[56715] = 29'b1_101110110001_011_0_111011000111;
      patterns[56716] = 29'b1_101110110001_100_1_110111011000;
      patterns[56717] = 29'b1_101110110001_101_0_111011101100;
      patterns[56718] = 29'b1_101110110001_110_1_101110110001;
      patterns[56719] = 29'b1_101110110001_111_1_101110110001;
      patterns[56720] = 29'b1_101110110010_000_1_101110110010;
      patterns[56721] = 29'b1_101110110010_001_1_110010101110;
      patterns[56722] = 29'b1_101110110010_010_1_011101100101;
      patterns[56723] = 29'b1_101110110010_011_0_111011001011;
      patterns[56724] = 29'b1_101110110010_100_0_110111011001;
      patterns[56725] = 29'b1_101110110010_101_1_011011101100;
      patterns[56726] = 29'b1_101110110010_110_1_101110110010;
      patterns[56727] = 29'b1_101110110010_111_1_101110110010;
      patterns[56728] = 29'b1_101110110011_000_1_101110110011;
      patterns[56729] = 29'b1_101110110011_001_1_110011101110;
      patterns[56730] = 29'b1_101110110011_010_1_011101100111;
      patterns[56731] = 29'b1_101110110011_011_0_111011001111;
      patterns[56732] = 29'b1_101110110011_100_1_110111011001;
      patterns[56733] = 29'b1_101110110011_101_1_111011101100;
      patterns[56734] = 29'b1_101110110011_110_1_101110110011;
      patterns[56735] = 29'b1_101110110011_111_1_101110110011;
      patterns[56736] = 29'b1_101110110100_000_1_101110110100;
      patterns[56737] = 29'b1_101110110100_001_1_110100101110;
      patterns[56738] = 29'b1_101110110100_010_1_011101101001;
      patterns[56739] = 29'b1_101110110100_011_0_111011010011;
      patterns[56740] = 29'b1_101110110100_100_0_110111011010;
      patterns[56741] = 29'b1_101110110100_101_0_011011101101;
      patterns[56742] = 29'b1_101110110100_110_1_101110110100;
      patterns[56743] = 29'b1_101110110100_111_1_101110110100;
      patterns[56744] = 29'b1_101110110101_000_1_101110110101;
      patterns[56745] = 29'b1_101110110101_001_1_110101101110;
      patterns[56746] = 29'b1_101110110101_010_1_011101101011;
      patterns[56747] = 29'b1_101110110101_011_0_111011010111;
      patterns[56748] = 29'b1_101110110101_100_1_110111011010;
      patterns[56749] = 29'b1_101110110101_101_0_111011101101;
      patterns[56750] = 29'b1_101110110101_110_1_101110110101;
      patterns[56751] = 29'b1_101110110101_111_1_101110110101;
      patterns[56752] = 29'b1_101110110110_000_1_101110110110;
      patterns[56753] = 29'b1_101110110110_001_1_110110101110;
      patterns[56754] = 29'b1_101110110110_010_1_011101101101;
      patterns[56755] = 29'b1_101110110110_011_0_111011011011;
      patterns[56756] = 29'b1_101110110110_100_0_110111011011;
      patterns[56757] = 29'b1_101110110110_101_1_011011101101;
      patterns[56758] = 29'b1_101110110110_110_1_101110110110;
      patterns[56759] = 29'b1_101110110110_111_1_101110110110;
      patterns[56760] = 29'b1_101110110111_000_1_101110110111;
      patterns[56761] = 29'b1_101110110111_001_1_110111101110;
      patterns[56762] = 29'b1_101110110111_010_1_011101101111;
      patterns[56763] = 29'b1_101110110111_011_0_111011011111;
      patterns[56764] = 29'b1_101110110111_100_1_110111011011;
      patterns[56765] = 29'b1_101110110111_101_1_111011101101;
      patterns[56766] = 29'b1_101110110111_110_1_101110110111;
      patterns[56767] = 29'b1_101110110111_111_1_101110110111;
      patterns[56768] = 29'b1_101110111000_000_1_101110111000;
      patterns[56769] = 29'b1_101110111000_001_1_111000101110;
      patterns[56770] = 29'b1_101110111000_010_1_011101110001;
      patterns[56771] = 29'b1_101110111000_011_0_111011100011;
      patterns[56772] = 29'b1_101110111000_100_0_110111011100;
      patterns[56773] = 29'b1_101110111000_101_0_011011101110;
      patterns[56774] = 29'b1_101110111000_110_1_101110111000;
      patterns[56775] = 29'b1_101110111000_111_1_101110111000;
      patterns[56776] = 29'b1_101110111001_000_1_101110111001;
      patterns[56777] = 29'b1_101110111001_001_1_111001101110;
      patterns[56778] = 29'b1_101110111001_010_1_011101110011;
      patterns[56779] = 29'b1_101110111001_011_0_111011100111;
      patterns[56780] = 29'b1_101110111001_100_1_110111011100;
      patterns[56781] = 29'b1_101110111001_101_0_111011101110;
      patterns[56782] = 29'b1_101110111001_110_1_101110111001;
      patterns[56783] = 29'b1_101110111001_111_1_101110111001;
      patterns[56784] = 29'b1_101110111010_000_1_101110111010;
      patterns[56785] = 29'b1_101110111010_001_1_111010101110;
      patterns[56786] = 29'b1_101110111010_010_1_011101110101;
      patterns[56787] = 29'b1_101110111010_011_0_111011101011;
      patterns[56788] = 29'b1_101110111010_100_0_110111011101;
      patterns[56789] = 29'b1_101110111010_101_1_011011101110;
      patterns[56790] = 29'b1_101110111010_110_1_101110111010;
      patterns[56791] = 29'b1_101110111010_111_1_101110111010;
      patterns[56792] = 29'b1_101110111011_000_1_101110111011;
      patterns[56793] = 29'b1_101110111011_001_1_111011101110;
      patterns[56794] = 29'b1_101110111011_010_1_011101110111;
      patterns[56795] = 29'b1_101110111011_011_0_111011101111;
      patterns[56796] = 29'b1_101110111011_100_1_110111011101;
      patterns[56797] = 29'b1_101110111011_101_1_111011101110;
      patterns[56798] = 29'b1_101110111011_110_1_101110111011;
      patterns[56799] = 29'b1_101110111011_111_1_101110111011;
      patterns[56800] = 29'b1_101110111100_000_1_101110111100;
      patterns[56801] = 29'b1_101110111100_001_1_111100101110;
      patterns[56802] = 29'b1_101110111100_010_1_011101111001;
      patterns[56803] = 29'b1_101110111100_011_0_111011110011;
      patterns[56804] = 29'b1_101110111100_100_0_110111011110;
      patterns[56805] = 29'b1_101110111100_101_0_011011101111;
      patterns[56806] = 29'b1_101110111100_110_1_101110111100;
      patterns[56807] = 29'b1_101110111100_111_1_101110111100;
      patterns[56808] = 29'b1_101110111101_000_1_101110111101;
      patterns[56809] = 29'b1_101110111101_001_1_111101101110;
      patterns[56810] = 29'b1_101110111101_010_1_011101111011;
      patterns[56811] = 29'b1_101110111101_011_0_111011110111;
      patterns[56812] = 29'b1_101110111101_100_1_110111011110;
      patterns[56813] = 29'b1_101110111101_101_0_111011101111;
      patterns[56814] = 29'b1_101110111101_110_1_101110111101;
      patterns[56815] = 29'b1_101110111101_111_1_101110111101;
      patterns[56816] = 29'b1_101110111110_000_1_101110111110;
      patterns[56817] = 29'b1_101110111110_001_1_111110101110;
      patterns[56818] = 29'b1_101110111110_010_1_011101111101;
      patterns[56819] = 29'b1_101110111110_011_0_111011111011;
      patterns[56820] = 29'b1_101110111110_100_0_110111011111;
      patterns[56821] = 29'b1_101110111110_101_1_011011101111;
      patterns[56822] = 29'b1_101110111110_110_1_101110111110;
      patterns[56823] = 29'b1_101110111110_111_1_101110111110;
      patterns[56824] = 29'b1_101110111111_000_1_101110111111;
      patterns[56825] = 29'b1_101110111111_001_1_111111101110;
      patterns[56826] = 29'b1_101110111111_010_1_011101111111;
      patterns[56827] = 29'b1_101110111111_011_0_111011111111;
      patterns[56828] = 29'b1_101110111111_100_1_110111011111;
      patterns[56829] = 29'b1_101110111111_101_1_111011101111;
      patterns[56830] = 29'b1_101110111111_110_1_101110111111;
      patterns[56831] = 29'b1_101110111111_111_1_101110111111;
      patterns[56832] = 29'b1_101111000000_000_1_101111000000;
      patterns[56833] = 29'b1_101111000000_001_1_000000101111;
      patterns[56834] = 29'b1_101111000000_010_1_011110000001;
      patterns[56835] = 29'b1_101111000000_011_0_111100000011;
      patterns[56836] = 29'b1_101111000000_100_0_110111100000;
      patterns[56837] = 29'b1_101111000000_101_0_011011110000;
      patterns[56838] = 29'b1_101111000000_110_1_101111000000;
      patterns[56839] = 29'b1_101111000000_111_1_101111000000;
      patterns[56840] = 29'b1_101111000001_000_1_101111000001;
      patterns[56841] = 29'b1_101111000001_001_1_000001101111;
      patterns[56842] = 29'b1_101111000001_010_1_011110000011;
      patterns[56843] = 29'b1_101111000001_011_0_111100000111;
      patterns[56844] = 29'b1_101111000001_100_1_110111100000;
      patterns[56845] = 29'b1_101111000001_101_0_111011110000;
      patterns[56846] = 29'b1_101111000001_110_1_101111000001;
      patterns[56847] = 29'b1_101111000001_111_1_101111000001;
      patterns[56848] = 29'b1_101111000010_000_1_101111000010;
      patterns[56849] = 29'b1_101111000010_001_1_000010101111;
      patterns[56850] = 29'b1_101111000010_010_1_011110000101;
      patterns[56851] = 29'b1_101111000010_011_0_111100001011;
      patterns[56852] = 29'b1_101111000010_100_0_110111100001;
      patterns[56853] = 29'b1_101111000010_101_1_011011110000;
      patterns[56854] = 29'b1_101111000010_110_1_101111000010;
      patterns[56855] = 29'b1_101111000010_111_1_101111000010;
      patterns[56856] = 29'b1_101111000011_000_1_101111000011;
      patterns[56857] = 29'b1_101111000011_001_1_000011101111;
      patterns[56858] = 29'b1_101111000011_010_1_011110000111;
      patterns[56859] = 29'b1_101111000011_011_0_111100001111;
      patterns[56860] = 29'b1_101111000011_100_1_110111100001;
      patterns[56861] = 29'b1_101111000011_101_1_111011110000;
      patterns[56862] = 29'b1_101111000011_110_1_101111000011;
      patterns[56863] = 29'b1_101111000011_111_1_101111000011;
      patterns[56864] = 29'b1_101111000100_000_1_101111000100;
      patterns[56865] = 29'b1_101111000100_001_1_000100101111;
      patterns[56866] = 29'b1_101111000100_010_1_011110001001;
      patterns[56867] = 29'b1_101111000100_011_0_111100010011;
      patterns[56868] = 29'b1_101111000100_100_0_110111100010;
      patterns[56869] = 29'b1_101111000100_101_0_011011110001;
      patterns[56870] = 29'b1_101111000100_110_1_101111000100;
      patterns[56871] = 29'b1_101111000100_111_1_101111000100;
      patterns[56872] = 29'b1_101111000101_000_1_101111000101;
      patterns[56873] = 29'b1_101111000101_001_1_000101101111;
      patterns[56874] = 29'b1_101111000101_010_1_011110001011;
      patterns[56875] = 29'b1_101111000101_011_0_111100010111;
      patterns[56876] = 29'b1_101111000101_100_1_110111100010;
      patterns[56877] = 29'b1_101111000101_101_0_111011110001;
      patterns[56878] = 29'b1_101111000101_110_1_101111000101;
      patterns[56879] = 29'b1_101111000101_111_1_101111000101;
      patterns[56880] = 29'b1_101111000110_000_1_101111000110;
      patterns[56881] = 29'b1_101111000110_001_1_000110101111;
      patterns[56882] = 29'b1_101111000110_010_1_011110001101;
      patterns[56883] = 29'b1_101111000110_011_0_111100011011;
      patterns[56884] = 29'b1_101111000110_100_0_110111100011;
      patterns[56885] = 29'b1_101111000110_101_1_011011110001;
      patterns[56886] = 29'b1_101111000110_110_1_101111000110;
      patterns[56887] = 29'b1_101111000110_111_1_101111000110;
      patterns[56888] = 29'b1_101111000111_000_1_101111000111;
      patterns[56889] = 29'b1_101111000111_001_1_000111101111;
      patterns[56890] = 29'b1_101111000111_010_1_011110001111;
      patterns[56891] = 29'b1_101111000111_011_0_111100011111;
      patterns[56892] = 29'b1_101111000111_100_1_110111100011;
      patterns[56893] = 29'b1_101111000111_101_1_111011110001;
      patterns[56894] = 29'b1_101111000111_110_1_101111000111;
      patterns[56895] = 29'b1_101111000111_111_1_101111000111;
      patterns[56896] = 29'b1_101111001000_000_1_101111001000;
      patterns[56897] = 29'b1_101111001000_001_1_001000101111;
      patterns[56898] = 29'b1_101111001000_010_1_011110010001;
      patterns[56899] = 29'b1_101111001000_011_0_111100100011;
      patterns[56900] = 29'b1_101111001000_100_0_110111100100;
      patterns[56901] = 29'b1_101111001000_101_0_011011110010;
      patterns[56902] = 29'b1_101111001000_110_1_101111001000;
      patterns[56903] = 29'b1_101111001000_111_1_101111001000;
      patterns[56904] = 29'b1_101111001001_000_1_101111001001;
      patterns[56905] = 29'b1_101111001001_001_1_001001101111;
      patterns[56906] = 29'b1_101111001001_010_1_011110010011;
      patterns[56907] = 29'b1_101111001001_011_0_111100100111;
      patterns[56908] = 29'b1_101111001001_100_1_110111100100;
      patterns[56909] = 29'b1_101111001001_101_0_111011110010;
      patterns[56910] = 29'b1_101111001001_110_1_101111001001;
      patterns[56911] = 29'b1_101111001001_111_1_101111001001;
      patterns[56912] = 29'b1_101111001010_000_1_101111001010;
      patterns[56913] = 29'b1_101111001010_001_1_001010101111;
      patterns[56914] = 29'b1_101111001010_010_1_011110010101;
      patterns[56915] = 29'b1_101111001010_011_0_111100101011;
      patterns[56916] = 29'b1_101111001010_100_0_110111100101;
      patterns[56917] = 29'b1_101111001010_101_1_011011110010;
      patterns[56918] = 29'b1_101111001010_110_1_101111001010;
      patterns[56919] = 29'b1_101111001010_111_1_101111001010;
      patterns[56920] = 29'b1_101111001011_000_1_101111001011;
      patterns[56921] = 29'b1_101111001011_001_1_001011101111;
      patterns[56922] = 29'b1_101111001011_010_1_011110010111;
      patterns[56923] = 29'b1_101111001011_011_0_111100101111;
      patterns[56924] = 29'b1_101111001011_100_1_110111100101;
      patterns[56925] = 29'b1_101111001011_101_1_111011110010;
      patterns[56926] = 29'b1_101111001011_110_1_101111001011;
      patterns[56927] = 29'b1_101111001011_111_1_101111001011;
      patterns[56928] = 29'b1_101111001100_000_1_101111001100;
      patterns[56929] = 29'b1_101111001100_001_1_001100101111;
      patterns[56930] = 29'b1_101111001100_010_1_011110011001;
      patterns[56931] = 29'b1_101111001100_011_0_111100110011;
      patterns[56932] = 29'b1_101111001100_100_0_110111100110;
      patterns[56933] = 29'b1_101111001100_101_0_011011110011;
      patterns[56934] = 29'b1_101111001100_110_1_101111001100;
      patterns[56935] = 29'b1_101111001100_111_1_101111001100;
      patterns[56936] = 29'b1_101111001101_000_1_101111001101;
      patterns[56937] = 29'b1_101111001101_001_1_001101101111;
      patterns[56938] = 29'b1_101111001101_010_1_011110011011;
      patterns[56939] = 29'b1_101111001101_011_0_111100110111;
      patterns[56940] = 29'b1_101111001101_100_1_110111100110;
      patterns[56941] = 29'b1_101111001101_101_0_111011110011;
      patterns[56942] = 29'b1_101111001101_110_1_101111001101;
      patterns[56943] = 29'b1_101111001101_111_1_101111001101;
      patterns[56944] = 29'b1_101111001110_000_1_101111001110;
      patterns[56945] = 29'b1_101111001110_001_1_001110101111;
      patterns[56946] = 29'b1_101111001110_010_1_011110011101;
      patterns[56947] = 29'b1_101111001110_011_0_111100111011;
      patterns[56948] = 29'b1_101111001110_100_0_110111100111;
      patterns[56949] = 29'b1_101111001110_101_1_011011110011;
      patterns[56950] = 29'b1_101111001110_110_1_101111001110;
      patterns[56951] = 29'b1_101111001110_111_1_101111001110;
      patterns[56952] = 29'b1_101111001111_000_1_101111001111;
      patterns[56953] = 29'b1_101111001111_001_1_001111101111;
      patterns[56954] = 29'b1_101111001111_010_1_011110011111;
      patterns[56955] = 29'b1_101111001111_011_0_111100111111;
      patterns[56956] = 29'b1_101111001111_100_1_110111100111;
      patterns[56957] = 29'b1_101111001111_101_1_111011110011;
      patterns[56958] = 29'b1_101111001111_110_1_101111001111;
      patterns[56959] = 29'b1_101111001111_111_1_101111001111;
      patterns[56960] = 29'b1_101111010000_000_1_101111010000;
      patterns[56961] = 29'b1_101111010000_001_1_010000101111;
      patterns[56962] = 29'b1_101111010000_010_1_011110100001;
      patterns[56963] = 29'b1_101111010000_011_0_111101000011;
      patterns[56964] = 29'b1_101111010000_100_0_110111101000;
      patterns[56965] = 29'b1_101111010000_101_0_011011110100;
      patterns[56966] = 29'b1_101111010000_110_1_101111010000;
      patterns[56967] = 29'b1_101111010000_111_1_101111010000;
      patterns[56968] = 29'b1_101111010001_000_1_101111010001;
      patterns[56969] = 29'b1_101111010001_001_1_010001101111;
      patterns[56970] = 29'b1_101111010001_010_1_011110100011;
      patterns[56971] = 29'b1_101111010001_011_0_111101000111;
      patterns[56972] = 29'b1_101111010001_100_1_110111101000;
      patterns[56973] = 29'b1_101111010001_101_0_111011110100;
      patterns[56974] = 29'b1_101111010001_110_1_101111010001;
      patterns[56975] = 29'b1_101111010001_111_1_101111010001;
      patterns[56976] = 29'b1_101111010010_000_1_101111010010;
      patterns[56977] = 29'b1_101111010010_001_1_010010101111;
      patterns[56978] = 29'b1_101111010010_010_1_011110100101;
      patterns[56979] = 29'b1_101111010010_011_0_111101001011;
      patterns[56980] = 29'b1_101111010010_100_0_110111101001;
      patterns[56981] = 29'b1_101111010010_101_1_011011110100;
      patterns[56982] = 29'b1_101111010010_110_1_101111010010;
      patterns[56983] = 29'b1_101111010010_111_1_101111010010;
      patterns[56984] = 29'b1_101111010011_000_1_101111010011;
      patterns[56985] = 29'b1_101111010011_001_1_010011101111;
      patterns[56986] = 29'b1_101111010011_010_1_011110100111;
      patterns[56987] = 29'b1_101111010011_011_0_111101001111;
      patterns[56988] = 29'b1_101111010011_100_1_110111101001;
      patterns[56989] = 29'b1_101111010011_101_1_111011110100;
      patterns[56990] = 29'b1_101111010011_110_1_101111010011;
      patterns[56991] = 29'b1_101111010011_111_1_101111010011;
      patterns[56992] = 29'b1_101111010100_000_1_101111010100;
      patterns[56993] = 29'b1_101111010100_001_1_010100101111;
      patterns[56994] = 29'b1_101111010100_010_1_011110101001;
      patterns[56995] = 29'b1_101111010100_011_0_111101010011;
      patterns[56996] = 29'b1_101111010100_100_0_110111101010;
      patterns[56997] = 29'b1_101111010100_101_0_011011110101;
      patterns[56998] = 29'b1_101111010100_110_1_101111010100;
      patterns[56999] = 29'b1_101111010100_111_1_101111010100;
      patterns[57000] = 29'b1_101111010101_000_1_101111010101;
      patterns[57001] = 29'b1_101111010101_001_1_010101101111;
      patterns[57002] = 29'b1_101111010101_010_1_011110101011;
      patterns[57003] = 29'b1_101111010101_011_0_111101010111;
      patterns[57004] = 29'b1_101111010101_100_1_110111101010;
      patterns[57005] = 29'b1_101111010101_101_0_111011110101;
      patterns[57006] = 29'b1_101111010101_110_1_101111010101;
      patterns[57007] = 29'b1_101111010101_111_1_101111010101;
      patterns[57008] = 29'b1_101111010110_000_1_101111010110;
      patterns[57009] = 29'b1_101111010110_001_1_010110101111;
      patterns[57010] = 29'b1_101111010110_010_1_011110101101;
      patterns[57011] = 29'b1_101111010110_011_0_111101011011;
      patterns[57012] = 29'b1_101111010110_100_0_110111101011;
      patterns[57013] = 29'b1_101111010110_101_1_011011110101;
      patterns[57014] = 29'b1_101111010110_110_1_101111010110;
      patterns[57015] = 29'b1_101111010110_111_1_101111010110;
      patterns[57016] = 29'b1_101111010111_000_1_101111010111;
      patterns[57017] = 29'b1_101111010111_001_1_010111101111;
      patterns[57018] = 29'b1_101111010111_010_1_011110101111;
      patterns[57019] = 29'b1_101111010111_011_0_111101011111;
      patterns[57020] = 29'b1_101111010111_100_1_110111101011;
      patterns[57021] = 29'b1_101111010111_101_1_111011110101;
      patterns[57022] = 29'b1_101111010111_110_1_101111010111;
      patterns[57023] = 29'b1_101111010111_111_1_101111010111;
      patterns[57024] = 29'b1_101111011000_000_1_101111011000;
      patterns[57025] = 29'b1_101111011000_001_1_011000101111;
      patterns[57026] = 29'b1_101111011000_010_1_011110110001;
      patterns[57027] = 29'b1_101111011000_011_0_111101100011;
      patterns[57028] = 29'b1_101111011000_100_0_110111101100;
      patterns[57029] = 29'b1_101111011000_101_0_011011110110;
      patterns[57030] = 29'b1_101111011000_110_1_101111011000;
      patterns[57031] = 29'b1_101111011000_111_1_101111011000;
      patterns[57032] = 29'b1_101111011001_000_1_101111011001;
      patterns[57033] = 29'b1_101111011001_001_1_011001101111;
      patterns[57034] = 29'b1_101111011001_010_1_011110110011;
      patterns[57035] = 29'b1_101111011001_011_0_111101100111;
      patterns[57036] = 29'b1_101111011001_100_1_110111101100;
      patterns[57037] = 29'b1_101111011001_101_0_111011110110;
      patterns[57038] = 29'b1_101111011001_110_1_101111011001;
      patterns[57039] = 29'b1_101111011001_111_1_101111011001;
      patterns[57040] = 29'b1_101111011010_000_1_101111011010;
      patterns[57041] = 29'b1_101111011010_001_1_011010101111;
      patterns[57042] = 29'b1_101111011010_010_1_011110110101;
      patterns[57043] = 29'b1_101111011010_011_0_111101101011;
      patterns[57044] = 29'b1_101111011010_100_0_110111101101;
      patterns[57045] = 29'b1_101111011010_101_1_011011110110;
      patterns[57046] = 29'b1_101111011010_110_1_101111011010;
      patterns[57047] = 29'b1_101111011010_111_1_101111011010;
      patterns[57048] = 29'b1_101111011011_000_1_101111011011;
      patterns[57049] = 29'b1_101111011011_001_1_011011101111;
      patterns[57050] = 29'b1_101111011011_010_1_011110110111;
      patterns[57051] = 29'b1_101111011011_011_0_111101101111;
      patterns[57052] = 29'b1_101111011011_100_1_110111101101;
      patterns[57053] = 29'b1_101111011011_101_1_111011110110;
      patterns[57054] = 29'b1_101111011011_110_1_101111011011;
      patterns[57055] = 29'b1_101111011011_111_1_101111011011;
      patterns[57056] = 29'b1_101111011100_000_1_101111011100;
      patterns[57057] = 29'b1_101111011100_001_1_011100101111;
      patterns[57058] = 29'b1_101111011100_010_1_011110111001;
      patterns[57059] = 29'b1_101111011100_011_0_111101110011;
      patterns[57060] = 29'b1_101111011100_100_0_110111101110;
      patterns[57061] = 29'b1_101111011100_101_0_011011110111;
      patterns[57062] = 29'b1_101111011100_110_1_101111011100;
      patterns[57063] = 29'b1_101111011100_111_1_101111011100;
      patterns[57064] = 29'b1_101111011101_000_1_101111011101;
      patterns[57065] = 29'b1_101111011101_001_1_011101101111;
      patterns[57066] = 29'b1_101111011101_010_1_011110111011;
      patterns[57067] = 29'b1_101111011101_011_0_111101110111;
      patterns[57068] = 29'b1_101111011101_100_1_110111101110;
      patterns[57069] = 29'b1_101111011101_101_0_111011110111;
      patterns[57070] = 29'b1_101111011101_110_1_101111011101;
      patterns[57071] = 29'b1_101111011101_111_1_101111011101;
      patterns[57072] = 29'b1_101111011110_000_1_101111011110;
      patterns[57073] = 29'b1_101111011110_001_1_011110101111;
      patterns[57074] = 29'b1_101111011110_010_1_011110111101;
      patterns[57075] = 29'b1_101111011110_011_0_111101111011;
      patterns[57076] = 29'b1_101111011110_100_0_110111101111;
      patterns[57077] = 29'b1_101111011110_101_1_011011110111;
      patterns[57078] = 29'b1_101111011110_110_1_101111011110;
      patterns[57079] = 29'b1_101111011110_111_1_101111011110;
      patterns[57080] = 29'b1_101111011111_000_1_101111011111;
      patterns[57081] = 29'b1_101111011111_001_1_011111101111;
      patterns[57082] = 29'b1_101111011111_010_1_011110111111;
      patterns[57083] = 29'b1_101111011111_011_0_111101111111;
      patterns[57084] = 29'b1_101111011111_100_1_110111101111;
      patterns[57085] = 29'b1_101111011111_101_1_111011110111;
      patterns[57086] = 29'b1_101111011111_110_1_101111011111;
      patterns[57087] = 29'b1_101111011111_111_1_101111011111;
      patterns[57088] = 29'b1_101111100000_000_1_101111100000;
      patterns[57089] = 29'b1_101111100000_001_1_100000101111;
      patterns[57090] = 29'b1_101111100000_010_1_011111000001;
      patterns[57091] = 29'b1_101111100000_011_0_111110000011;
      patterns[57092] = 29'b1_101111100000_100_0_110111110000;
      patterns[57093] = 29'b1_101111100000_101_0_011011111000;
      patterns[57094] = 29'b1_101111100000_110_1_101111100000;
      patterns[57095] = 29'b1_101111100000_111_1_101111100000;
      patterns[57096] = 29'b1_101111100001_000_1_101111100001;
      patterns[57097] = 29'b1_101111100001_001_1_100001101111;
      patterns[57098] = 29'b1_101111100001_010_1_011111000011;
      patterns[57099] = 29'b1_101111100001_011_0_111110000111;
      patterns[57100] = 29'b1_101111100001_100_1_110111110000;
      patterns[57101] = 29'b1_101111100001_101_0_111011111000;
      patterns[57102] = 29'b1_101111100001_110_1_101111100001;
      patterns[57103] = 29'b1_101111100001_111_1_101111100001;
      patterns[57104] = 29'b1_101111100010_000_1_101111100010;
      patterns[57105] = 29'b1_101111100010_001_1_100010101111;
      patterns[57106] = 29'b1_101111100010_010_1_011111000101;
      patterns[57107] = 29'b1_101111100010_011_0_111110001011;
      patterns[57108] = 29'b1_101111100010_100_0_110111110001;
      patterns[57109] = 29'b1_101111100010_101_1_011011111000;
      patterns[57110] = 29'b1_101111100010_110_1_101111100010;
      patterns[57111] = 29'b1_101111100010_111_1_101111100010;
      patterns[57112] = 29'b1_101111100011_000_1_101111100011;
      patterns[57113] = 29'b1_101111100011_001_1_100011101111;
      patterns[57114] = 29'b1_101111100011_010_1_011111000111;
      patterns[57115] = 29'b1_101111100011_011_0_111110001111;
      patterns[57116] = 29'b1_101111100011_100_1_110111110001;
      patterns[57117] = 29'b1_101111100011_101_1_111011111000;
      patterns[57118] = 29'b1_101111100011_110_1_101111100011;
      patterns[57119] = 29'b1_101111100011_111_1_101111100011;
      patterns[57120] = 29'b1_101111100100_000_1_101111100100;
      patterns[57121] = 29'b1_101111100100_001_1_100100101111;
      patterns[57122] = 29'b1_101111100100_010_1_011111001001;
      patterns[57123] = 29'b1_101111100100_011_0_111110010011;
      patterns[57124] = 29'b1_101111100100_100_0_110111110010;
      patterns[57125] = 29'b1_101111100100_101_0_011011111001;
      patterns[57126] = 29'b1_101111100100_110_1_101111100100;
      patterns[57127] = 29'b1_101111100100_111_1_101111100100;
      patterns[57128] = 29'b1_101111100101_000_1_101111100101;
      patterns[57129] = 29'b1_101111100101_001_1_100101101111;
      patterns[57130] = 29'b1_101111100101_010_1_011111001011;
      patterns[57131] = 29'b1_101111100101_011_0_111110010111;
      patterns[57132] = 29'b1_101111100101_100_1_110111110010;
      patterns[57133] = 29'b1_101111100101_101_0_111011111001;
      patterns[57134] = 29'b1_101111100101_110_1_101111100101;
      patterns[57135] = 29'b1_101111100101_111_1_101111100101;
      patterns[57136] = 29'b1_101111100110_000_1_101111100110;
      patterns[57137] = 29'b1_101111100110_001_1_100110101111;
      patterns[57138] = 29'b1_101111100110_010_1_011111001101;
      patterns[57139] = 29'b1_101111100110_011_0_111110011011;
      patterns[57140] = 29'b1_101111100110_100_0_110111110011;
      patterns[57141] = 29'b1_101111100110_101_1_011011111001;
      patterns[57142] = 29'b1_101111100110_110_1_101111100110;
      patterns[57143] = 29'b1_101111100110_111_1_101111100110;
      patterns[57144] = 29'b1_101111100111_000_1_101111100111;
      patterns[57145] = 29'b1_101111100111_001_1_100111101111;
      patterns[57146] = 29'b1_101111100111_010_1_011111001111;
      patterns[57147] = 29'b1_101111100111_011_0_111110011111;
      patterns[57148] = 29'b1_101111100111_100_1_110111110011;
      patterns[57149] = 29'b1_101111100111_101_1_111011111001;
      patterns[57150] = 29'b1_101111100111_110_1_101111100111;
      patterns[57151] = 29'b1_101111100111_111_1_101111100111;
      patterns[57152] = 29'b1_101111101000_000_1_101111101000;
      patterns[57153] = 29'b1_101111101000_001_1_101000101111;
      patterns[57154] = 29'b1_101111101000_010_1_011111010001;
      patterns[57155] = 29'b1_101111101000_011_0_111110100011;
      patterns[57156] = 29'b1_101111101000_100_0_110111110100;
      patterns[57157] = 29'b1_101111101000_101_0_011011111010;
      patterns[57158] = 29'b1_101111101000_110_1_101111101000;
      patterns[57159] = 29'b1_101111101000_111_1_101111101000;
      patterns[57160] = 29'b1_101111101001_000_1_101111101001;
      patterns[57161] = 29'b1_101111101001_001_1_101001101111;
      patterns[57162] = 29'b1_101111101001_010_1_011111010011;
      patterns[57163] = 29'b1_101111101001_011_0_111110100111;
      patterns[57164] = 29'b1_101111101001_100_1_110111110100;
      patterns[57165] = 29'b1_101111101001_101_0_111011111010;
      patterns[57166] = 29'b1_101111101001_110_1_101111101001;
      patterns[57167] = 29'b1_101111101001_111_1_101111101001;
      patterns[57168] = 29'b1_101111101010_000_1_101111101010;
      patterns[57169] = 29'b1_101111101010_001_1_101010101111;
      patterns[57170] = 29'b1_101111101010_010_1_011111010101;
      patterns[57171] = 29'b1_101111101010_011_0_111110101011;
      patterns[57172] = 29'b1_101111101010_100_0_110111110101;
      patterns[57173] = 29'b1_101111101010_101_1_011011111010;
      patterns[57174] = 29'b1_101111101010_110_1_101111101010;
      patterns[57175] = 29'b1_101111101010_111_1_101111101010;
      patterns[57176] = 29'b1_101111101011_000_1_101111101011;
      patterns[57177] = 29'b1_101111101011_001_1_101011101111;
      patterns[57178] = 29'b1_101111101011_010_1_011111010111;
      patterns[57179] = 29'b1_101111101011_011_0_111110101111;
      patterns[57180] = 29'b1_101111101011_100_1_110111110101;
      patterns[57181] = 29'b1_101111101011_101_1_111011111010;
      patterns[57182] = 29'b1_101111101011_110_1_101111101011;
      patterns[57183] = 29'b1_101111101011_111_1_101111101011;
      patterns[57184] = 29'b1_101111101100_000_1_101111101100;
      patterns[57185] = 29'b1_101111101100_001_1_101100101111;
      patterns[57186] = 29'b1_101111101100_010_1_011111011001;
      patterns[57187] = 29'b1_101111101100_011_0_111110110011;
      patterns[57188] = 29'b1_101111101100_100_0_110111110110;
      patterns[57189] = 29'b1_101111101100_101_0_011011111011;
      patterns[57190] = 29'b1_101111101100_110_1_101111101100;
      patterns[57191] = 29'b1_101111101100_111_1_101111101100;
      patterns[57192] = 29'b1_101111101101_000_1_101111101101;
      patterns[57193] = 29'b1_101111101101_001_1_101101101111;
      patterns[57194] = 29'b1_101111101101_010_1_011111011011;
      patterns[57195] = 29'b1_101111101101_011_0_111110110111;
      patterns[57196] = 29'b1_101111101101_100_1_110111110110;
      patterns[57197] = 29'b1_101111101101_101_0_111011111011;
      patterns[57198] = 29'b1_101111101101_110_1_101111101101;
      patterns[57199] = 29'b1_101111101101_111_1_101111101101;
      patterns[57200] = 29'b1_101111101110_000_1_101111101110;
      patterns[57201] = 29'b1_101111101110_001_1_101110101111;
      patterns[57202] = 29'b1_101111101110_010_1_011111011101;
      patterns[57203] = 29'b1_101111101110_011_0_111110111011;
      patterns[57204] = 29'b1_101111101110_100_0_110111110111;
      patterns[57205] = 29'b1_101111101110_101_1_011011111011;
      patterns[57206] = 29'b1_101111101110_110_1_101111101110;
      patterns[57207] = 29'b1_101111101110_111_1_101111101110;
      patterns[57208] = 29'b1_101111101111_000_1_101111101111;
      patterns[57209] = 29'b1_101111101111_001_1_101111101111;
      patterns[57210] = 29'b1_101111101111_010_1_011111011111;
      patterns[57211] = 29'b1_101111101111_011_0_111110111111;
      patterns[57212] = 29'b1_101111101111_100_1_110111110111;
      patterns[57213] = 29'b1_101111101111_101_1_111011111011;
      patterns[57214] = 29'b1_101111101111_110_1_101111101111;
      patterns[57215] = 29'b1_101111101111_111_1_101111101111;
      patterns[57216] = 29'b1_101111110000_000_1_101111110000;
      patterns[57217] = 29'b1_101111110000_001_1_110000101111;
      patterns[57218] = 29'b1_101111110000_010_1_011111100001;
      patterns[57219] = 29'b1_101111110000_011_0_111111000011;
      patterns[57220] = 29'b1_101111110000_100_0_110111111000;
      patterns[57221] = 29'b1_101111110000_101_0_011011111100;
      patterns[57222] = 29'b1_101111110000_110_1_101111110000;
      patterns[57223] = 29'b1_101111110000_111_1_101111110000;
      patterns[57224] = 29'b1_101111110001_000_1_101111110001;
      patterns[57225] = 29'b1_101111110001_001_1_110001101111;
      patterns[57226] = 29'b1_101111110001_010_1_011111100011;
      patterns[57227] = 29'b1_101111110001_011_0_111111000111;
      patterns[57228] = 29'b1_101111110001_100_1_110111111000;
      patterns[57229] = 29'b1_101111110001_101_0_111011111100;
      patterns[57230] = 29'b1_101111110001_110_1_101111110001;
      patterns[57231] = 29'b1_101111110001_111_1_101111110001;
      patterns[57232] = 29'b1_101111110010_000_1_101111110010;
      patterns[57233] = 29'b1_101111110010_001_1_110010101111;
      patterns[57234] = 29'b1_101111110010_010_1_011111100101;
      patterns[57235] = 29'b1_101111110010_011_0_111111001011;
      patterns[57236] = 29'b1_101111110010_100_0_110111111001;
      patterns[57237] = 29'b1_101111110010_101_1_011011111100;
      patterns[57238] = 29'b1_101111110010_110_1_101111110010;
      patterns[57239] = 29'b1_101111110010_111_1_101111110010;
      patterns[57240] = 29'b1_101111110011_000_1_101111110011;
      patterns[57241] = 29'b1_101111110011_001_1_110011101111;
      patterns[57242] = 29'b1_101111110011_010_1_011111100111;
      patterns[57243] = 29'b1_101111110011_011_0_111111001111;
      patterns[57244] = 29'b1_101111110011_100_1_110111111001;
      patterns[57245] = 29'b1_101111110011_101_1_111011111100;
      patterns[57246] = 29'b1_101111110011_110_1_101111110011;
      patterns[57247] = 29'b1_101111110011_111_1_101111110011;
      patterns[57248] = 29'b1_101111110100_000_1_101111110100;
      patterns[57249] = 29'b1_101111110100_001_1_110100101111;
      patterns[57250] = 29'b1_101111110100_010_1_011111101001;
      patterns[57251] = 29'b1_101111110100_011_0_111111010011;
      patterns[57252] = 29'b1_101111110100_100_0_110111111010;
      patterns[57253] = 29'b1_101111110100_101_0_011011111101;
      patterns[57254] = 29'b1_101111110100_110_1_101111110100;
      patterns[57255] = 29'b1_101111110100_111_1_101111110100;
      patterns[57256] = 29'b1_101111110101_000_1_101111110101;
      patterns[57257] = 29'b1_101111110101_001_1_110101101111;
      patterns[57258] = 29'b1_101111110101_010_1_011111101011;
      patterns[57259] = 29'b1_101111110101_011_0_111111010111;
      patterns[57260] = 29'b1_101111110101_100_1_110111111010;
      patterns[57261] = 29'b1_101111110101_101_0_111011111101;
      patterns[57262] = 29'b1_101111110101_110_1_101111110101;
      patterns[57263] = 29'b1_101111110101_111_1_101111110101;
      patterns[57264] = 29'b1_101111110110_000_1_101111110110;
      patterns[57265] = 29'b1_101111110110_001_1_110110101111;
      patterns[57266] = 29'b1_101111110110_010_1_011111101101;
      patterns[57267] = 29'b1_101111110110_011_0_111111011011;
      patterns[57268] = 29'b1_101111110110_100_0_110111111011;
      patterns[57269] = 29'b1_101111110110_101_1_011011111101;
      patterns[57270] = 29'b1_101111110110_110_1_101111110110;
      patterns[57271] = 29'b1_101111110110_111_1_101111110110;
      patterns[57272] = 29'b1_101111110111_000_1_101111110111;
      patterns[57273] = 29'b1_101111110111_001_1_110111101111;
      patterns[57274] = 29'b1_101111110111_010_1_011111101111;
      patterns[57275] = 29'b1_101111110111_011_0_111111011111;
      patterns[57276] = 29'b1_101111110111_100_1_110111111011;
      patterns[57277] = 29'b1_101111110111_101_1_111011111101;
      patterns[57278] = 29'b1_101111110111_110_1_101111110111;
      patterns[57279] = 29'b1_101111110111_111_1_101111110111;
      patterns[57280] = 29'b1_101111111000_000_1_101111111000;
      patterns[57281] = 29'b1_101111111000_001_1_111000101111;
      patterns[57282] = 29'b1_101111111000_010_1_011111110001;
      patterns[57283] = 29'b1_101111111000_011_0_111111100011;
      patterns[57284] = 29'b1_101111111000_100_0_110111111100;
      patterns[57285] = 29'b1_101111111000_101_0_011011111110;
      patterns[57286] = 29'b1_101111111000_110_1_101111111000;
      patterns[57287] = 29'b1_101111111000_111_1_101111111000;
      patterns[57288] = 29'b1_101111111001_000_1_101111111001;
      patterns[57289] = 29'b1_101111111001_001_1_111001101111;
      patterns[57290] = 29'b1_101111111001_010_1_011111110011;
      patterns[57291] = 29'b1_101111111001_011_0_111111100111;
      patterns[57292] = 29'b1_101111111001_100_1_110111111100;
      patterns[57293] = 29'b1_101111111001_101_0_111011111110;
      patterns[57294] = 29'b1_101111111001_110_1_101111111001;
      patterns[57295] = 29'b1_101111111001_111_1_101111111001;
      patterns[57296] = 29'b1_101111111010_000_1_101111111010;
      patterns[57297] = 29'b1_101111111010_001_1_111010101111;
      patterns[57298] = 29'b1_101111111010_010_1_011111110101;
      patterns[57299] = 29'b1_101111111010_011_0_111111101011;
      patterns[57300] = 29'b1_101111111010_100_0_110111111101;
      patterns[57301] = 29'b1_101111111010_101_1_011011111110;
      patterns[57302] = 29'b1_101111111010_110_1_101111111010;
      patterns[57303] = 29'b1_101111111010_111_1_101111111010;
      patterns[57304] = 29'b1_101111111011_000_1_101111111011;
      patterns[57305] = 29'b1_101111111011_001_1_111011101111;
      patterns[57306] = 29'b1_101111111011_010_1_011111110111;
      patterns[57307] = 29'b1_101111111011_011_0_111111101111;
      patterns[57308] = 29'b1_101111111011_100_1_110111111101;
      patterns[57309] = 29'b1_101111111011_101_1_111011111110;
      patterns[57310] = 29'b1_101111111011_110_1_101111111011;
      patterns[57311] = 29'b1_101111111011_111_1_101111111011;
      patterns[57312] = 29'b1_101111111100_000_1_101111111100;
      patterns[57313] = 29'b1_101111111100_001_1_111100101111;
      patterns[57314] = 29'b1_101111111100_010_1_011111111001;
      patterns[57315] = 29'b1_101111111100_011_0_111111110011;
      patterns[57316] = 29'b1_101111111100_100_0_110111111110;
      patterns[57317] = 29'b1_101111111100_101_0_011011111111;
      patterns[57318] = 29'b1_101111111100_110_1_101111111100;
      patterns[57319] = 29'b1_101111111100_111_1_101111111100;
      patterns[57320] = 29'b1_101111111101_000_1_101111111101;
      patterns[57321] = 29'b1_101111111101_001_1_111101101111;
      patterns[57322] = 29'b1_101111111101_010_1_011111111011;
      patterns[57323] = 29'b1_101111111101_011_0_111111110111;
      patterns[57324] = 29'b1_101111111101_100_1_110111111110;
      patterns[57325] = 29'b1_101111111101_101_0_111011111111;
      patterns[57326] = 29'b1_101111111101_110_1_101111111101;
      patterns[57327] = 29'b1_101111111101_111_1_101111111101;
      patterns[57328] = 29'b1_101111111110_000_1_101111111110;
      patterns[57329] = 29'b1_101111111110_001_1_111110101111;
      patterns[57330] = 29'b1_101111111110_010_1_011111111101;
      patterns[57331] = 29'b1_101111111110_011_0_111111111011;
      patterns[57332] = 29'b1_101111111110_100_0_110111111111;
      patterns[57333] = 29'b1_101111111110_101_1_011011111111;
      patterns[57334] = 29'b1_101111111110_110_1_101111111110;
      patterns[57335] = 29'b1_101111111110_111_1_101111111110;
      patterns[57336] = 29'b1_101111111111_000_1_101111111111;
      patterns[57337] = 29'b1_101111111111_001_1_111111101111;
      patterns[57338] = 29'b1_101111111111_010_1_011111111111;
      patterns[57339] = 29'b1_101111111111_011_0_111111111111;
      patterns[57340] = 29'b1_101111111111_100_1_110111111111;
      patterns[57341] = 29'b1_101111111111_101_1_111011111111;
      patterns[57342] = 29'b1_101111111111_110_1_101111111111;
      patterns[57343] = 29'b1_101111111111_111_1_101111111111;
      patterns[57344] = 29'b1_110000000000_000_1_110000000000;
      patterns[57345] = 29'b1_110000000000_001_1_000000110000;
      patterns[57346] = 29'b1_110000000000_010_1_100000000001;
      patterns[57347] = 29'b1_110000000000_011_1_000000000011;
      patterns[57348] = 29'b1_110000000000_100_0_111000000000;
      patterns[57349] = 29'b1_110000000000_101_0_011100000000;
      patterns[57350] = 29'b1_110000000000_110_1_110000000000;
      patterns[57351] = 29'b1_110000000000_111_1_110000000000;
      patterns[57352] = 29'b1_110000000001_000_1_110000000001;
      patterns[57353] = 29'b1_110000000001_001_1_000001110000;
      patterns[57354] = 29'b1_110000000001_010_1_100000000011;
      patterns[57355] = 29'b1_110000000001_011_1_000000000111;
      patterns[57356] = 29'b1_110000000001_100_1_111000000000;
      patterns[57357] = 29'b1_110000000001_101_0_111100000000;
      patterns[57358] = 29'b1_110000000001_110_1_110000000001;
      patterns[57359] = 29'b1_110000000001_111_1_110000000001;
      patterns[57360] = 29'b1_110000000010_000_1_110000000010;
      patterns[57361] = 29'b1_110000000010_001_1_000010110000;
      patterns[57362] = 29'b1_110000000010_010_1_100000000101;
      patterns[57363] = 29'b1_110000000010_011_1_000000001011;
      patterns[57364] = 29'b1_110000000010_100_0_111000000001;
      patterns[57365] = 29'b1_110000000010_101_1_011100000000;
      patterns[57366] = 29'b1_110000000010_110_1_110000000010;
      patterns[57367] = 29'b1_110000000010_111_1_110000000010;
      patterns[57368] = 29'b1_110000000011_000_1_110000000011;
      patterns[57369] = 29'b1_110000000011_001_1_000011110000;
      patterns[57370] = 29'b1_110000000011_010_1_100000000111;
      patterns[57371] = 29'b1_110000000011_011_1_000000001111;
      patterns[57372] = 29'b1_110000000011_100_1_111000000001;
      patterns[57373] = 29'b1_110000000011_101_1_111100000000;
      patterns[57374] = 29'b1_110000000011_110_1_110000000011;
      patterns[57375] = 29'b1_110000000011_111_1_110000000011;
      patterns[57376] = 29'b1_110000000100_000_1_110000000100;
      patterns[57377] = 29'b1_110000000100_001_1_000100110000;
      patterns[57378] = 29'b1_110000000100_010_1_100000001001;
      patterns[57379] = 29'b1_110000000100_011_1_000000010011;
      patterns[57380] = 29'b1_110000000100_100_0_111000000010;
      patterns[57381] = 29'b1_110000000100_101_0_011100000001;
      patterns[57382] = 29'b1_110000000100_110_1_110000000100;
      patterns[57383] = 29'b1_110000000100_111_1_110000000100;
      patterns[57384] = 29'b1_110000000101_000_1_110000000101;
      patterns[57385] = 29'b1_110000000101_001_1_000101110000;
      patterns[57386] = 29'b1_110000000101_010_1_100000001011;
      patterns[57387] = 29'b1_110000000101_011_1_000000010111;
      patterns[57388] = 29'b1_110000000101_100_1_111000000010;
      patterns[57389] = 29'b1_110000000101_101_0_111100000001;
      patterns[57390] = 29'b1_110000000101_110_1_110000000101;
      patterns[57391] = 29'b1_110000000101_111_1_110000000101;
      patterns[57392] = 29'b1_110000000110_000_1_110000000110;
      patterns[57393] = 29'b1_110000000110_001_1_000110110000;
      patterns[57394] = 29'b1_110000000110_010_1_100000001101;
      patterns[57395] = 29'b1_110000000110_011_1_000000011011;
      patterns[57396] = 29'b1_110000000110_100_0_111000000011;
      patterns[57397] = 29'b1_110000000110_101_1_011100000001;
      patterns[57398] = 29'b1_110000000110_110_1_110000000110;
      patterns[57399] = 29'b1_110000000110_111_1_110000000110;
      patterns[57400] = 29'b1_110000000111_000_1_110000000111;
      patterns[57401] = 29'b1_110000000111_001_1_000111110000;
      patterns[57402] = 29'b1_110000000111_010_1_100000001111;
      patterns[57403] = 29'b1_110000000111_011_1_000000011111;
      patterns[57404] = 29'b1_110000000111_100_1_111000000011;
      patterns[57405] = 29'b1_110000000111_101_1_111100000001;
      patterns[57406] = 29'b1_110000000111_110_1_110000000111;
      patterns[57407] = 29'b1_110000000111_111_1_110000000111;
      patterns[57408] = 29'b1_110000001000_000_1_110000001000;
      patterns[57409] = 29'b1_110000001000_001_1_001000110000;
      patterns[57410] = 29'b1_110000001000_010_1_100000010001;
      patterns[57411] = 29'b1_110000001000_011_1_000000100011;
      patterns[57412] = 29'b1_110000001000_100_0_111000000100;
      patterns[57413] = 29'b1_110000001000_101_0_011100000010;
      patterns[57414] = 29'b1_110000001000_110_1_110000001000;
      patterns[57415] = 29'b1_110000001000_111_1_110000001000;
      patterns[57416] = 29'b1_110000001001_000_1_110000001001;
      patterns[57417] = 29'b1_110000001001_001_1_001001110000;
      patterns[57418] = 29'b1_110000001001_010_1_100000010011;
      patterns[57419] = 29'b1_110000001001_011_1_000000100111;
      patterns[57420] = 29'b1_110000001001_100_1_111000000100;
      patterns[57421] = 29'b1_110000001001_101_0_111100000010;
      patterns[57422] = 29'b1_110000001001_110_1_110000001001;
      patterns[57423] = 29'b1_110000001001_111_1_110000001001;
      patterns[57424] = 29'b1_110000001010_000_1_110000001010;
      patterns[57425] = 29'b1_110000001010_001_1_001010110000;
      patterns[57426] = 29'b1_110000001010_010_1_100000010101;
      patterns[57427] = 29'b1_110000001010_011_1_000000101011;
      patterns[57428] = 29'b1_110000001010_100_0_111000000101;
      patterns[57429] = 29'b1_110000001010_101_1_011100000010;
      patterns[57430] = 29'b1_110000001010_110_1_110000001010;
      patterns[57431] = 29'b1_110000001010_111_1_110000001010;
      patterns[57432] = 29'b1_110000001011_000_1_110000001011;
      patterns[57433] = 29'b1_110000001011_001_1_001011110000;
      patterns[57434] = 29'b1_110000001011_010_1_100000010111;
      patterns[57435] = 29'b1_110000001011_011_1_000000101111;
      patterns[57436] = 29'b1_110000001011_100_1_111000000101;
      patterns[57437] = 29'b1_110000001011_101_1_111100000010;
      patterns[57438] = 29'b1_110000001011_110_1_110000001011;
      patterns[57439] = 29'b1_110000001011_111_1_110000001011;
      patterns[57440] = 29'b1_110000001100_000_1_110000001100;
      patterns[57441] = 29'b1_110000001100_001_1_001100110000;
      patterns[57442] = 29'b1_110000001100_010_1_100000011001;
      patterns[57443] = 29'b1_110000001100_011_1_000000110011;
      patterns[57444] = 29'b1_110000001100_100_0_111000000110;
      patterns[57445] = 29'b1_110000001100_101_0_011100000011;
      patterns[57446] = 29'b1_110000001100_110_1_110000001100;
      patterns[57447] = 29'b1_110000001100_111_1_110000001100;
      patterns[57448] = 29'b1_110000001101_000_1_110000001101;
      patterns[57449] = 29'b1_110000001101_001_1_001101110000;
      patterns[57450] = 29'b1_110000001101_010_1_100000011011;
      patterns[57451] = 29'b1_110000001101_011_1_000000110111;
      patterns[57452] = 29'b1_110000001101_100_1_111000000110;
      patterns[57453] = 29'b1_110000001101_101_0_111100000011;
      patterns[57454] = 29'b1_110000001101_110_1_110000001101;
      patterns[57455] = 29'b1_110000001101_111_1_110000001101;
      patterns[57456] = 29'b1_110000001110_000_1_110000001110;
      patterns[57457] = 29'b1_110000001110_001_1_001110110000;
      patterns[57458] = 29'b1_110000001110_010_1_100000011101;
      patterns[57459] = 29'b1_110000001110_011_1_000000111011;
      patterns[57460] = 29'b1_110000001110_100_0_111000000111;
      patterns[57461] = 29'b1_110000001110_101_1_011100000011;
      patterns[57462] = 29'b1_110000001110_110_1_110000001110;
      patterns[57463] = 29'b1_110000001110_111_1_110000001110;
      patterns[57464] = 29'b1_110000001111_000_1_110000001111;
      patterns[57465] = 29'b1_110000001111_001_1_001111110000;
      patterns[57466] = 29'b1_110000001111_010_1_100000011111;
      patterns[57467] = 29'b1_110000001111_011_1_000000111111;
      patterns[57468] = 29'b1_110000001111_100_1_111000000111;
      patterns[57469] = 29'b1_110000001111_101_1_111100000011;
      patterns[57470] = 29'b1_110000001111_110_1_110000001111;
      patterns[57471] = 29'b1_110000001111_111_1_110000001111;
      patterns[57472] = 29'b1_110000010000_000_1_110000010000;
      patterns[57473] = 29'b1_110000010000_001_1_010000110000;
      patterns[57474] = 29'b1_110000010000_010_1_100000100001;
      patterns[57475] = 29'b1_110000010000_011_1_000001000011;
      patterns[57476] = 29'b1_110000010000_100_0_111000001000;
      patterns[57477] = 29'b1_110000010000_101_0_011100000100;
      patterns[57478] = 29'b1_110000010000_110_1_110000010000;
      patterns[57479] = 29'b1_110000010000_111_1_110000010000;
      patterns[57480] = 29'b1_110000010001_000_1_110000010001;
      patterns[57481] = 29'b1_110000010001_001_1_010001110000;
      patterns[57482] = 29'b1_110000010001_010_1_100000100011;
      patterns[57483] = 29'b1_110000010001_011_1_000001000111;
      patterns[57484] = 29'b1_110000010001_100_1_111000001000;
      patterns[57485] = 29'b1_110000010001_101_0_111100000100;
      patterns[57486] = 29'b1_110000010001_110_1_110000010001;
      patterns[57487] = 29'b1_110000010001_111_1_110000010001;
      patterns[57488] = 29'b1_110000010010_000_1_110000010010;
      patterns[57489] = 29'b1_110000010010_001_1_010010110000;
      patterns[57490] = 29'b1_110000010010_010_1_100000100101;
      patterns[57491] = 29'b1_110000010010_011_1_000001001011;
      patterns[57492] = 29'b1_110000010010_100_0_111000001001;
      patterns[57493] = 29'b1_110000010010_101_1_011100000100;
      patterns[57494] = 29'b1_110000010010_110_1_110000010010;
      patterns[57495] = 29'b1_110000010010_111_1_110000010010;
      patterns[57496] = 29'b1_110000010011_000_1_110000010011;
      patterns[57497] = 29'b1_110000010011_001_1_010011110000;
      patterns[57498] = 29'b1_110000010011_010_1_100000100111;
      patterns[57499] = 29'b1_110000010011_011_1_000001001111;
      patterns[57500] = 29'b1_110000010011_100_1_111000001001;
      patterns[57501] = 29'b1_110000010011_101_1_111100000100;
      patterns[57502] = 29'b1_110000010011_110_1_110000010011;
      patterns[57503] = 29'b1_110000010011_111_1_110000010011;
      patterns[57504] = 29'b1_110000010100_000_1_110000010100;
      patterns[57505] = 29'b1_110000010100_001_1_010100110000;
      patterns[57506] = 29'b1_110000010100_010_1_100000101001;
      patterns[57507] = 29'b1_110000010100_011_1_000001010011;
      patterns[57508] = 29'b1_110000010100_100_0_111000001010;
      patterns[57509] = 29'b1_110000010100_101_0_011100000101;
      patterns[57510] = 29'b1_110000010100_110_1_110000010100;
      patterns[57511] = 29'b1_110000010100_111_1_110000010100;
      patterns[57512] = 29'b1_110000010101_000_1_110000010101;
      patterns[57513] = 29'b1_110000010101_001_1_010101110000;
      patterns[57514] = 29'b1_110000010101_010_1_100000101011;
      patterns[57515] = 29'b1_110000010101_011_1_000001010111;
      patterns[57516] = 29'b1_110000010101_100_1_111000001010;
      patterns[57517] = 29'b1_110000010101_101_0_111100000101;
      patterns[57518] = 29'b1_110000010101_110_1_110000010101;
      patterns[57519] = 29'b1_110000010101_111_1_110000010101;
      patterns[57520] = 29'b1_110000010110_000_1_110000010110;
      patterns[57521] = 29'b1_110000010110_001_1_010110110000;
      patterns[57522] = 29'b1_110000010110_010_1_100000101101;
      patterns[57523] = 29'b1_110000010110_011_1_000001011011;
      patterns[57524] = 29'b1_110000010110_100_0_111000001011;
      patterns[57525] = 29'b1_110000010110_101_1_011100000101;
      patterns[57526] = 29'b1_110000010110_110_1_110000010110;
      patterns[57527] = 29'b1_110000010110_111_1_110000010110;
      patterns[57528] = 29'b1_110000010111_000_1_110000010111;
      patterns[57529] = 29'b1_110000010111_001_1_010111110000;
      patterns[57530] = 29'b1_110000010111_010_1_100000101111;
      patterns[57531] = 29'b1_110000010111_011_1_000001011111;
      patterns[57532] = 29'b1_110000010111_100_1_111000001011;
      patterns[57533] = 29'b1_110000010111_101_1_111100000101;
      patterns[57534] = 29'b1_110000010111_110_1_110000010111;
      patterns[57535] = 29'b1_110000010111_111_1_110000010111;
      patterns[57536] = 29'b1_110000011000_000_1_110000011000;
      patterns[57537] = 29'b1_110000011000_001_1_011000110000;
      patterns[57538] = 29'b1_110000011000_010_1_100000110001;
      patterns[57539] = 29'b1_110000011000_011_1_000001100011;
      patterns[57540] = 29'b1_110000011000_100_0_111000001100;
      patterns[57541] = 29'b1_110000011000_101_0_011100000110;
      patterns[57542] = 29'b1_110000011000_110_1_110000011000;
      patterns[57543] = 29'b1_110000011000_111_1_110000011000;
      patterns[57544] = 29'b1_110000011001_000_1_110000011001;
      patterns[57545] = 29'b1_110000011001_001_1_011001110000;
      patterns[57546] = 29'b1_110000011001_010_1_100000110011;
      patterns[57547] = 29'b1_110000011001_011_1_000001100111;
      patterns[57548] = 29'b1_110000011001_100_1_111000001100;
      patterns[57549] = 29'b1_110000011001_101_0_111100000110;
      patterns[57550] = 29'b1_110000011001_110_1_110000011001;
      patterns[57551] = 29'b1_110000011001_111_1_110000011001;
      patterns[57552] = 29'b1_110000011010_000_1_110000011010;
      patterns[57553] = 29'b1_110000011010_001_1_011010110000;
      patterns[57554] = 29'b1_110000011010_010_1_100000110101;
      patterns[57555] = 29'b1_110000011010_011_1_000001101011;
      patterns[57556] = 29'b1_110000011010_100_0_111000001101;
      patterns[57557] = 29'b1_110000011010_101_1_011100000110;
      patterns[57558] = 29'b1_110000011010_110_1_110000011010;
      patterns[57559] = 29'b1_110000011010_111_1_110000011010;
      patterns[57560] = 29'b1_110000011011_000_1_110000011011;
      patterns[57561] = 29'b1_110000011011_001_1_011011110000;
      patterns[57562] = 29'b1_110000011011_010_1_100000110111;
      patterns[57563] = 29'b1_110000011011_011_1_000001101111;
      patterns[57564] = 29'b1_110000011011_100_1_111000001101;
      patterns[57565] = 29'b1_110000011011_101_1_111100000110;
      patterns[57566] = 29'b1_110000011011_110_1_110000011011;
      patterns[57567] = 29'b1_110000011011_111_1_110000011011;
      patterns[57568] = 29'b1_110000011100_000_1_110000011100;
      patterns[57569] = 29'b1_110000011100_001_1_011100110000;
      patterns[57570] = 29'b1_110000011100_010_1_100000111001;
      patterns[57571] = 29'b1_110000011100_011_1_000001110011;
      patterns[57572] = 29'b1_110000011100_100_0_111000001110;
      patterns[57573] = 29'b1_110000011100_101_0_011100000111;
      patterns[57574] = 29'b1_110000011100_110_1_110000011100;
      patterns[57575] = 29'b1_110000011100_111_1_110000011100;
      patterns[57576] = 29'b1_110000011101_000_1_110000011101;
      patterns[57577] = 29'b1_110000011101_001_1_011101110000;
      patterns[57578] = 29'b1_110000011101_010_1_100000111011;
      patterns[57579] = 29'b1_110000011101_011_1_000001110111;
      patterns[57580] = 29'b1_110000011101_100_1_111000001110;
      patterns[57581] = 29'b1_110000011101_101_0_111100000111;
      patterns[57582] = 29'b1_110000011101_110_1_110000011101;
      patterns[57583] = 29'b1_110000011101_111_1_110000011101;
      patterns[57584] = 29'b1_110000011110_000_1_110000011110;
      patterns[57585] = 29'b1_110000011110_001_1_011110110000;
      patterns[57586] = 29'b1_110000011110_010_1_100000111101;
      patterns[57587] = 29'b1_110000011110_011_1_000001111011;
      patterns[57588] = 29'b1_110000011110_100_0_111000001111;
      patterns[57589] = 29'b1_110000011110_101_1_011100000111;
      patterns[57590] = 29'b1_110000011110_110_1_110000011110;
      patterns[57591] = 29'b1_110000011110_111_1_110000011110;
      patterns[57592] = 29'b1_110000011111_000_1_110000011111;
      patterns[57593] = 29'b1_110000011111_001_1_011111110000;
      patterns[57594] = 29'b1_110000011111_010_1_100000111111;
      patterns[57595] = 29'b1_110000011111_011_1_000001111111;
      patterns[57596] = 29'b1_110000011111_100_1_111000001111;
      patterns[57597] = 29'b1_110000011111_101_1_111100000111;
      patterns[57598] = 29'b1_110000011111_110_1_110000011111;
      patterns[57599] = 29'b1_110000011111_111_1_110000011111;
      patterns[57600] = 29'b1_110000100000_000_1_110000100000;
      patterns[57601] = 29'b1_110000100000_001_1_100000110000;
      patterns[57602] = 29'b1_110000100000_010_1_100001000001;
      patterns[57603] = 29'b1_110000100000_011_1_000010000011;
      patterns[57604] = 29'b1_110000100000_100_0_111000010000;
      patterns[57605] = 29'b1_110000100000_101_0_011100001000;
      patterns[57606] = 29'b1_110000100000_110_1_110000100000;
      patterns[57607] = 29'b1_110000100000_111_1_110000100000;
      patterns[57608] = 29'b1_110000100001_000_1_110000100001;
      patterns[57609] = 29'b1_110000100001_001_1_100001110000;
      patterns[57610] = 29'b1_110000100001_010_1_100001000011;
      patterns[57611] = 29'b1_110000100001_011_1_000010000111;
      patterns[57612] = 29'b1_110000100001_100_1_111000010000;
      patterns[57613] = 29'b1_110000100001_101_0_111100001000;
      patterns[57614] = 29'b1_110000100001_110_1_110000100001;
      patterns[57615] = 29'b1_110000100001_111_1_110000100001;
      patterns[57616] = 29'b1_110000100010_000_1_110000100010;
      patterns[57617] = 29'b1_110000100010_001_1_100010110000;
      patterns[57618] = 29'b1_110000100010_010_1_100001000101;
      patterns[57619] = 29'b1_110000100010_011_1_000010001011;
      patterns[57620] = 29'b1_110000100010_100_0_111000010001;
      patterns[57621] = 29'b1_110000100010_101_1_011100001000;
      patterns[57622] = 29'b1_110000100010_110_1_110000100010;
      patterns[57623] = 29'b1_110000100010_111_1_110000100010;
      patterns[57624] = 29'b1_110000100011_000_1_110000100011;
      patterns[57625] = 29'b1_110000100011_001_1_100011110000;
      patterns[57626] = 29'b1_110000100011_010_1_100001000111;
      patterns[57627] = 29'b1_110000100011_011_1_000010001111;
      patterns[57628] = 29'b1_110000100011_100_1_111000010001;
      patterns[57629] = 29'b1_110000100011_101_1_111100001000;
      patterns[57630] = 29'b1_110000100011_110_1_110000100011;
      patterns[57631] = 29'b1_110000100011_111_1_110000100011;
      patterns[57632] = 29'b1_110000100100_000_1_110000100100;
      patterns[57633] = 29'b1_110000100100_001_1_100100110000;
      patterns[57634] = 29'b1_110000100100_010_1_100001001001;
      patterns[57635] = 29'b1_110000100100_011_1_000010010011;
      patterns[57636] = 29'b1_110000100100_100_0_111000010010;
      patterns[57637] = 29'b1_110000100100_101_0_011100001001;
      patterns[57638] = 29'b1_110000100100_110_1_110000100100;
      patterns[57639] = 29'b1_110000100100_111_1_110000100100;
      patterns[57640] = 29'b1_110000100101_000_1_110000100101;
      patterns[57641] = 29'b1_110000100101_001_1_100101110000;
      patterns[57642] = 29'b1_110000100101_010_1_100001001011;
      patterns[57643] = 29'b1_110000100101_011_1_000010010111;
      patterns[57644] = 29'b1_110000100101_100_1_111000010010;
      patterns[57645] = 29'b1_110000100101_101_0_111100001001;
      patterns[57646] = 29'b1_110000100101_110_1_110000100101;
      patterns[57647] = 29'b1_110000100101_111_1_110000100101;
      patterns[57648] = 29'b1_110000100110_000_1_110000100110;
      patterns[57649] = 29'b1_110000100110_001_1_100110110000;
      patterns[57650] = 29'b1_110000100110_010_1_100001001101;
      patterns[57651] = 29'b1_110000100110_011_1_000010011011;
      patterns[57652] = 29'b1_110000100110_100_0_111000010011;
      patterns[57653] = 29'b1_110000100110_101_1_011100001001;
      patterns[57654] = 29'b1_110000100110_110_1_110000100110;
      patterns[57655] = 29'b1_110000100110_111_1_110000100110;
      patterns[57656] = 29'b1_110000100111_000_1_110000100111;
      patterns[57657] = 29'b1_110000100111_001_1_100111110000;
      patterns[57658] = 29'b1_110000100111_010_1_100001001111;
      patterns[57659] = 29'b1_110000100111_011_1_000010011111;
      patterns[57660] = 29'b1_110000100111_100_1_111000010011;
      patterns[57661] = 29'b1_110000100111_101_1_111100001001;
      patterns[57662] = 29'b1_110000100111_110_1_110000100111;
      patterns[57663] = 29'b1_110000100111_111_1_110000100111;
      patterns[57664] = 29'b1_110000101000_000_1_110000101000;
      patterns[57665] = 29'b1_110000101000_001_1_101000110000;
      patterns[57666] = 29'b1_110000101000_010_1_100001010001;
      patterns[57667] = 29'b1_110000101000_011_1_000010100011;
      patterns[57668] = 29'b1_110000101000_100_0_111000010100;
      patterns[57669] = 29'b1_110000101000_101_0_011100001010;
      patterns[57670] = 29'b1_110000101000_110_1_110000101000;
      patterns[57671] = 29'b1_110000101000_111_1_110000101000;
      patterns[57672] = 29'b1_110000101001_000_1_110000101001;
      patterns[57673] = 29'b1_110000101001_001_1_101001110000;
      patterns[57674] = 29'b1_110000101001_010_1_100001010011;
      patterns[57675] = 29'b1_110000101001_011_1_000010100111;
      patterns[57676] = 29'b1_110000101001_100_1_111000010100;
      patterns[57677] = 29'b1_110000101001_101_0_111100001010;
      patterns[57678] = 29'b1_110000101001_110_1_110000101001;
      patterns[57679] = 29'b1_110000101001_111_1_110000101001;
      patterns[57680] = 29'b1_110000101010_000_1_110000101010;
      patterns[57681] = 29'b1_110000101010_001_1_101010110000;
      patterns[57682] = 29'b1_110000101010_010_1_100001010101;
      patterns[57683] = 29'b1_110000101010_011_1_000010101011;
      patterns[57684] = 29'b1_110000101010_100_0_111000010101;
      patterns[57685] = 29'b1_110000101010_101_1_011100001010;
      patterns[57686] = 29'b1_110000101010_110_1_110000101010;
      patterns[57687] = 29'b1_110000101010_111_1_110000101010;
      patterns[57688] = 29'b1_110000101011_000_1_110000101011;
      patterns[57689] = 29'b1_110000101011_001_1_101011110000;
      patterns[57690] = 29'b1_110000101011_010_1_100001010111;
      patterns[57691] = 29'b1_110000101011_011_1_000010101111;
      patterns[57692] = 29'b1_110000101011_100_1_111000010101;
      patterns[57693] = 29'b1_110000101011_101_1_111100001010;
      patterns[57694] = 29'b1_110000101011_110_1_110000101011;
      patterns[57695] = 29'b1_110000101011_111_1_110000101011;
      patterns[57696] = 29'b1_110000101100_000_1_110000101100;
      patterns[57697] = 29'b1_110000101100_001_1_101100110000;
      patterns[57698] = 29'b1_110000101100_010_1_100001011001;
      patterns[57699] = 29'b1_110000101100_011_1_000010110011;
      patterns[57700] = 29'b1_110000101100_100_0_111000010110;
      patterns[57701] = 29'b1_110000101100_101_0_011100001011;
      patterns[57702] = 29'b1_110000101100_110_1_110000101100;
      patterns[57703] = 29'b1_110000101100_111_1_110000101100;
      patterns[57704] = 29'b1_110000101101_000_1_110000101101;
      patterns[57705] = 29'b1_110000101101_001_1_101101110000;
      patterns[57706] = 29'b1_110000101101_010_1_100001011011;
      patterns[57707] = 29'b1_110000101101_011_1_000010110111;
      patterns[57708] = 29'b1_110000101101_100_1_111000010110;
      patterns[57709] = 29'b1_110000101101_101_0_111100001011;
      patterns[57710] = 29'b1_110000101101_110_1_110000101101;
      patterns[57711] = 29'b1_110000101101_111_1_110000101101;
      patterns[57712] = 29'b1_110000101110_000_1_110000101110;
      patterns[57713] = 29'b1_110000101110_001_1_101110110000;
      patterns[57714] = 29'b1_110000101110_010_1_100001011101;
      patterns[57715] = 29'b1_110000101110_011_1_000010111011;
      patterns[57716] = 29'b1_110000101110_100_0_111000010111;
      patterns[57717] = 29'b1_110000101110_101_1_011100001011;
      patterns[57718] = 29'b1_110000101110_110_1_110000101110;
      patterns[57719] = 29'b1_110000101110_111_1_110000101110;
      patterns[57720] = 29'b1_110000101111_000_1_110000101111;
      patterns[57721] = 29'b1_110000101111_001_1_101111110000;
      patterns[57722] = 29'b1_110000101111_010_1_100001011111;
      patterns[57723] = 29'b1_110000101111_011_1_000010111111;
      patterns[57724] = 29'b1_110000101111_100_1_111000010111;
      patterns[57725] = 29'b1_110000101111_101_1_111100001011;
      patterns[57726] = 29'b1_110000101111_110_1_110000101111;
      patterns[57727] = 29'b1_110000101111_111_1_110000101111;
      patterns[57728] = 29'b1_110000110000_000_1_110000110000;
      patterns[57729] = 29'b1_110000110000_001_1_110000110000;
      patterns[57730] = 29'b1_110000110000_010_1_100001100001;
      patterns[57731] = 29'b1_110000110000_011_1_000011000011;
      patterns[57732] = 29'b1_110000110000_100_0_111000011000;
      patterns[57733] = 29'b1_110000110000_101_0_011100001100;
      patterns[57734] = 29'b1_110000110000_110_1_110000110000;
      patterns[57735] = 29'b1_110000110000_111_1_110000110000;
      patterns[57736] = 29'b1_110000110001_000_1_110000110001;
      patterns[57737] = 29'b1_110000110001_001_1_110001110000;
      patterns[57738] = 29'b1_110000110001_010_1_100001100011;
      patterns[57739] = 29'b1_110000110001_011_1_000011000111;
      patterns[57740] = 29'b1_110000110001_100_1_111000011000;
      patterns[57741] = 29'b1_110000110001_101_0_111100001100;
      patterns[57742] = 29'b1_110000110001_110_1_110000110001;
      patterns[57743] = 29'b1_110000110001_111_1_110000110001;
      patterns[57744] = 29'b1_110000110010_000_1_110000110010;
      patterns[57745] = 29'b1_110000110010_001_1_110010110000;
      patterns[57746] = 29'b1_110000110010_010_1_100001100101;
      patterns[57747] = 29'b1_110000110010_011_1_000011001011;
      patterns[57748] = 29'b1_110000110010_100_0_111000011001;
      patterns[57749] = 29'b1_110000110010_101_1_011100001100;
      patterns[57750] = 29'b1_110000110010_110_1_110000110010;
      patterns[57751] = 29'b1_110000110010_111_1_110000110010;
      patterns[57752] = 29'b1_110000110011_000_1_110000110011;
      patterns[57753] = 29'b1_110000110011_001_1_110011110000;
      patterns[57754] = 29'b1_110000110011_010_1_100001100111;
      patterns[57755] = 29'b1_110000110011_011_1_000011001111;
      patterns[57756] = 29'b1_110000110011_100_1_111000011001;
      patterns[57757] = 29'b1_110000110011_101_1_111100001100;
      patterns[57758] = 29'b1_110000110011_110_1_110000110011;
      patterns[57759] = 29'b1_110000110011_111_1_110000110011;
      patterns[57760] = 29'b1_110000110100_000_1_110000110100;
      patterns[57761] = 29'b1_110000110100_001_1_110100110000;
      patterns[57762] = 29'b1_110000110100_010_1_100001101001;
      patterns[57763] = 29'b1_110000110100_011_1_000011010011;
      patterns[57764] = 29'b1_110000110100_100_0_111000011010;
      patterns[57765] = 29'b1_110000110100_101_0_011100001101;
      patterns[57766] = 29'b1_110000110100_110_1_110000110100;
      patterns[57767] = 29'b1_110000110100_111_1_110000110100;
      patterns[57768] = 29'b1_110000110101_000_1_110000110101;
      patterns[57769] = 29'b1_110000110101_001_1_110101110000;
      patterns[57770] = 29'b1_110000110101_010_1_100001101011;
      patterns[57771] = 29'b1_110000110101_011_1_000011010111;
      patterns[57772] = 29'b1_110000110101_100_1_111000011010;
      patterns[57773] = 29'b1_110000110101_101_0_111100001101;
      patterns[57774] = 29'b1_110000110101_110_1_110000110101;
      patterns[57775] = 29'b1_110000110101_111_1_110000110101;
      patterns[57776] = 29'b1_110000110110_000_1_110000110110;
      patterns[57777] = 29'b1_110000110110_001_1_110110110000;
      patterns[57778] = 29'b1_110000110110_010_1_100001101101;
      patterns[57779] = 29'b1_110000110110_011_1_000011011011;
      patterns[57780] = 29'b1_110000110110_100_0_111000011011;
      patterns[57781] = 29'b1_110000110110_101_1_011100001101;
      patterns[57782] = 29'b1_110000110110_110_1_110000110110;
      patterns[57783] = 29'b1_110000110110_111_1_110000110110;
      patterns[57784] = 29'b1_110000110111_000_1_110000110111;
      patterns[57785] = 29'b1_110000110111_001_1_110111110000;
      patterns[57786] = 29'b1_110000110111_010_1_100001101111;
      patterns[57787] = 29'b1_110000110111_011_1_000011011111;
      patterns[57788] = 29'b1_110000110111_100_1_111000011011;
      patterns[57789] = 29'b1_110000110111_101_1_111100001101;
      patterns[57790] = 29'b1_110000110111_110_1_110000110111;
      patterns[57791] = 29'b1_110000110111_111_1_110000110111;
      patterns[57792] = 29'b1_110000111000_000_1_110000111000;
      patterns[57793] = 29'b1_110000111000_001_1_111000110000;
      patterns[57794] = 29'b1_110000111000_010_1_100001110001;
      patterns[57795] = 29'b1_110000111000_011_1_000011100011;
      patterns[57796] = 29'b1_110000111000_100_0_111000011100;
      patterns[57797] = 29'b1_110000111000_101_0_011100001110;
      patterns[57798] = 29'b1_110000111000_110_1_110000111000;
      patterns[57799] = 29'b1_110000111000_111_1_110000111000;
      patterns[57800] = 29'b1_110000111001_000_1_110000111001;
      patterns[57801] = 29'b1_110000111001_001_1_111001110000;
      patterns[57802] = 29'b1_110000111001_010_1_100001110011;
      patterns[57803] = 29'b1_110000111001_011_1_000011100111;
      patterns[57804] = 29'b1_110000111001_100_1_111000011100;
      patterns[57805] = 29'b1_110000111001_101_0_111100001110;
      patterns[57806] = 29'b1_110000111001_110_1_110000111001;
      patterns[57807] = 29'b1_110000111001_111_1_110000111001;
      patterns[57808] = 29'b1_110000111010_000_1_110000111010;
      patterns[57809] = 29'b1_110000111010_001_1_111010110000;
      patterns[57810] = 29'b1_110000111010_010_1_100001110101;
      patterns[57811] = 29'b1_110000111010_011_1_000011101011;
      patterns[57812] = 29'b1_110000111010_100_0_111000011101;
      patterns[57813] = 29'b1_110000111010_101_1_011100001110;
      patterns[57814] = 29'b1_110000111010_110_1_110000111010;
      patterns[57815] = 29'b1_110000111010_111_1_110000111010;
      patterns[57816] = 29'b1_110000111011_000_1_110000111011;
      patterns[57817] = 29'b1_110000111011_001_1_111011110000;
      patterns[57818] = 29'b1_110000111011_010_1_100001110111;
      patterns[57819] = 29'b1_110000111011_011_1_000011101111;
      patterns[57820] = 29'b1_110000111011_100_1_111000011101;
      patterns[57821] = 29'b1_110000111011_101_1_111100001110;
      patterns[57822] = 29'b1_110000111011_110_1_110000111011;
      patterns[57823] = 29'b1_110000111011_111_1_110000111011;
      patterns[57824] = 29'b1_110000111100_000_1_110000111100;
      patterns[57825] = 29'b1_110000111100_001_1_111100110000;
      patterns[57826] = 29'b1_110000111100_010_1_100001111001;
      patterns[57827] = 29'b1_110000111100_011_1_000011110011;
      patterns[57828] = 29'b1_110000111100_100_0_111000011110;
      patterns[57829] = 29'b1_110000111100_101_0_011100001111;
      patterns[57830] = 29'b1_110000111100_110_1_110000111100;
      patterns[57831] = 29'b1_110000111100_111_1_110000111100;
      patterns[57832] = 29'b1_110000111101_000_1_110000111101;
      patterns[57833] = 29'b1_110000111101_001_1_111101110000;
      patterns[57834] = 29'b1_110000111101_010_1_100001111011;
      patterns[57835] = 29'b1_110000111101_011_1_000011110111;
      patterns[57836] = 29'b1_110000111101_100_1_111000011110;
      patterns[57837] = 29'b1_110000111101_101_0_111100001111;
      patterns[57838] = 29'b1_110000111101_110_1_110000111101;
      patterns[57839] = 29'b1_110000111101_111_1_110000111101;
      patterns[57840] = 29'b1_110000111110_000_1_110000111110;
      patterns[57841] = 29'b1_110000111110_001_1_111110110000;
      patterns[57842] = 29'b1_110000111110_010_1_100001111101;
      patterns[57843] = 29'b1_110000111110_011_1_000011111011;
      patterns[57844] = 29'b1_110000111110_100_0_111000011111;
      patterns[57845] = 29'b1_110000111110_101_1_011100001111;
      patterns[57846] = 29'b1_110000111110_110_1_110000111110;
      patterns[57847] = 29'b1_110000111110_111_1_110000111110;
      patterns[57848] = 29'b1_110000111111_000_1_110000111111;
      patterns[57849] = 29'b1_110000111111_001_1_111111110000;
      patterns[57850] = 29'b1_110000111111_010_1_100001111111;
      patterns[57851] = 29'b1_110000111111_011_1_000011111111;
      patterns[57852] = 29'b1_110000111111_100_1_111000011111;
      patterns[57853] = 29'b1_110000111111_101_1_111100001111;
      patterns[57854] = 29'b1_110000111111_110_1_110000111111;
      patterns[57855] = 29'b1_110000111111_111_1_110000111111;
      patterns[57856] = 29'b1_110001000000_000_1_110001000000;
      patterns[57857] = 29'b1_110001000000_001_1_000000110001;
      patterns[57858] = 29'b1_110001000000_010_1_100010000001;
      patterns[57859] = 29'b1_110001000000_011_1_000100000011;
      patterns[57860] = 29'b1_110001000000_100_0_111000100000;
      patterns[57861] = 29'b1_110001000000_101_0_011100010000;
      patterns[57862] = 29'b1_110001000000_110_1_110001000000;
      patterns[57863] = 29'b1_110001000000_111_1_110001000000;
      patterns[57864] = 29'b1_110001000001_000_1_110001000001;
      patterns[57865] = 29'b1_110001000001_001_1_000001110001;
      patterns[57866] = 29'b1_110001000001_010_1_100010000011;
      patterns[57867] = 29'b1_110001000001_011_1_000100000111;
      patterns[57868] = 29'b1_110001000001_100_1_111000100000;
      patterns[57869] = 29'b1_110001000001_101_0_111100010000;
      patterns[57870] = 29'b1_110001000001_110_1_110001000001;
      patterns[57871] = 29'b1_110001000001_111_1_110001000001;
      patterns[57872] = 29'b1_110001000010_000_1_110001000010;
      patterns[57873] = 29'b1_110001000010_001_1_000010110001;
      patterns[57874] = 29'b1_110001000010_010_1_100010000101;
      patterns[57875] = 29'b1_110001000010_011_1_000100001011;
      patterns[57876] = 29'b1_110001000010_100_0_111000100001;
      patterns[57877] = 29'b1_110001000010_101_1_011100010000;
      patterns[57878] = 29'b1_110001000010_110_1_110001000010;
      patterns[57879] = 29'b1_110001000010_111_1_110001000010;
      patterns[57880] = 29'b1_110001000011_000_1_110001000011;
      patterns[57881] = 29'b1_110001000011_001_1_000011110001;
      patterns[57882] = 29'b1_110001000011_010_1_100010000111;
      patterns[57883] = 29'b1_110001000011_011_1_000100001111;
      patterns[57884] = 29'b1_110001000011_100_1_111000100001;
      patterns[57885] = 29'b1_110001000011_101_1_111100010000;
      patterns[57886] = 29'b1_110001000011_110_1_110001000011;
      patterns[57887] = 29'b1_110001000011_111_1_110001000011;
      patterns[57888] = 29'b1_110001000100_000_1_110001000100;
      patterns[57889] = 29'b1_110001000100_001_1_000100110001;
      patterns[57890] = 29'b1_110001000100_010_1_100010001001;
      patterns[57891] = 29'b1_110001000100_011_1_000100010011;
      patterns[57892] = 29'b1_110001000100_100_0_111000100010;
      patterns[57893] = 29'b1_110001000100_101_0_011100010001;
      patterns[57894] = 29'b1_110001000100_110_1_110001000100;
      patterns[57895] = 29'b1_110001000100_111_1_110001000100;
      patterns[57896] = 29'b1_110001000101_000_1_110001000101;
      patterns[57897] = 29'b1_110001000101_001_1_000101110001;
      patterns[57898] = 29'b1_110001000101_010_1_100010001011;
      patterns[57899] = 29'b1_110001000101_011_1_000100010111;
      patterns[57900] = 29'b1_110001000101_100_1_111000100010;
      patterns[57901] = 29'b1_110001000101_101_0_111100010001;
      patterns[57902] = 29'b1_110001000101_110_1_110001000101;
      patterns[57903] = 29'b1_110001000101_111_1_110001000101;
      patterns[57904] = 29'b1_110001000110_000_1_110001000110;
      patterns[57905] = 29'b1_110001000110_001_1_000110110001;
      patterns[57906] = 29'b1_110001000110_010_1_100010001101;
      patterns[57907] = 29'b1_110001000110_011_1_000100011011;
      patterns[57908] = 29'b1_110001000110_100_0_111000100011;
      patterns[57909] = 29'b1_110001000110_101_1_011100010001;
      patterns[57910] = 29'b1_110001000110_110_1_110001000110;
      patterns[57911] = 29'b1_110001000110_111_1_110001000110;
      patterns[57912] = 29'b1_110001000111_000_1_110001000111;
      patterns[57913] = 29'b1_110001000111_001_1_000111110001;
      patterns[57914] = 29'b1_110001000111_010_1_100010001111;
      patterns[57915] = 29'b1_110001000111_011_1_000100011111;
      patterns[57916] = 29'b1_110001000111_100_1_111000100011;
      patterns[57917] = 29'b1_110001000111_101_1_111100010001;
      patterns[57918] = 29'b1_110001000111_110_1_110001000111;
      patterns[57919] = 29'b1_110001000111_111_1_110001000111;
      patterns[57920] = 29'b1_110001001000_000_1_110001001000;
      patterns[57921] = 29'b1_110001001000_001_1_001000110001;
      patterns[57922] = 29'b1_110001001000_010_1_100010010001;
      patterns[57923] = 29'b1_110001001000_011_1_000100100011;
      patterns[57924] = 29'b1_110001001000_100_0_111000100100;
      patterns[57925] = 29'b1_110001001000_101_0_011100010010;
      patterns[57926] = 29'b1_110001001000_110_1_110001001000;
      patterns[57927] = 29'b1_110001001000_111_1_110001001000;
      patterns[57928] = 29'b1_110001001001_000_1_110001001001;
      patterns[57929] = 29'b1_110001001001_001_1_001001110001;
      patterns[57930] = 29'b1_110001001001_010_1_100010010011;
      patterns[57931] = 29'b1_110001001001_011_1_000100100111;
      patterns[57932] = 29'b1_110001001001_100_1_111000100100;
      patterns[57933] = 29'b1_110001001001_101_0_111100010010;
      patterns[57934] = 29'b1_110001001001_110_1_110001001001;
      patterns[57935] = 29'b1_110001001001_111_1_110001001001;
      patterns[57936] = 29'b1_110001001010_000_1_110001001010;
      patterns[57937] = 29'b1_110001001010_001_1_001010110001;
      patterns[57938] = 29'b1_110001001010_010_1_100010010101;
      patterns[57939] = 29'b1_110001001010_011_1_000100101011;
      patterns[57940] = 29'b1_110001001010_100_0_111000100101;
      patterns[57941] = 29'b1_110001001010_101_1_011100010010;
      patterns[57942] = 29'b1_110001001010_110_1_110001001010;
      patterns[57943] = 29'b1_110001001010_111_1_110001001010;
      patterns[57944] = 29'b1_110001001011_000_1_110001001011;
      patterns[57945] = 29'b1_110001001011_001_1_001011110001;
      patterns[57946] = 29'b1_110001001011_010_1_100010010111;
      patterns[57947] = 29'b1_110001001011_011_1_000100101111;
      patterns[57948] = 29'b1_110001001011_100_1_111000100101;
      patterns[57949] = 29'b1_110001001011_101_1_111100010010;
      patterns[57950] = 29'b1_110001001011_110_1_110001001011;
      patterns[57951] = 29'b1_110001001011_111_1_110001001011;
      patterns[57952] = 29'b1_110001001100_000_1_110001001100;
      patterns[57953] = 29'b1_110001001100_001_1_001100110001;
      patterns[57954] = 29'b1_110001001100_010_1_100010011001;
      patterns[57955] = 29'b1_110001001100_011_1_000100110011;
      patterns[57956] = 29'b1_110001001100_100_0_111000100110;
      patterns[57957] = 29'b1_110001001100_101_0_011100010011;
      patterns[57958] = 29'b1_110001001100_110_1_110001001100;
      patterns[57959] = 29'b1_110001001100_111_1_110001001100;
      patterns[57960] = 29'b1_110001001101_000_1_110001001101;
      patterns[57961] = 29'b1_110001001101_001_1_001101110001;
      patterns[57962] = 29'b1_110001001101_010_1_100010011011;
      patterns[57963] = 29'b1_110001001101_011_1_000100110111;
      patterns[57964] = 29'b1_110001001101_100_1_111000100110;
      patterns[57965] = 29'b1_110001001101_101_0_111100010011;
      patterns[57966] = 29'b1_110001001101_110_1_110001001101;
      patterns[57967] = 29'b1_110001001101_111_1_110001001101;
      patterns[57968] = 29'b1_110001001110_000_1_110001001110;
      patterns[57969] = 29'b1_110001001110_001_1_001110110001;
      patterns[57970] = 29'b1_110001001110_010_1_100010011101;
      patterns[57971] = 29'b1_110001001110_011_1_000100111011;
      patterns[57972] = 29'b1_110001001110_100_0_111000100111;
      patterns[57973] = 29'b1_110001001110_101_1_011100010011;
      patterns[57974] = 29'b1_110001001110_110_1_110001001110;
      patterns[57975] = 29'b1_110001001110_111_1_110001001110;
      patterns[57976] = 29'b1_110001001111_000_1_110001001111;
      patterns[57977] = 29'b1_110001001111_001_1_001111110001;
      patterns[57978] = 29'b1_110001001111_010_1_100010011111;
      patterns[57979] = 29'b1_110001001111_011_1_000100111111;
      patterns[57980] = 29'b1_110001001111_100_1_111000100111;
      patterns[57981] = 29'b1_110001001111_101_1_111100010011;
      patterns[57982] = 29'b1_110001001111_110_1_110001001111;
      patterns[57983] = 29'b1_110001001111_111_1_110001001111;
      patterns[57984] = 29'b1_110001010000_000_1_110001010000;
      patterns[57985] = 29'b1_110001010000_001_1_010000110001;
      patterns[57986] = 29'b1_110001010000_010_1_100010100001;
      patterns[57987] = 29'b1_110001010000_011_1_000101000011;
      patterns[57988] = 29'b1_110001010000_100_0_111000101000;
      patterns[57989] = 29'b1_110001010000_101_0_011100010100;
      patterns[57990] = 29'b1_110001010000_110_1_110001010000;
      patterns[57991] = 29'b1_110001010000_111_1_110001010000;
      patterns[57992] = 29'b1_110001010001_000_1_110001010001;
      patterns[57993] = 29'b1_110001010001_001_1_010001110001;
      patterns[57994] = 29'b1_110001010001_010_1_100010100011;
      patterns[57995] = 29'b1_110001010001_011_1_000101000111;
      patterns[57996] = 29'b1_110001010001_100_1_111000101000;
      patterns[57997] = 29'b1_110001010001_101_0_111100010100;
      patterns[57998] = 29'b1_110001010001_110_1_110001010001;
      patterns[57999] = 29'b1_110001010001_111_1_110001010001;
      patterns[58000] = 29'b1_110001010010_000_1_110001010010;
      patterns[58001] = 29'b1_110001010010_001_1_010010110001;
      patterns[58002] = 29'b1_110001010010_010_1_100010100101;
      patterns[58003] = 29'b1_110001010010_011_1_000101001011;
      patterns[58004] = 29'b1_110001010010_100_0_111000101001;
      patterns[58005] = 29'b1_110001010010_101_1_011100010100;
      patterns[58006] = 29'b1_110001010010_110_1_110001010010;
      patterns[58007] = 29'b1_110001010010_111_1_110001010010;
      patterns[58008] = 29'b1_110001010011_000_1_110001010011;
      patterns[58009] = 29'b1_110001010011_001_1_010011110001;
      patterns[58010] = 29'b1_110001010011_010_1_100010100111;
      patterns[58011] = 29'b1_110001010011_011_1_000101001111;
      patterns[58012] = 29'b1_110001010011_100_1_111000101001;
      patterns[58013] = 29'b1_110001010011_101_1_111100010100;
      patterns[58014] = 29'b1_110001010011_110_1_110001010011;
      patterns[58015] = 29'b1_110001010011_111_1_110001010011;
      patterns[58016] = 29'b1_110001010100_000_1_110001010100;
      patterns[58017] = 29'b1_110001010100_001_1_010100110001;
      patterns[58018] = 29'b1_110001010100_010_1_100010101001;
      patterns[58019] = 29'b1_110001010100_011_1_000101010011;
      patterns[58020] = 29'b1_110001010100_100_0_111000101010;
      patterns[58021] = 29'b1_110001010100_101_0_011100010101;
      patterns[58022] = 29'b1_110001010100_110_1_110001010100;
      patterns[58023] = 29'b1_110001010100_111_1_110001010100;
      patterns[58024] = 29'b1_110001010101_000_1_110001010101;
      patterns[58025] = 29'b1_110001010101_001_1_010101110001;
      patterns[58026] = 29'b1_110001010101_010_1_100010101011;
      patterns[58027] = 29'b1_110001010101_011_1_000101010111;
      patterns[58028] = 29'b1_110001010101_100_1_111000101010;
      patterns[58029] = 29'b1_110001010101_101_0_111100010101;
      patterns[58030] = 29'b1_110001010101_110_1_110001010101;
      patterns[58031] = 29'b1_110001010101_111_1_110001010101;
      patterns[58032] = 29'b1_110001010110_000_1_110001010110;
      patterns[58033] = 29'b1_110001010110_001_1_010110110001;
      patterns[58034] = 29'b1_110001010110_010_1_100010101101;
      patterns[58035] = 29'b1_110001010110_011_1_000101011011;
      patterns[58036] = 29'b1_110001010110_100_0_111000101011;
      patterns[58037] = 29'b1_110001010110_101_1_011100010101;
      patterns[58038] = 29'b1_110001010110_110_1_110001010110;
      patterns[58039] = 29'b1_110001010110_111_1_110001010110;
      patterns[58040] = 29'b1_110001010111_000_1_110001010111;
      patterns[58041] = 29'b1_110001010111_001_1_010111110001;
      patterns[58042] = 29'b1_110001010111_010_1_100010101111;
      patterns[58043] = 29'b1_110001010111_011_1_000101011111;
      patterns[58044] = 29'b1_110001010111_100_1_111000101011;
      patterns[58045] = 29'b1_110001010111_101_1_111100010101;
      patterns[58046] = 29'b1_110001010111_110_1_110001010111;
      patterns[58047] = 29'b1_110001010111_111_1_110001010111;
      patterns[58048] = 29'b1_110001011000_000_1_110001011000;
      patterns[58049] = 29'b1_110001011000_001_1_011000110001;
      patterns[58050] = 29'b1_110001011000_010_1_100010110001;
      patterns[58051] = 29'b1_110001011000_011_1_000101100011;
      patterns[58052] = 29'b1_110001011000_100_0_111000101100;
      patterns[58053] = 29'b1_110001011000_101_0_011100010110;
      patterns[58054] = 29'b1_110001011000_110_1_110001011000;
      patterns[58055] = 29'b1_110001011000_111_1_110001011000;
      patterns[58056] = 29'b1_110001011001_000_1_110001011001;
      patterns[58057] = 29'b1_110001011001_001_1_011001110001;
      patterns[58058] = 29'b1_110001011001_010_1_100010110011;
      patterns[58059] = 29'b1_110001011001_011_1_000101100111;
      patterns[58060] = 29'b1_110001011001_100_1_111000101100;
      patterns[58061] = 29'b1_110001011001_101_0_111100010110;
      patterns[58062] = 29'b1_110001011001_110_1_110001011001;
      patterns[58063] = 29'b1_110001011001_111_1_110001011001;
      patterns[58064] = 29'b1_110001011010_000_1_110001011010;
      patterns[58065] = 29'b1_110001011010_001_1_011010110001;
      patterns[58066] = 29'b1_110001011010_010_1_100010110101;
      patterns[58067] = 29'b1_110001011010_011_1_000101101011;
      patterns[58068] = 29'b1_110001011010_100_0_111000101101;
      patterns[58069] = 29'b1_110001011010_101_1_011100010110;
      patterns[58070] = 29'b1_110001011010_110_1_110001011010;
      patterns[58071] = 29'b1_110001011010_111_1_110001011010;
      patterns[58072] = 29'b1_110001011011_000_1_110001011011;
      patterns[58073] = 29'b1_110001011011_001_1_011011110001;
      patterns[58074] = 29'b1_110001011011_010_1_100010110111;
      patterns[58075] = 29'b1_110001011011_011_1_000101101111;
      patterns[58076] = 29'b1_110001011011_100_1_111000101101;
      patterns[58077] = 29'b1_110001011011_101_1_111100010110;
      patterns[58078] = 29'b1_110001011011_110_1_110001011011;
      patterns[58079] = 29'b1_110001011011_111_1_110001011011;
      patterns[58080] = 29'b1_110001011100_000_1_110001011100;
      patterns[58081] = 29'b1_110001011100_001_1_011100110001;
      patterns[58082] = 29'b1_110001011100_010_1_100010111001;
      patterns[58083] = 29'b1_110001011100_011_1_000101110011;
      patterns[58084] = 29'b1_110001011100_100_0_111000101110;
      patterns[58085] = 29'b1_110001011100_101_0_011100010111;
      patterns[58086] = 29'b1_110001011100_110_1_110001011100;
      patterns[58087] = 29'b1_110001011100_111_1_110001011100;
      patterns[58088] = 29'b1_110001011101_000_1_110001011101;
      patterns[58089] = 29'b1_110001011101_001_1_011101110001;
      patterns[58090] = 29'b1_110001011101_010_1_100010111011;
      patterns[58091] = 29'b1_110001011101_011_1_000101110111;
      patterns[58092] = 29'b1_110001011101_100_1_111000101110;
      patterns[58093] = 29'b1_110001011101_101_0_111100010111;
      patterns[58094] = 29'b1_110001011101_110_1_110001011101;
      patterns[58095] = 29'b1_110001011101_111_1_110001011101;
      patterns[58096] = 29'b1_110001011110_000_1_110001011110;
      patterns[58097] = 29'b1_110001011110_001_1_011110110001;
      patterns[58098] = 29'b1_110001011110_010_1_100010111101;
      patterns[58099] = 29'b1_110001011110_011_1_000101111011;
      patterns[58100] = 29'b1_110001011110_100_0_111000101111;
      patterns[58101] = 29'b1_110001011110_101_1_011100010111;
      patterns[58102] = 29'b1_110001011110_110_1_110001011110;
      patterns[58103] = 29'b1_110001011110_111_1_110001011110;
      patterns[58104] = 29'b1_110001011111_000_1_110001011111;
      patterns[58105] = 29'b1_110001011111_001_1_011111110001;
      patterns[58106] = 29'b1_110001011111_010_1_100010111111;
      patterns[58107] = 29'b1_110001011111_011_1_000101111111;
      patterns[58108] = 29'b1_110001011111_100_1_111000101111;
      patterns[58109] = 29'b1_110001011111_101_1_111100010111;
      patterns[58110] = 29'b1_110001011111_110_1_110001011111;
      patterns[58111] = 29'b1_110001011111_111_1_110001011111;
      patterns[58112] = 29'b1_110001100000_000_1_110001100000;
      patterns[58113] = 29'b1_110001100000_001_1_100000110001;
      patterns[58114] = 29'b1_110001100000_010_1_100011000001;
      patterns[58115] = 29'b1_110001100000_011_1_000110000011;
      patterns[58116] = 29'b1_110001100000_100_0_111000110000;
      patterns[58117] = 29'b1_110001100000_101_0_011100011000;
      patterns[58118] = 29'b1_110001100000_110_1_110001100000;
      patterns[58119] = 29'b1_110001100000_111_1_110001100000;
      patterns[58120] = 29'b1_110001100001_000_1_110001100001;
      patterns[58121] = 29'b1_110001100001_001_1_100001110001;
      patterns[58122] = 29'b1_110001100001_010_1_100011000011;
      patterns[58123] = 29'b1_110001100001_011_1_000110000111;
      patterns[58124] = 29'b1_110001100001_100_1_111000110000;
      patterns[58125] = 29'b1_110001100001_101_0_111100011000;
      patterns[58126] = 29'b1_110001100001_110_1_110001100001;
      patterns[58127] = 29'b1_110001100001_111_1_110001100001;
      patterns[58128] = 29'b1_110001100010_000_1_110001100010;
      patterns[58129] = 29'b1_110001100010_001_1_100010110001;
      patterns[58130] = 29'b1_110001100010_010_1_100011000101;
      patterns[58131] = 29'b1_110001100010_011_1_000110001011;
      patterns[58132] = 29'b1_110001100010_100_0_111000110001;
      patterns[58133] = 29'b1_110001100010_101_1_011100011000;
      patterns[58134] = 29'b1_110001100010_110_1_110001100010;
      patterns[58135] = 29'b1_110001100010_111_1_110001100010;
      patterns[58136] = 29'b1_110001100011_000_1_110001100011;
      patterns[58137] = 29'b1_110001100011_001_1_100011110001;
      patterns[58138] = 29'b1_110001100011_010_1_100011000111;
      patterns[58139] = 29'b1_110001100011_011_1_000110001111;
      patterns[58140] = 29'b1_110001100011_100_1_111000110001;
      patterns[58141] = 29'b1_110001100011_101_1_111100011000;
      patterns[58142] = 29'b1_110001100011_110_1_110001100011;
      patterns[58143] = 29'b1_110001100011_111_1_110001100011;
      patterns[58144] = 29'b1_110001100100_000_1_110001100100;
      patterns[58145] = 29'b1_110001100100_001_1_100100110001;
      patterns[58146] = 29'b1_110001100100_010_1_100011001001;
      patterns[58147] = 29'b1_110001100100_011_1_000110010011;
      patterns[58148] = 29'b1_110001100100_100_0_111000110010;
      patterns[58149] = 29'b1_110001100100_101_0_011100011001;
      patterns[58150] = 29'b1_110001100100_110_1_110001100100;
      patterns[58151] = 29'b1_110001100100_111_1_110001100100;
      patterns[58152] = 29'b1_110001100101_000_1_110001100101;
      patterns[58153] = 29'b1_110001100101_001_1_100101110001;
      patterns[58154] = 29'b1_110001100101_010_1_100011001011;
      patterns[58155] = 29'b1_110001100101_011_1_000110010111;
      patterns[58156] = 29'b1_110001100101_100_1_111000110010;
      patterns[58157] = 29'b1_110001100101_101_0_111100011001;
      patterns[58158] = 29'b1_110001100101_110_1_110001100101;
      patterns[58159] = 29'b1_110001100101_111_1_110001100101;
      patterns[58160] = 29'b1_110001100110_000_1_110001100110;
      patterns[58161] = 29'b1_110001100110_001_1_100110110001;
      patterns[58162] = 29'b1_110001100110_010_1_100011001101;
      patterns[58163] = 29'b1_110001100110_011_1_000110011011;
      patterns[58164] = 29'b1_110001100110_100_0_111000110011;
      patterns[58165] = 29'b1_110001100110_101_1_011100011001;
      patterns[58166] = 29'b1_110001100110_110_1_110001100110;
      patterns[58167] = 29'b1_110001100110_111_1_110001100110;
      patterns[58168] = 29'b1_110001100111_000_1_110001100111;
      patterns[58169] = 29'b1_110001100111_001_1_100111110001;
      patterns[58170] = 29'b1_110001100111_010_1_100011001111;
      patterns[58171] = 29'b1_110001100111_011_1_000110011111;
      patterns[58172] = 29'b1_110001100111_100_1_111000110011;
      patterns[58173] = 29'b1_110001100111_101_1_111100011001;
      patterns[58174] = 29'b1_110001100111_110_1_110001100111;
      patterns[58175] = 29'b1_110001100111_111_1_110001100111;
      patterns[58176] = 29'b1_110001101000_000_1_110001101000;
      patterns[58177] = 29'b1_110001101000_001_1_101000110001;
      patterns[58178] = 29'b1_110001101000_010_1_100011010001;
      patterns[58179] = 29'b1_110001101000_011_1_000110100011;
      patterns[58180] = 29'b1_110001101000_100_0_111000110100;
      patterns[58181] = 29'b1_110001101000_101_0_011100011010;
      patterns[58182] = 29'b1_110001101000_110_1_110001101000;
      patterns[58183] = 29'b1_110001101000_111_1_110001101000;
      patterns[58184] = 29'b1_110001101001_000_1_110001101001;
      patterns[58185] = 29'b1_110001101001_001_1_101001110001;
      patterns[58186] = 29'b1_110001101001_010_1_100011010011;
      patterns[58187] = 29'b1_110001101001_011_1_000110100111;
      patterns[58188] = 29'b1_110001101001_100_1_111000110100;
      patterns[58189] = 29'b1_110001101001_101_0_111100011010;
      patterns[58190] = 29'b1_110001101001_110_1_110001101001;
      patterns[58191] = 29'b1_110001101001_111_1_110001101001;
      patterns[58192] = 29'b1_110001101010_000_1_110001101010;
      patterns[58193] = 29'b1_110001101010_001_1_101010110001;
      patterns[58194] = 29'b1_110001101010_010_1_100011010101;
      patterns[58195] = 29'b1_110001101010_011_1_000110101011;
      patterns[58196] = 29'b1_110001101010_100_0_111000110101;
      patterns[58197] = 29'b1_110001101010_101_1_011100011010;
      patterns[58198] = 29'b1_110001101010_110_1_110001101010;
      patterns[58199] = 29'b1_110001101010_111_1_110001101010;
      patterns[58200] = 29'b1_110001101011_000_1_110001101011;
      patterns[58201] = 29'b1_110001101011_001_1_101011110001;
      patterns[58202] = 29'b1_110001101011_010_1_100011010111;
      patterns[58203] = 29'b1_110001101011_011_1_000110101111;
      patterns[58204] = 29'b1_110001101011_100_1_111000110101;
      patterns[58205] = 29'b1_110001101011_101_1_111100011010;
      patterns[58206] = 29'b1_110001101011_110_1_110001101011;
      patterns[58207] = 29'b1_110001101011_111_1_110001101011;
      patterns[58208] = 29'b1_110001101100_000_1_110001101100;
      patterns[58209] = 29'b1_110001101100_001_1_101100110001;
      patterns[58210] = 29'b1_110001101100_010_1_100011011001;
      patterns[58211] = 29'b1_110001101100_011_1_000110110011;
      patterns[58212] = 29'b1_110001101100_100_0_111000110110;
      patterns[58213] = 29'b1_110001101100_101_0_011100011011;
      patterns[58214] = 29'b1_110001101100_110_1_110001101100;
      patterns[58215] = 29'b1_110001101100_111_1_110001101100;
      patterns[58216] = 29'b1_110001101101_000_1_110001101101;
      patterns[58217] = 29'b1_110001101101_001_1_101101110001;
      patterns[58218] = 29'b1_110001101101_010_1_100011011011;
      patterns[58219] = 29'b1_110001101101_011_1_000110110111;
      patterns[58220] = 29'b1_110001101101_100_1_111000110110;
      patterns[58221] = 29'b1_110001101101_101_0_111100011011;
      patterns[58222] = 29'b1_110001101101_110_1_110001101101;
      patterns[58223] = 29'b1_110001101101_111_1_110001101101;
      patterns[58224] = 29'b1_110001101110_000_1_110001101110;
      patterns[58225] = 29'b1_110001101110_001_1_101110110001;
      patterns[58226] = 29'b1_110001101110_010_1_100011011101;
      patterns[58227] = 29'b1_110001101110_011_1_000110111011;
      patterns[58228] = 29'b1_110001101110_100_0_111000110111;
      patterns[58229] = 29'b1_110001101110_101_1_011100011011;
      patterns[58230] = 29'b1_110001101110_110_1_110001101110;
      patterns[58231] = 29'b1_110001101110_111_1_110001101110;
      patterns[58232] = 29'b1_110001101111_000_1_110001101111;
      patterns[58233] = 29'b1_110001101111_001_1_101111110001;
      patterns[58234] = 29'b1_110001101111_010_1_100011011111;
      patterns[58235] = 29'b1_110001101111_011_1_000110111111;
      patterns[58236] = 29'b1_110001101111_100_1_111000110111;
      patterns[58237] = 29'b1_110001101111_101_1_111100011011;
      patterns[58238] = 29'b1_110001101111_110_1_110001101111;
      patterns[58239] = 29'b1_110001101111_111_1_110001101111;
      patterns[58240] = 29'b1_110001110000_000_1_110001110000;
      patterns[58241] = 29'b1_110001110000_001_1_110000110001;
      patterns[58242] = 29'b1_110001110000_010_1_100011100001;
      patterns[58243] = 29'b1_110001110000_011_1_000111000011;
      patterns[58244] = 29'b1_110001110000_100_0_111000111000;
      patterns[58245] = 29'b1_110001110000_101_0_011100011100;
      patterns[58246] = 29'b1_110001110000_110_1_110001110000;
      patterns[58247] = 29'b1_110001110000_111_1_110001110000;
      patterns[58248] = 29'b1_110001110001_000_1_110001110001;
      patterns[58249] = 29'b1_110001110001_001_1_110001110001;
      patterns[58250] = 29'b1_110001110001_010_1_100011100011;
      patterns[58251] = 29'b1_110001110001_011_1_000111000111;
      patterns[58252] = 29'b1_110001110001_100_1_111000111000;
      patterns[58253] = 29'b1_110001110001_101_0_111100011100;
      patterns[58254] = 29'b1_110001110001_110_1_110001110001;
      patterns[58255] = 29'b1_110001110001_111_1_110001110001;
      patterns[58256] = 29'b1_110001110010_000_1_110001110010;
      patterns[58257] = 29'b1_110001110010_001_1_110010110001;
      patterns[58258] = 29'b1_110001110010_010_1_100011100101;
      patterns[58259] = 29'b1_110001110010_011_1_000111001011;
      patterns[58260] = 29'b1_110001110010_100_0_111000111001;
      patterns[58261] = 29'b1_110001110010_101_1_011100011100;
      patterns[58262] = 29'b1_110001110010_110_1_110001110010;
      patterns[58263] = 29'b1_110001110010_111_1_110001110010;
      patterns[58264] = 29'b1_110001110011_000_1_110001110011;
      patterns[58265] = 29'b1_110001110011_001_1_110011110001;
      patterns[58266] = 29'b1_110001110011_010_1_100011100111;
      patterns[58267] = 29'b1_110001110011_011_1_000111001111;
      patterns[58268] = 29'b1_110001110011_100_1_111000111001;
      patterns[58269] = 29'b1_110001110011_101_1_111100011100;
      patterns[58270] = 29'b1_110001110011_110_1_110001110011;
      patterns[58271] = 29'b1_110001110011_111_1_110001110011;
      patterns[58272] = 29'b1_110001110100_000_1_110001110100;
      patterns[58273] = 29'b1_110001110100_001_1_110100110001;
      patterns[58274] = 29'b1_110001110100_010_1_100011101001;
      patterns[58275] = 29'b1_110001110100_011_1_000111010011;
      patterns[58276] = 29'b1_110001110100_100_0_111000111010;
      patterns[58277] = 29'b1_110001110100_101_0_011100011101;
      patterns[58278] = 29'b1_110001110100_110_1_110001110100;
      patterns[58279] = 29'b1_110001110100_111_1_110001110100;
      patterns[58280] = 29'b1_110001110101_000_1_110001110101;
      patterns[58281] = 29'b1_110001110101_001_1_110101110001;
      patterns[58282] = 29'b1_110001110101_010_1_100011101011;
      patterns[58283] = 29'b1_110001110101_011_1_000111010111;
      patterns[58284] = 29'b1_110001110101_100_1_111000111010;
      patterns[58285] = 29'b1_110001110101_101_0_111100011101;
      patterns[58286] = 29'b1_110001110101_110_1_110001110101;
      patterns[58287] = 29'b1_110001110101_111_1_110001110101;
      patterns[58288] = 29'b1_110001110110_000_1_110001110110;
      patterns[58289] = 29'b1_110001110110_001_1_110110110001;
      patterns[58290] = 29'b1_110001110110_010_1_100011101101;
      patterns[58291] = 29'b1_110001110110_011_1_000111011011;
      patterns[58292] = 29'b1_110001110110_100_0_111000111011;
      patterns[58293] = 29'b1_110001110110_101_1_011100011101;
      patterns[58294] = 29'b1_110001110110_110_1_110001110110;
      patterns[58295] = 29'b1_110001110110_111_1_110001110110;
      patterns[58296] = 29'b1_110001110111_000_1_110001110111;
      patterns[58297] = 29'b1_110001110111_001_1_110111110001;
      patterns[58298] = 29'b1_110001110111_010_1_100011101111;
      patterns[58299] = 29'b1_110001110111_011_1_000111011111;
      patterns[58300] = 29'b1_110001110111_100_1_111000111011;
      patterns[58301] = 29'b1_110001110111_101_1_111100011101;
      patterns[58302] = 29'b1_110001110111_110_1_110001110111;
      patterns[58303] = 29'b1_110001110111_111_1_110001110111;
      patterns[58304] = 29'b1_110001111000_000_1_110001111000;
      patterns[58305] = 29'b1_110001111000_001_1_111000110001;
      patterns[58306] = 29'b1_110001111000_010_1_100011110001;
      patterns[58307] = 29'b1_110001111000_011_1_000111100011;
      patterns[58308] = 29'b1_110001111000_100_0_111000111100;
      patterns[58309] = 29'b1_110001111000_101_0_011100011110;
      patterns[58310] = 29'b1_110001111000_110_1_110001111000;
      patterns[58311] = 29'b1_110001111000_111_1_110001111000;
      patterns[58312] = 29'b1_110001111001_000_1_110001111001;
      patterns[58313] = 29'b1_110001111001_001_1_111001110001;
      patterns[58314] = 29'b1_110001111001_010_1_100011110011;
      patterns[58315] = 29'b1_110001111001_011_1_000111100111;
      patterns[58316] = 29'b1_110001111001_100_1_111000111100;
      patterns[58317] = 29'b1_110001111001_101_0_111100011110;
      patterns[58318] = 29'b1_110001111001_110_1_110001111001;
      patterns[58319] = 29'b1_110001111001_111_1_110001111001;
      patterns[58320] = 29'b1_110001111010_000_1_110001111010;
      patterns[58321] = 29'b1_110001111010_001_1_111010110001;
      patterns[58322] = 29'b1_110001111010_010_1_100011110101;
      patterns[58323] = 29'b1_110001111010_011_1_000111101011;
      patterns[58324] = 29'b1_110001111010_100_0_111000111101;
      patterns[58325] = 29'b1_110001111010_101_1_011100011110;
      patterns[58326] = 29'b1_110001111010_110_1_110001111010;
      patterns[58327] = 29'b1_110001111010_111_1_110001111010;
      patterns[58328] = 29'b1_110001111011_000_1_110001111011;
      patterns[58329] = 29'b1_110001111011_001_1_111011110001;
      patterns[58330] = 29'b1_110001111011_010_1_100011110111;
      patterns[58331] = 29'b1_110001111011_011_1_000111101111;
      patterns[58332] = 29'b1_110001111011_100_1_111000111101;
      patterns[58333] = 29'b1_110001111011_101_1_111100011110;
      patterns[58334] = 29'b1_110001111011_110_1_110001111011;
      patterns[58335] = 29'b1_110001111011_111_1_110001111011;
      patterns[58336] = 29'b1_110001111100_000_1_110001111100;
      patterns[58337] = 29'b1_110001111100_001_1_111100110001;
      patterns[58338] = 29'b1_110001111100_010_1_100011111001;
      patterns[58339] = 29'b1_110001111100_011_1_000111110011;
      patterns[58340] = 29'b1_110001111100_100_0_111000111110;
      patterns[58341] = 29'b1_110001111100_101_0_011100011111;
      patterns[58342] = 29'b1_110001111100_110_1_110001111100;
      patterns[58343] = 29'b1_110001111100_111_1_110001111100;
      patterns[58344] = 29'b1_110001111101_000_1_110001111101;
      patterns[58345] = 29'b1_110001111101_001_1_111101110001;
      patterns[58346] = 29'b1_110001111101_010_1_100011111011;
      patterns[58347] = 29'b1_110001111101_011_1_000111110111;
      patterns[58348] = 29'b1_110001111101_100_1_111000111110;
      patterns[58349] = 29'b1_110001111101_101_0_111100011111;
      patterns[58350] = 29'b1_110001111101_110_1_110001111101;
      patterns[58351] = 29'b1_110001111101_111_1_110001111101;
      patterns[58352] = 29'b1_110001111110_000_1_110001111110;
      patterns[58353] = 29'b1_110001111110_001_1_111110110001;
      patterns[58354] = 29'b1_110001111110_010_1_100011111101;
      patterns[58355] = 29'b1_110001111110_011_1_000111111011;
      patterns[58356] = 29'b1_110001111110_100_0_111000111111;
      patterns[58357] = 29'b1_110001111110_101_1_011100011111;
      patterns[58358] = 29'b1_110001111110_110_1_110001111110;
      patterns[58359] = 29'b1_110001111110_111_1_110001111110;
      patterns[58360] = 29'b1_110001111111_000_1_110001111111;
      patterns[58361] = 29'b1_110001111111_001_1_111111110001;
      patterns[58362] = 29'b1_110001111111_010_1_100011111111;
      patterns[58363] = 29'b1_110001111111_011_1_000111111111;
      patterns[58364] = 29'b1_110001111111_100_1_111000111111;
      patterns[58365] = 29'b1_110001111111_101_1_111100011111;
      patterns[58366] = 29'b1_110001111111_110_1_110001111111;
      patterns[58367] = 29'b1_110001111111_111_1_110001111111;
      patterns[58368] = 29'b1_110010000000_000_1_110010000000;
      patterns[58369] = 29'b1_110010000000_001_1_000000110010;
      patterns[58370] = 29'b1_110010000000_010_1_100100000001;
      patterns[58371] = 29'b1_110010000000_011_1_001000000011;
      patterns[58372] = 29'b1_110010000000_100_0_111001000000;
      patterns[58373] = 29'b1_110010000000_101_0_011100100000;
      patterns[58374] = 29'b1_110010000000_110_1_110010000000;
      patterns[58375] = 29'b1_110010000000_111_1_110010000000;
      patterns[58376] = 29'b1_110010000001_000_1_110010000001;
      patterns[58377] = 29'b1_110010000001_001_1_000001110010;
      patterns[58378] = 29'b1_110010000001_010_1_100100000011;
      patterns[58379] = 29'b1_110010000001_011_1_001000000111;
      patterns[58380] = 29'b1_110010000001_100_1_111001000000;
      patterns[58381] = 29'b1_110010000001_101_0_111100100000;
      patterns[58382] = 29'b1_110010000001_110_1_110010000001;
      patterns[58383] = 29'b1_110010000001_111_1_110010000001;
      patterns[58384] = 29'b1_110010000010_000_1_110010000010;
      patterns[58385] = 29'b1_110010000010_001_1_000010110010;
      patterns[58386] = 29'b1_110010000010_010_1_100100000101;
      patterns[58387] = 29'b1_110010000010_011_1_001000001011;
      patterns[58388] = 29'b1_110010000010_100_0_111001000001;
      patterns[58389] = 29'b1_110010000010_101_1_011100100000;
      patterns[58390] = 29'b1_110010000010_110_1_110010000010;
      patterns[58391] = 29'b1_110010000010_111_1_110010000010;
      patterns[58392] = 29'b1_110010000011_000_1_110010000011;
      patterns[58393] = 29'b1_110010000011_001_1_000011110010;
      patterns[58394] = 29'b1_110010000011_010_1_100100000111;
      patterns[58395] = 29'b1_110010000011_011_1_001000001111;
      patterns[58396] = 29'b1_110010000011_100_1_111001000001;
      patterns[58397] = 29'b1_110010000011_101_1_111100100000;
      patterns[58398] = 29'b1_110010000011_110_1_110010000011;
      patterns[58399] = 29'b1_110010000011_111_1_110010000011;
      patterns[58400] = 29'b1_110010000100_000_1_110010000100;
      patterns[58401] = 29'b1_110010000100_001_1_000100110010;
      patterns[58402] = 29'b1_110010000100_010_1_100100001001;
      patterns[58403] = 29'b1_110010000100_011_1_001000010011;
      patterns[58404] = 29'b1_110010000100_100_0_111001000010;
      patterns[58405] = 29'b1_110010000100_101_0_011100100001;
      patterns[58406] = 29'b1_110010000100_110_1_110010000100;
      patterns[58407] = 29'b1_110010000100_111_1_110010000100;
      patterns[58408] = 29'b1_110010000101_000_1_110010000101;
      patterns[58409] = 29'b1_110010000101_001_1_000101110010;
      patterns[58410] = 29'b1_110010000101_010_1_100100001011;
      patterns[58411] = 29'b1_110010000101_011_1_001000010111;
      patterns[58412] = 29'b1_110010000101_100_1_111001000010;
      patterns[58413] = 29'b1_110010000101_101_0_111100100001;
      patterns[58414] = 29'b1_110010000101_110_1_110010000101;
      patterns[58415] = 29'b1_110010000101_111_1_110010000101;
      patterns[58416] = 29'b1_110010000110_000_1_110010000110;
      patterns[58417] = 29'b1_110010000110_001_1_000110110010;
      patterns[58418] = 29'b1_110010000110_010_1_100100001101;
      patterns[58419] = 29'b1_110010000110_011_1_001000011011;
      patterns[58420] = 29'b1_110010000110_100_0_111001000011;
      patterns[58421] = 29'b1_110010000110_101_1_011100100001;
      patterns[58422] = 29'b1_110010000110_110_1_110010000110;
      patterns[58423] = 29'b1_110010000110_111_1_110010000110;
      patterns[58424] = 29'b1_110010000111_000_1_110010000111;
      patterns[58425] = 29'b1_110010000111_001_1_000111110010;
      patterns[58426] = 29'b1_110010000111_010_1_100100001111;
      patterns[58427] = 29'b1_110010000111_011_1_001000011111;
      patterns[58428] = 29'b1_110010000111_100_1_111001000011;
      patterns[58429] = 29'b1_110010000111_101_1_111100100001;
      patterns[58430] = 29'b1_110010000111_110_1_110010000111;
      patterns[58431] = 29'b1_110010000111_111_1_110010000111;
      patterns[58432] = 29'b1_110010001000_000_1_110010001000;
      patterns[58433] = 29'b1_110010001000_001_1_001000110010;
      patterns[58434] = 29'b1_110010001000_010_1_100100010001;
      patterns[58435] = 29'b1_110010001000_011_1_001000100011;
      patterns[58436] = 29'b1_110010001000_100_0_111001000100;
      patterns[58437] = 29'b1_110010001000_101_0_011100100010;
      patterns[58438] = 29'b1_110010001000_110_1_110010001000;
      patterns[58439] = 29'b1_110010001000_111_1_110010001000;
      patterns[58440] = 29'b1_110010001001_000_1_110010001001;
      patterns[58441] = 29'b1_110010001001_001_1_001001110010;
      patterns[58442] = 29'b1_110010001001_010_1_100100010011;
      patterns[58443] = 29'b1_110010001001_011_1_001000100111;
      patterns[58444] = 29'b1_110010001001_100_1_111001000100;
      patterns[58445] = 29'b1_110010001001_101_0_111100100010;
      patterns[58446] = 29'b1_110010001001_110_1_110010001001;
      patterns[58447] = 29'b1_110010001001_111_1_110010001001;
      patterns[58448] = 29'b1_110010001010_000_1_110010001010;
      patterns[58449] = 29'b1_110010001010_001_1_001010110010;
      patterns[58450] = 29'b1_110010001010_010_1_100100010101;
      patterns[58451] = 29'b1_110010001010_011_1_001000101011;
      patterns[58452] = 29'b1_110010001010_100_0_111001000101;
      patterns[58453] = 29'b1_110010001010_101_1_011100100010;
      patterns[58454] = 29'b1_110010001010_110_1_110010001010;
      patterns[58455] = 29'b1_110010001010_111_1_110010001010;
      patterns[58456] = 29'b1_110010001011_000_1_110010001011;
      patterns[58457] = 29'b1_110010001011_001_1_001011110010;
      patterns[58458] = 29'b1_110010001011_010_1_100100010111;
      patterns[58459] = 29'b1_110010001011_011_1_001000101111;
      patterns[58460] = 29'b1_110010001011_100_1_111001000101;
      patterns[58461] = 29'b1_110010001011_101_1_111100100010;
      patterns[58462] = 29'b1_110010001011_110_1_110010001011;
      patterns[58463] = 29'b1_110010001011_111_1_110010001011;
      patterns[58464] = 29'b1_110010001100_000_1_110010001100;
      patterns[58465] = 29'b1_110010001100_001_1_001100110010;
      patterns[58466] = 29'b1_110010001100_010_1_100100011001;
      patterns[58467] = 29'b1_110010001100_011_1_001000110011;
      patterns[58468] = 29'b1_110010001100_100_0_111001000110;
      patterns[58469] = 29'b1_110010001100_101_0_011100100011;
      patterns[58470] = 29'b1_110010001100_110_1_110010001100;
      patterns[58471] = 29'b1_110010001100_111_1_110010001100;
      patterns[58472] = 29'b1_110010001101_000_1_110010001101;
      patterns[58473] = 29'b1_110010001101_001_1_001101110010;
      patterns[58474] = 29'b1_110010001101_010_1_100100011011;
      patterns[58475] = 29'b1_110010001101_011_1_001000110111;
      patterns[58476] = 29'b1_110010001101_100_1_111001000110;
      patterns[58477] = 29'b1_110010001101_101_0_111100100011;
      patterns[58478] = 29'b1_110010001101_110_1_110010001101;
      patterns[58479] = 29'b1_110010001101_111_1_110010001101;
      patterns[58480] = 29'b1_110010001110_000_1_110010001110;
      patterns[58481] = 29'b1_110010001110_001_1_001110110010;
      patterns[58482] = 29'b1_110010001110_010_1_100100011101;
      patterns[58483] = 29'b1_110010001110_011_1_001000111011;
      patterns[58484] = 29'b1_110010001110_100_0_111001000111;
      patterns[58485] = 29'b1_110010001110_101_1_011100100011;
      patterns[58486] = 29'b1_110010001110_110_1_110010001110;
      patterns[58487] = 29'b1_110010001110_111_1_110010001110;
      patterns[58488] = 29'b1_110010001111_000_1_110010001111;
      patterns[58489] = 29'b1_110010001111_001_1_001111110010;
      patterns[58490] = 29'b1_110010001111_010_1_100100011111;
      patterns[58491] = 29'b1_110010001111_011_1_001000111111;
      patterns[58492] = 29'b1_110010001111_100_1_111001000111;
      patterns[58493] = 29'b1_110010001111_101_1_111100100011;
      patterns[58494] = 29'b1_110010001111_110_1_110010001111;
      patterns[58495] = 29'b1_110010001111_111_1_110010001111;
      patterns[58496] = 29'b1_110010010000_000_1_110010010000;
      patterns[58497] = 29'b1_110010010000_001_1_010000110010;
      patterns[58498] = 29'b1_110010010000_010_1_100100100001;
      patterns[58499] = 29'b1_110010010000_011_1_001001000011;
      patterns[58500] = 29'b1_110010010000_100_0_111001001000;
      patterns[58501] = 29'b1_110010010000_101_0_011100100100;
      patterns[58502] = 29'b1_110010010000_110_1_110010010000;
      patterns[58503] = 29'b1_110010010000_111_1_110010010000;
      patterns[58504] = 29'b1_110010010001_000_1_110010010001;
      patterns[58505] = 29'b1_110010010001_001_1_010001110010;
      patterns[58506] = 29'b1_110010010001_010_1_100100100011;
      patterns[58507] = 29'b1_110010010001_011_1_001001000111;
      patterns[58508] = 29'b1_110010010001_100_1_111001001000;
      patterns[58509] = 29'b1_110010010001_101_0_111100100100;
      patterns[58510] = 29'b1_110010010001_110_1_110010010001;
      patterns[58511] = 29'b1_110010010001_111_1_110010010001;
      patterns[58512] = 29'b1_110010010010_000_1_110010010010;
      patterns[58513] = 29'b1_110010010010_001_1_010010110010;
      patterns[58514] = 29'b1_110010010010_010_1_100100100101;
      patterns[58515] = 29'b1_110010010010_011_1_001001001011;
      patterns[58516] = 29'b1_110010010010_100_0_111001001001;
      patterns[58517] = 29'b1_110010010010_101_1_011100100100;
      patterns[58518] = 29'b1_110010010010_110_1_110010010010;
      patterns[58519] = 29'b1_110010010010_111_1_110010010010;
      patterns[58520] = 29'b1_110010010011_000_1_110010010011;
      patterns[58521] = 29'b1_110010010011_001_1_010011110010;
      patterns[58522] = 29'b1_110010010011_010_1_100100100111;
      patterns[58523] = 29'b1_110010010011_011_1_001001001111;
      patterns[58524] = 29'b1_110010010011_100_1_111001001001;
      patterns[58525] = 29'b1_110010010011_101_1_111100100100;
      patterns[58526] = 29'b1_110010010011_110_1_110010010011;
      patterns[58527] = 29'b1_110010010011_111_1_110010010011;
      patterns[58528] = 29'b1_110010010100_000_1_110010010100;
      patterns[58529] = 29'b1_110010010100_001_1_010100110010;
      patterns[58530] = 29'b1_110010010100_010_1_100100101001;
      patterns[58531] = 29'b1_110010010100_011_1_001001010011;
      patterns[58532] = 29'b1_110010010100_100_0_111001001010;
      patterns[58533] = 29'b1_110010010100_101_0_011100100101;
      patterns[58534] = 29'b1_110010010100_110_1_110010010100;
      patterns[58535] = 29'b1_110010010100_111_1_110010010100;
      patterns[58536] = 29'b1_110010010101_000_1_110010010101;
      patterns[58537] = 29'b1_110010010101_001_1_010101110010;
      patterns[58538] = 29'b1_110010010101_010_1_100100101011;
      patterns[58539] = 29'b1_110010010101_011_1_001001010111;
      patterns[58540] = 29'b1_110010010101_100_1_111001001010;
      patterns[58541] = 29'b1_110010010101_101_0_111100100101;
      patterns[58542] = 29'b1_110010010101_110_1_110010010101;
      patterns[58543] = 29'b1_110010010101_111_1_110010010101;
      patterns[58544] = 29'b1_110010010110_000_1_110010010110;
      patterns[58545] = 29'b1_110010010110_001_1_010110110010;
      patterns[58546] = 29'b1_110010010110_010_1_100100101101;
      patterns[58547] = 29'b1_110010010110_011_1_001001011011;
      patterns[58548] = 29'b1_110010010110_100_0_111001001011;
      patterns[58549] = 29'b1_110010010110_101_1_011100100101;
      patterns[58550] = 29'b1_110010010110_110_1_110010010110;
      patterns[58551] = 29'b1_110010010110_111_1_110010010110;
      patterns[58552] = 29'b1_110010010111_000_1_110010010111;
      patterns[58553] = 29'b1_110010010111_001_1_010111110010;
      patterns[58554] = 29'b1_110010010111_010_1_100100101111;
      patterns[58555] = 29'b1_110010010111_011_1_001001011111;
      patterns[58556] = 29'b1_110010010111_100_1_111001001011;
      patterns[58557] = 29'b1_110010010111_101_1_111100100101;
      patterns[58558] = 29'b1_110010010111_110_1_110010010111;
      patterns[58559] = 29'b1_110010010111_111_1_110010010111;
      patterns[58560] = 29'b1_110010011000_000_1_110010011000;
      patterns[58561] = 29'b1_110010011000_001_1_011000110010;
      patterns[58562] = 29'b1_110010011000_010_1_100100110001;
      patterns[58563] = 29'b1_110010011000_011_1_001001100011;
      patterns[58564] = 29'b1_110010011000_100_0_111001001100;
      patterns[58565] = 29'b1_110010011000_101_0_011100100110;
      patterns[58566] = 29'b1_110010011000_110_1_110010011000;
      patterns[58567] = 29'b1_110010011000_111_1_110010011000;
      patterns[58568] = 29'b1_110010011001_000_1_110010011001;
      patterns[58569] = 29'b1_110010011001_001_1_011001110010;
      patterns[58570] = 29'b1_110010011001_010_1_100100110011;
      patterns[58571] = 29'b1_110010011001_011_1_001001100111;
      patterns[58572] = 29'b1_110010011001_100_1_111001001100;
      patterns[58573] = 29'b1_110010011001_101_0_111100100110;
      patterns[58574] = 29'b1_110010011001_110_1_110010011001;
      patterns[58575] = 29'b1_110010011001_111_1_110010011001;
      patterns[58576] = 29'b1_110010011010_000_1_110010011010;
      patterns[58577] = 29'b1_110010011010_001_1_011010110010;
      patterns[58578] = 29'b1_110010011010_010_1_100100110101;
      patterns[58579] = 29'b1_110010011010_011_1_001001101011;
      patterns[58580] = 29'b1_110010011010_100_0_111001001101;
      patterns[58581] = 29'b1_110010011010_101_1_011100100110;
      patterns[58582] = 29'b1_110010011010_110_1_110010011010;
      patterns[58583] = 29'b1_110010011010_111_1_110010011010;
      patterns[58584] = 29'b1_110010011011_000_1_110010011011;
      patterns[58585] = 29'b1_110010011011_001_1_011011110010;
      patterns[58586] = 29'b1_110010011011_010_1_100100110111;
      patterns[58587] = 29'b1_110010011011_011_1_001001101111;
      patterns[58588] = 29'b1_110010011011_100_1_111001001101;
      patterns[58589] = 29'b1_110010011011_101_1_111100100110;
      patterns[58590] = 29'b1_110010011011_110_1_110010011011;
      patterns[58591] = 29'b1_110010011011_111_1_110010011011;
      patterns[58592] = 29'b1_110010011100_000_1_110010011100;
      patterns[58593] = 29'b1_110010011100_001_1_011100110010;
      patterns[58594] = 29'b1_110010011100_010_1_100100111001;
      patterns[58595] = 29'b1_110010011100_011_1_001001110011;
      patterns[58596] = 29'b1_110010011100_100_0_111001001110;
      patterns[58597] = 29'b1_110010011100_101_0_011100100111;
      patterns[58598] = 29'b1_110010011100_110_1_110010011100;
      patterns[58599] = 29'b1_110010011100_111_1_110010011100;
      patterns[58600] = 29'b1_110010011101_000_1_110010011101;
      patterns[58601] = 29'b1_110010011101_001_1_011101110010;
      patterns[58602] = 29'b1_110010011101_010_1_100100111011;
      patterns[58603] = 29'b1_110010011101_011_1_001001110111;
      patterns[58604] = 29'b1_110010011101_100_1_111001001110;
      patterns[58605] = 29'b1_110010011101_101_0_111100100111;
      patterns[58606] = 29'b1_110010011101_110_1_110010011101;
      patterns[58607] = 29'b1_110010011101_111_1_110010011101;
      patterns[58608] = 29'b1_110010011110_000_1_110010011110;
      patterns[58609] = 29'b1_110010011110_001_1_011110110010;
      patterns[58610] = 29'b1_110010011110_010_1_100100111101;
      patterns[58611] = 29'b1_110010011110_011_1_001001111011;
      patterns[58612] = 29'b1_110010011110_100_0_111001001111;
      patterns[58613] = 29'b1_110010011110_101_1_011100100111;
      patterns[58614] = 29'b1_110010011110_110_1_110010011110;
      patterns[58615] = 29'b1_110010011110_111_1_110010011110;
      patterns[58616] = 29'b1_110010011111_000_1_110010011111;
      patterns[58617] = 29'b1_110010011111_001_1_011111110010;
      patterns[58618] = 29'b1_110010011111_010_1_100100111111;
      patterns[58619] = 29'b1_110010011111_011_1_001001111111;
      patterns[58620] = 29'b1_110010011111_100_1_111001001111;
      patterns[58621] = 29'b1_110010011111_101_1_111100100111;
      patterns[58622] = 29'b1_110010011111_110_1_110010011111;
      patterns[58623] = 29'b1_110010011111_111_1_110010011111;
      patterns[58624] = 29'b1_110010100000_000_1_110010100000;
      patterns[58625] = 29'b1_110010100000_001_1_100000110010;
      patterns[58626] = 29'b1_110010100000_010_1_100101000001;
      patterns[58627] = 29'b1_110010100000_011_1_001010000011;
      patterns[58628] = 29'b1_110010100000_100_0_111001010000;
      patterns[58629] = 29'b1_110010100000_101_0_011100101000;
      patterns[58630] = 29'b1_110010100000_110_1_110010100000;
      patterns[58631] = 29'b1_110010100000_111_1_110010100000;
      patterns[58632] = 29'b1_110010100001_000_1_110010100001;
      patterns[58633] = 29'b1_110010100001_001_1_100001110010;
      patterns[58634] = 29'b1_110010100001_010_1_100101000011;
      patterns[58635] = 29'b1_110010100001_011_1_001010000111;
      patterns[58636] = 29'b1_110010100001_100_1_111001010000;
      patterns[58637] = 29'b1_110010100001_101_0_111100101000;
      patterns[58638] = 29'b1_110010100001_110_1_110010100001;
      patterns[58639] = 29'b1_110010100001_111_1_110010100001;
      patterns[58640] = 29'b1_110010100010_000_1_110010100010;
      patterns[58641] = 29'b1_110010100010_001_1_100010110010;
      patterns[58642] = 29'b1_110010100010_010_1_100101000101;
      patterns[58643] = 29'b1_110010100010_011_1_001010001011;
      patterns[58644] = 29'b1_110010100010_100_0_111001010001;
      patterns[58645] = 29'b1_110010100010_101_1_011100101000;
      patterns[58646] = 29'b1_110010100010_110_1_110010100010;
      patterns[58647] = 29'b1_110010100010_111_1_110010100010;
      patterns[58648] = 29'b1_110010100011_000_1_110010100011;
      patterns[58649] = 29'b1_110010100011_001_1_100011110010;
      patterns[58650] = 29'b1_110010100011_010_1_100101000111;
      patterns[58651] = 29'b1_110010100011_011_1_001010001111;
      patterns[58652] = 29'b1_110010100011_100_1_111001010001;
      patterns[58653] = 29'b1_110010100011_101_1_111100101000;
      patterns[58654] = 29'b1_110010100011_110_1_110010100011;
      patterns[58655] = 29'b1_110010100011_111_1_110010100011;
      patterns[58656] = 29'b1_110010100100_000_1_110010100100;
      patterns[58657] = 29'b1_110010100100_001_1_100100110010;
      patterns[58658] = 29'b1_110010100100_010_1_100101001001;
      patterns[58659] = 29'b1_110010100100_011_1_001010010011;
      patterns[58660] = 29'b1_110010100100_100_0_111001010010;
      patterns[58661] = 29'b1_110010100100_101_0_011100101001;
      patterns[58662] = 29'b1_110010100100_110_1_110010100100;
      patterns[58663] = 29'b1_110010100100_111_1_110010100100;
      patterns[58664] = 29'b1_110010100101_000_1_110010100101;
      patterns[58665] = 29'b1_110010100101_001_1_100101110010;
      patterns[58666] = 29'b1_110010100101_010_1_100101001011;
      patterns[58667] = 29'b1_110010100101_011_1_001010010111;
      patterns[58668] = 29'b1_110010100101_100_1_111001010010;
      patterns[58669] = 29'b1_110010100101_101_0_111100101001;
      patterns[58670] = 29'b1_110010100101_110_1_110010100101;
      patterns[58671] = 29'b1_110010100101_111_1_110010100101;
      patterns[58672] = 29'b1_110010100110_000_1_110010100110;
      patterns[58673] = 29'b1_110010100110_001_1_100110110010;
      patterns[58674] = 29'b1_110010100110_010_1_100101001101;
      patterns[58675] = 29'b1_110010100110_011_1_001010011011;
      patterns[58676] = 29'b1_110010100110_100_0_111001010011;
      patterns[58677] = 29'b1_110010100110_101_1_011100101001;
      patterns[58678] = 29'b1_110010100110_110_1_110010100110;
      patterns[58679] = 29'b1_110010100110_111_1_110010100110;
      patterns[58680] = 29'b1_110010100111_000_1_110010100111;
      patterns[58681] = 29'b1_110010100111_001_1_100111110010;
      patterns[58682] = 29'b1_110010100111_010_1_100101001111;
      patterns[58683] = 29'b1_110010100111_011_1_001010011111;
      patterns[58684] = 29'b1_110010100111_100_1_111001010011;
      patterns[58685] = 29'b1_110010100111_101_1_111100101001;
      patterns[58686] = 29'b1_110010100111_110_1_110010100111;
      patterns[58687] = 29'b1_110010100111_111_1_110010100111;
      patterns[58688] = 29'b1_110010101000_000_1_110010101000;
      patterns[58689] = 29'b1_110010101000_001_1_101000110010;
      patterns[58690] = 29'b1_110010101000_010_1_100101010001;
      patterns[58691] = 29'b1_110010101000_011_1_001010100011;
      patterns[58692] = 29'b1_110010101000_100_0_111001010100;
      patterns[58693] = 29'b1_110010101000_101_0_011100101010;
      patterns[58694] = 29'b1_110010101000_110_1_110010101000;
      patterns[58695] = 29'b1_110010101000_111_1_110010101000;
      patterns[58696] = 29'b1_110010101001_000_1_110010101001;
      patterns[58697] = 29'b1_110010101001_001_1_101001110010;
      patterns[58698] = 29'b1_110010101001_010_1_100101010011;
      patterns[58699] = 29'b1_110010101001_011_1_001010100111;
      patterns[58700] = 29'b1_110010101001_100_1_111001010100;
      patterns[58701] = 29'b1_110010101001_101_0_111100101010;
      patterns[58702] = 29'b1_110010101001_110_1_110010101001;
      patterns[58703] = 29'b1_110010101001_111_1_110010101001;
      patterns[58704] = 29'b1_110010101010_000_1_110010101010;
      patterns[58705] = 29'b1_110010101010_001_1_101010110010;
      patterns[58706] = 29'b1_110010101010_010_1_100101010101;
      patterns[58707] = 29'b1_110010101010_011_1_001010101011;
      patterns[58708] = 29'b1_110010101010_100_0_111001010101;
      patterns[58709] = 29'b1_110010101010_101_1_011100101010;
      patterns[58710] = 29'b1_110010101010_110_1_110010101010;
      patterns[58711] = 29'b1_110010101010_111_1_110010101010;
      patterns[58712] = 29'b1_110010101011_000_1_110010101011;
      patterns[58713] = 29'b1_110010101011_001_1_101011110010;
      patterns[58714] = 29'b1_110010101011_010_1_100101010111;
      patterns[58715] = 29'b1_110010101011_011_1_001010101111;
      patterns[58716] = 29'b1_110010101011_100_1_111001010101;
      patterns[58717] = 29'b1_110010101011_101_1_111100101010;
      patterns[58718] = 29'b1_110010101011_110_1_110010101011;
      patterns[58719] = 29'b1_110010101011_111_1_110010101011;
      patterns[58720] = 29'b1_110010101100_000_1_110010101100;
      patterns[58721] = 29'b1_110010101100_001_1_101100110010;
      patterns[58722] = 29'b1_110010101100_010_1_100101011001;
      patterns[58723] = 29'b1_110010101100_011_1_001010110011;
      patterns[58724] = 29'b1_110010101100_100_0_111001010110;
      patterns[58725] = 29'b1_110010101100_101_0_011100101011;
      patterns[58726] = 29'b1_110010101100_110_1_110010101100;
      patterns[58727] = 29'b1_110010101100_111_1_110010101100;
      patterns[58728] = 29'b1_110010101101_000_1_110010101101;
      patterns[58729] = 29'b1_110010101101_001_1_101101110010;
      patterns[58730] = 29'b1_110010101101_010_1_100101011011;
      patterns[58731] = 29'b1_110010101101_011_1_001010110111;
      patterns[58732] = 29'b1_110010101101_100_1_111001010110;
      patterns[58733] = 29'b1_110010101101_101_0_111100101011;
      patterns[58734] = 29'b1_110010101101_110_1_110010101101;
      patterns[58735] = 29'b1_110010101101_111_1_110010101101;
      patterns[58736] = 29'b1_110010101110_000_1_110010101110;
      patterns[58737] = 29'b1_110010101110_001_1_101110110010;
      patterns[58738] = 29'b1_110010101110_010_1_100101011101;
      patterns[58739] = 29'b1_110010101110_011_1_001010111011;
      patterns[58740] = 29'b1_110010101110_100_0_111001010111;
      patterns[58741] = 29'b1_110010101110_101_1_011100101011;
      patterns[58742] = 29'b1_110010101110_110_1_110010101110;
      patterns[58743] = 29'b1_110010101110_111_1_110010101110;
      patterns[58744] = 29'b1_110010101111_000_1_110010101111;
      patterns[58745] = 29'b1_110010101111_001_1_101111110010;
      patterns[58746] = 29'b1_110010101111_010_1_100101011111;
      patterns[58747] = 29'b1_110010101111_011_1_001010111111;
      patterns[58748] = 29'b1_110010101111_100_1_111001010111;
      patterns[58749] = 29'b1_110010101111_101_1_111100101011;
      patterns[58750] = 29'b1_110010101111_110_1_110010101111;
      patterns[58751] = 29'b1_110010101111_111_1_110010101111;
      patterns[58752] = 29'b1_110010110000_000_1_110010110000;
      patterns[58753] = 29'b1_110010110000_001_1_110000110010;
      patterns[58754] = 29'b1_110010110000_010_1_100101100001;
      patterns[58755] = 29'b1_110010110000_011_1_001011000011;
      patterns[58756] = 29'b1_110010110000_100_0_111001011000;
      patterns[58757] = 29'b1_110010110000_101_0_011100101100;
      patterns[58758] = 29'b1_110010110000_110_1_110010110000;
      patterns[58759] = 29'b1_110010110000_111_1_110010110000;
      patterns[58760] = 29'b1_110010110001_000_1_110010110001;
      patterns[58761] = 29'b1_110010110001_001_1_110001110010;
      patterns[58762] = 29'b1_110010110001_010_1_100101100011;
      patterns[58763] = 29'b1_110010110001_011_1_001011000111;
      patterns[58764] = 29'b1_110010110001_100_1_111001011000;
      patterns[58765] = 29'b1_110010110001_101_0_111100101100;
      patterns[58766] = 29'b1_110010110001_110_1_110010110001;
      patterns[58767] = 29'b1_110010110001_111_1_110010110001;
      patterns[58768] = 29'b1_110010110010_000_1_110010110010;
      patterns[58769] = 29'b1_110010110010_001_1_110010110010;
      patterns[58770] = 29'b1_110010110010_010_1_100101100101;
      patterns[58771] = 29'b1_110010110010_011_1_001011001011;
      patterns[58772] = 29'b1_110010110010_100_0_111001011001;
      patterns[58773] = 29'b1_110010110010_101_1_011100101100;
      patterns[58774] = 29'b1_110010110010_110_1_110010110010;
      patterns[58775] = 29'b1_110010110010_111_1_110010110010;
      patterns[58776] = 29'b1_110010110011_000_1_110010110011;
      patterns[58777] = 29'b1_110010110011_001_1_110011110010;
      patterns[58778] = 29'b1_110010110011_010_1_100101100111;
      patterns[58779] = 29'b1_110010110011_011_1_001011001111;
      patterns[58780] = 29'b1_110010110011_100_1_111001011001;
      patterns[58781] = 29'b1_110010110011_101_1_111100101100;
      patterns[58782] = 29'b1_110010110011_110_1_110010110011;
      patterns[58783] = 29'b1_110010110011_111_1_110010110011;
      patterns[58784] = 29'b1_110010110100_000_1_110010110100;
      patterns[58785] = 29'b1_110010110100_001_1_110100110010;
      patterns[58786] = 29'b1_110010110100_010_1_100101101001;
      patterns[58787] = 29'b1_110010110100_011_1_001011010011;
      patterns[58788] = 29'b1_110010110100_100_0_111001011010;
      patterns[58789] = 29'b1_110010110100_101_0_011100101101;
      patterns[58790] = 29'b1_110010110100_110_1_110010110100;
      patterns[58791] = 29'b1_110010110100_111_1_110010110100;
      patterns[58792] = 29'b1_110010110101_000_1_110010110101;
      patterns[58793] = 29'b1_110010110101_001_1_110101110010;
      patterns[58794] = 29'b1_110010110101_010_1_100101101011;
      patterns[58795] = 29'b1_110010110101_011_1_001011010111;
      patterns[58796] = 29'b1_110010110101_100_1_111001011010;
      patterns[58797] = 29'b1_110010110101_101_0_111100101101;
      patterns[58798] = 29'b1_110010110101_110_1_110010110101;
      patterns[58799] = 29'b1_110010110101_111_1_110010110101;
      patterns[58800] = 29'b1_110010110110_000_1_110010110110;
      patterns[58801] = 29'b1_110010110110_001_1_110110110010;
      patterns[58802] = 29'b1_110010110110_010_1_100101101101;
      patterns[58803] = 29'b1_110010110110_011_1_001011011011;
      patterns[58804] = 29'b1_110010110110_100_0_111001011011;
      patterns[58805] = 29'b1_110010110110_101_1_011100101101;
      patterns[58806] = 29'b1_110010110110_110_1_110010110110;
      patterns[58807] = 29'b1_110010110110_111_1_110010110110;
      patterns[58808] = 29'b1_110010110111_000_1_110010110111;
      patterns[58809] = 29'b1_110010110111_001_1_110111110010;
      patterns[58810] = 29'b1_110010110111_010_1_100101101111;
      patterns[58811] = 29'b1_110010110111_011_1_001011011111;
      patterns[58812] = 29'b1_110010110111_100_1_111001011011;
      patterns[58813] = 29'b1_110010110111_101_1_111100101101;
      patterns[58814] = 29'b1_110010110111_110_1_110010110111;
      patterns[58815] = 29'b1_110010110111_111_1_110010110111;
      patterns[58816] = 29'b1_110010111000_000_1_110010111000;
      patterns[58817] = 29'b1_110010111000_001_1_111000110010;
      patterns[58818] = 29'b1_110010111000_010_1_100101110001;
      patterns[58819] = 29'b1_110010111000_011_1_001011100011;
      patterns[58820] = 29'b1_110010111000_100_0_111001011100;
      patterns[58821] = 29'b1_110010111000_101_0_011100101110;
      patterns[58822] = 29'b1_110010111000_110_1_110010111000;
      patterns[58823] = 29'b1_110010111000_111_1_110010111000;
      patterns[58824] = 29'b1_110010111001_000_1_110010111001;
      patterns[58825] = 29'b1_110010111001_001_1_111001110010;
      patterns[58826] = 29'b1_110010111001_010_1_100101110011;
      patterns[58827] = 29'b1_110010111001_011_1_001011100111;
      patterns[58828] = 29'b1_110010111001_100_1_111001011100;
      patterns[58829] = 29'b1_110010111001_101_0_111100101110;
      patterns[58830] = 29'b1_110010111001_110_1_110010111001;
      patterns[58831] = 29'b1_110010111001_111_1_110010111001;
      patterns[58832] = 29'b1_110010111010_000_1_110010111010;
      patterns[58833] = 29'b1_110010111010_001_1_111010110010;
      patterns[58834] = 29'b1_110010111010_010_1_100101110101;
      patterns[58835] = 29'b1_110010111010_011_1_001011101011;
      patterns[58836] = 29'b1_110010111010_100_0_111001011101;
      patterns[58837] = 29'b1_110010111010_101_1_011100101110;
      patterns[58838] = 29'b1_110010111010_110_1_110010111010;
      patterns[58839] = 29'b1_110010111010_111_1_110010111010;
      patterns[58840] = 29'b1_110010111011_000_1_110010111011;
      patterns[58841] = 29'b1_110010111011_001_1_111011110010;
      patterns[58842] = 29'b1_110010111011_010_1_100101110111;
      patterns[58843] = 29'b1_110010111011_011_1_001011101111;
      patterns[58844] = 29'b1_110010111011_100_1_111001011101;
      patterns[58845] = 29'b1_110010111011_101_1_111100101110;
      patterns[58846] = 29'b1_110010111011_110_1_110010111011;
      patterns[58847] = 29'b1_110010111011_111_1_110010111011;
      patterns[58848] = 29'b1_110010111100_000_1_110010111100;
      patterns[58849] = 29'b1_110010111100_001_1_111100110010;
      patterns[58850] = 29'b1_110010111100_010_1_100101111001;
      patterns[58851] = 29'b1_110010111100_011_1_001011110011;
      patterns[58852] = 29'b1_110010111100_100_0_111001011110;
      patterns[58853] = 29'b1_110010111100_101_0_011100101111;
      patterns[58854] = 29'b1_110010111100_110_1_110010111100;
      patterns[58855] = 29'b1_110010111100_111_1_110010111100;
      patterns[58856] = 29'b1_110010111101_000_1_110010111101;
      patterns[58857] = 29'b1_110010111101_001_1_111101110010;
      patterns[58858] = 29'b1_110010111101_010_1_100101111011;
      patterns[58859] = 29'b1_110010111101_011_1_001011110111;
      patterns[58860] = 29'b1_110010111101_100_1_111001011110;
      patterns[58861] = 29'b1_110010111101_101_0_111100101111;
      patterns[58862] = 29'b1_110010111101_110_1_110010111101;
      patterns[58863] = 29'b1_110010111101_111_1_110010111101;
      patterns[58864] = 29'b1_110010111110_000_1_110010111110;
      patterns[58865] = 29'b1_110010111110_001_1_111110110010;
      patterns[58866] = 29'b1_110010111110_010_1_100101111101;
      patterns[58867] = 29'b1_110010111110_011_1_001011111011;
      patterns[58868] = 29'b1_110010111110_100_0_111001011111;
      patterns[58869] = 29'b1_110010111110_101_1_011100101111;
      patterns[58870] = 29'b1_110010111110_110_1_110010111110;
      patterns[58871] = 29'b1_110010111110_111_1_110010111110;
      patterns[58872] = 29'b1_110010111111_000_1_110010111111;
      patterns[58873] = 29'b1_110010111111_001_1_111111110010;
      patterns[58874] = 29'b1_110010111111_010_1_100101111111;
      patterns[58875] = 29'b1_110010111111_011_1_001011111111;
      patterns[58876] = 29'b1_110010111111_100_1_111001011111;
      patterns[58877] = 29'b1_110010111111_101_1_111100101111;
      patterns[58878] = 29'b1_110010111111_110_1_110010111111;
      patterns[58879] = 29'b1_110010111111_111_1_110010111111;
      patterns[58880] = 29'b1_110011000000_000_1_110011000000;
      patterns[58881] = 29'b1_110011000000_001_1_000000110011;
      patterns[58882] = 29'b1_110011000000_010_1_100110000001;
      patterns[58883] = 29'b1_110011000000_011_1_001100000011;
      patterns[58884] = 29'b1_110011000000_100_0_111001100000;
      patterns[58885] = 29'b1_110011000000_101_0_011100110000;
      patterns[58886] = 29'b1_110011000000_110_1_110011000000;
      patterns[58887] = 29'b1_110011000000_111_1_110011000000;
      patterns[58888] = 29'b1_110011000001_000_1_110011000001;
      patterns[58889] = 29'b1_110011000001_001_1_000001110011;
      patterns[58890] = 29'b1_110011000001_010_1_100110000011;
      patterns[58891] = 29'b1_110011000001_011_1_001100000111;
      patterns[58892] = 29'b1_110011000001_100_1_111001100000;
      patterns[58893] = 29'b1_110011000001_101_0_111100110000;
      patterns[58894] = 29'b1_110011000001_110_1_110011000001;
      patterns[58895] = 29'b1_110011000001_111_1_110011000001;
      patterns[58896] = 29'b1_110011000010_000_1_110011000010;
      patterns[58897] = 29'b1_110011000010_001_1_000010110011;
      patterns[58898] = 29'b1_110011000010_010_1_100110000101;
      patterns[58899] = 29'b1_110011000010_011_1_001100001011;
      patterns[58900] = 29'b1_110011000010_100_0_111001100001;
      patterns[58901] = 29'b1_110011000010_101_1_011100110000;
      patterns[58902] = 29'b1_110011000010_110_1_110011000010;
      patterns[58903] = 29'b1_110011000010_111_1_110011000010;
      patterns[58904] = 29'b1_110011000011_000_1_110011000011;
      patterns[58905] = 29'b1_110011000011_001_1_000011110011;
      patterns[58906] = 29'b1_110011000011_010_1_100110000111;
      patterns[58907] = 29'b1_110011000011_011_1_001100001111;
      patterns[58908] = 29'b1_110011000011_100_1_111001100001;
      patterns[58909] = 29'b1_110011000011_101_1_111100110000;
      patterns[58910] = 29'b1_110011000011_110_1_110011000011;
      patterns[58911] = 29'b1_110011000011_111_1_110011000011;
      patterns[58912] = 29'b1_110011000100_000_1_110011000100;
      patterns[58913] = 29'b1_110011000100_001_1_000100110011;
      patterns[58914] = 29'b1_110011000100_010_1_100110001001;
      patterns[58915] = 29'b1_110011000100_011_1_001100010011;
      patterns[58916] = 29'b1_110011000100_100_0_111001100010;
      patterns[58917] = 29'b1_110011000100_101_0_011100110001;
      patterns[58918] = 29'b1_110011000100_110_1_110011000100;
      patterns[58919] = 29'b1_110011000100_111_1_110011000100;
      patterns[58920] = 29'b1_110011000101_000_1_110011000101;
      patterns[58921] = 29'b1_110011000101_001_1_000101110011;
      patterns[58922] = 29'b1_110011000101_010_1_100110001011;
      patterns[58923] = 29'b1_110011000101_011_1_001100010111;
      patterns[58924] = 29'b1_110011000101_100_1_111001100010;
      patterns[58925] = 29'b1_110011000101_101_0_111100110001;
      patterns[58926] = 29'b1_110011000101_110_1_110011000101;
      patterns[58927] = 29'b1_110011000101_111_1_110011000101;
      patterns[58928] = 29'b1_110011000110_000_1_110011000110;
      patterns[58929] = 29'b1_110011000110_001_1_000110110011;
      patterns[58930] = 29'b1_110011000110_010_1_100110001101;
      patterns[58931] = 29'b1_110011000110_011_1_001100011011;
      patterns[58932] = 29'b1_110011000110_100_0_111001100011;
      patterns[58933] = 29'b1_110011000110_101_1_011100110001;
      patterns[58934] = 29'b1_110011000110_110_1_110011000110;
      patterns[58935] = 29'b1_110011000110_111_1_110011000110;
      patterns[58936] = 29'b1_110011000111_000_1_110011000111;
      patterns[58937] = 29'b1_110011000111_001_1_000111110011;
      patterns[58938] = 29'b1_110011000111_010_1_100110001111;
      patterns[58939] = 29'b1_110011000111_011_1_001100011111;
      patterns[58940] = 29'b1_110011000111_100_1_111001100011;
      patterns[58941] = 29'b1_110011000111_101_1_111100110001;
      patterns[58942] = 29'b1_110011000111_110_1_110011000111;
      patterns[58943] = 29'b1_110011000111_111_1_110011000111;
      patterns[58944] = 29'b1_110011001000_000_1_110011001000;
      patterns[58945] = 29'b1_110011001000_001_1_001000110011;
      patterns[58946] = 29'b1_110011001000_010_1_100110010001;
      patterns[58947] = 29'b1_110011001000_011_1_001100100011;
      patterns[58948] = 29'b1_110011001000_100_0_111001100100;
      patterns[58949] = 29'b1_110011001000_101_0_011100110010;
      patterns[58950] = 29'b1_110011001000_110_1_110011001000;
      patterns[58951] = 29'b1_110011001000_111_1_110011001000;
      patterns[58952] = 29'b1_110011001001_000_1_110011001001;
      patterns[58953] = 29'b1_110011001001_001_1_001001110011;
      patterns[58954] = 29'b1_110011001001_010_1_100110010011;
      patterns[58955] = 29'b1_110011001001_011_1_001100100111;
      patterns[58956] = 29'b1_110011001001_100_1_111001100100;
      patterns[58957] = 29'b1_110011001001_101_0_111100110010;
      patterns[58958] = 29'b1_110011001001_110_1_110011001001;
      patterns[58959] = 29'b1_110011001001_111_1_110011001001;
      patterns[58960] = 29'b1_110011001010_000_1_110011001010;
      patterns[58961] = 29'b1_110011001010_001_1_001010110011;
      patterns[58962] = 29'b1_110011001010_010_1_100110010101;
      patterns[58963] = 29'b1_110011001010_011_1_001100101011;
      patterns[58964] = 29'b1_110011001010_100_0_111001100101;
      patterns[58965] = 29'b1_110011001010_101_1_011100110010;
      patterns[58966] = 29'b1_110011001010_110_1_110011001010;
      patterns[58967] = 29'b1_110011001010_111_1_110011001010;
      patterns[58968] = 29'b1_110011001011_000_1_110011001011;
      patterns[58969] = 29'b1_110011001011_001_1_001011110011;
      patterns[58970] = 29'b1_110011001011_010_1_100110010111;
      patterns[58971] = 29'b1_110011001011_011_1_001100101111;
      patterns[58972] = 29'b1_110011001011_100_1_111001100101;
      patterns[58973] = 29'b1_110011001011_101_1_111100110010;
      patterns[58974] = 29'b1_110011001011_110_1_110011001011;
      patterns[58975] = 29'b1_110011001011_111_1_110011001011;
      patterns[58976] = 29'b1_110011001100_000_1_110011001100;
      patterns[58977] = 29'b1_110011001100_001_1_001100110011;
      patterns[58978] = 29'b1_110011001100_010_1_100110011001;
      patterns[58979] = 29'b1_110011001100_011_1_001100110011;
      patterns[58980] = 29'b1_110011001100_100_0_111001100110;
      patterns[58981] = 29'b1_110011001100_101_0_011100110011;
      patterns[58982] = 29'b1_110011001100_110_1_110011001100;
      patterns[58983] = 29'b1_110011001100_111_1_110011001100;
      patterns[58984] = 29'b1_110011001101_000_1_110011001101;
      patterns[58985] = 29'b1_110011001101_001_1_001101110011;
      patterns[58986] = 29'b1_110011001101_010_1_100110011011;
      patterns[58987] = 29'b1_110011001101_011_1_001100110111;
      patterns[58988] = 29'b1_110011001101_100_1_111001100110;
      patterns[58989] = 29'b1_110011001101_101_0_111100110011;
      patterns[58990] = 29'b1_110011001101_110_1_110011001101;
      patterns[58991] = 29'b1_110011001101_111_1_110011001101;
      patterns[58992] = 29'b1_110011001110_000_1_110011001110;
      patterns[58993] = 29'b1_110011001110_001_1_001110110011;
      patterns[58994] = 29'b1_110011001110_010_1_100110011101;
      patterns[58995] = 29'b1_110011001110_011_1_001100111011;
      patterns[58996] = 29'b1_110011001110_100_0_111001100111;
      patterns[58997] = 29'b1_110011001110_101_1_011100110011;
      patterns[58998] = 29'b1_110011001110_110_1_110011001110;
      patterns[58999] = 29'b1_110011001110_111_1_110011001110;
      patterns[59000] = 29'b1_110011001111_000_1_110011001111;
      patterns[59001] = 29'b1_110011001111_001_1_001111110011;
      patterns[59002] = 29'b1_110011001111_010_1_100110011111;
      patterns[59003] = 29'b1_110011001111_011_1_001100111111;
      patterns[59004] = 29'b1_110011001111_100_1_111001100111;
      patterns[59005] = 29'b1_110011001111_101_1_111100110011;
      patterns[59006] = 29'b1_110011001111_110_1_110011001111;
      patterns[59007] = 29'b1_110011001111_111_1_110011001111;
      patterns[59008] = 29'b1_110011010000_000_1_110011010000;
      patterns[59009] = 29'b1_110011010000_001_1_010000110011;
      patterns[59010] = 29'b1_110011010000_010_1_100110100001;
      patterns[59011] = 29'b1_110011010000_011_1_001101000011;
      patterns[59012] = 29'b1_110011010000_100_0_111001101000;
      patterns[59013] = 29'b1_110011010000_101_0_011100110100;
      patterns[59014] = 29'b1_110011010000_110_1_110011010000;
      patterns[59015] = 29'b1_110011010000_111_1_110011010000;
      patterns[59016] = 29'b1_110011010001_000_1_110011010001;
      patterns[59017] = 29'b1_110011010001_001_1_010001110011;
      patterns[59018] = 29'b1_110011010001_010_1_100110100011;
      patterns[59019] = 29'b1_110011010001_011_1_001101000111;
      patterns[59020] = 29'b1_110011010001_100_1_111001101000;
      patterns[59021] = 29'b1_110011010001_101_0_111100110100;
      patterns[59022] = 29'b1_110011010001_110_1_110011010001;
      patterns[59023] = 29'b1_110011010001_111_1_110011010001;
      patterns[59024] = 29'b1_110011010010_000_1_110011010010;
      patterns[59025] = 29'b1_110011010010_001_1_010010110011;
      patterns[59026] = 29'b1_110011010010_010_1_100110100101;
      patterns[59027] = 29'b1_110011010010_011_1_001101001011;
      patterns[59028] = 29'b1_110011010010_100_0_111001101001;
      patterns[59029] = 29'b1_110011010010_101_1_011100110100;
      patterns[59030] = 29'b1_110011010010_110_1_110011010010;
      patterns[59031] = 29'b1_110011010010_111_1_110011010010;
      patterns[59032] = 29'b1_110011010011_000_1_110011010011;
      patterns[59033] = 29'b1_110011010011_001_1_010011110011;
      patterns[59034] = 29'b1_110011010011_010_1_100110100111;
      patterns[59035] = 29'b1_110011010011_011_1_001101001111;
      patterns[59036] = 29'b1_110011010011_100_1_111001101001;
      patterns[59037] = 29'b1_110011010011_101_1_111100110100;
      patterns[59038] = 29'b1_110011010011_110_1_110011010011;
      patterns[59039] = 29'b1_110011010011_111_1_110011010011;
      patterns[59040] = 29'b1_110011010100_000_1_110011010100;
      patterns[59041] = 29'b1_110011010100_001_1_010100110011;
      patterns[59042] = 29'b1_110011010100_010_1_100110101001;
      patterns[59043] = 29'b1_110011010100_011_1_001101010011;
      patterns[59044] = 29'b1_110011010100_100_0_111001101010;
      patterns[59045] = 29'b1_110011010100_101_0_011100110101;
      patterns[59046] = 29'b1_110011010100_110_1_110011010100;
      patterns[59047] = 29'b1_110011010100_111_1_110011010100;
      patterns[59048] = 29'b1_110011010101_000_1_110011010101;
      patterns[59049] = 29'b1_110011010101_001_1_010101110011;
      patterns[59050] = 29'b1_110011010101_010_1_100110101011;
      patterns[59051] = 29'b1_110011010101_011_1_001101010111;
      patterns[59052] = 29'b1_110011010101_100_1_111001101010;
      patterns[59053] = 29'b1_110011010101_101_0_111100110101;
      patterns[59054] = 29'b1_110011010101_110_1_110011010101;
      patterns[59055] = 29'b1_110011010101_111_1_110011010101;
      patterns[59056] = 29'b1_110011010110_000_1_110011010110;
      patterns[59057] = 29'b1_110011010110_001_1_010110110011;
      patterns[59058] = 29'b1_110011010110_010_1_100110101101;
      patterns[59059] = 29'b1_110011010110_011_1_001101011011;
      patterns[59060] = 29'b1_110011010110_100_0_111001101011;
      patterns[59061] = 29'b1_110011010110_101_1_011100110101;
      patterns[59062] = 29'b1_110011010110_110_1_110011010110;
      patterns[59063] = 29'b1_110011010110_111_1_110011010110;
      patterns[59064] = 29'b1_110011010111_000_1_110011010111;
      patterns[59065] = 29'b1_110011010111_001_1_010111110011;
      patterns[59066] = 29'b1_110011010111_010_1_100110101111;
      patterns[59067] = 29'b1_110011010111_011_1_001101011111;
      patterns[59068] = 29'b1_110011010111_100_1_111001101011;
      patterns[59069] = 29'b1_110011010111_101_1_111100110101;
      patterns[59070] = 29'b1_110011010111_110_1_110011010111;
      patterns[59071] = 29'b1_110011010111_111_1_110011010111;
      patterns[59072] = 29'b1_110011011000_000_1_110011011000;
      patterns[59073] = 29'b1_110011011000_001_1_011000110011;
      patterns[59074] = 29'b1_110011011000_010_1_100110110001;
      patterns[59075] = 29'b1_110011011000_011_1_001101100011;
      patterns[59076] = 29'b1_110011011000_100_0_111001101100;
      patterns[59077] = 29'b1_110011011000_101_0_011100110110;
      patterns[59078] = 29'b1_110011011000_110_1_110011011000;
      patterns[59079] = 29'b1_110011011000_111_1_110011011000;
      patterns[59080] = 29'b1_110011011001_000_1_110011011001;
      patterns[59081] = 29'b1_110011011001_001_1_011001110011;
      patterns[59082] = 29'b1_110011011001_010_1_100110110011;
      patterns[59083] = 29'b1_110011011001_011_1_001101100111;
      patterns[59084] = 29'b1_110011011001_100_1_111001101100;
      patterns[59085] = 29'b1_110011011001_101_0_111100110110;
      patterns[59086] = 29'b1_110011011001_110_1_110011011001;
      patterns[59087] = 29'b1_110011011001_111_1_110011011001;
      patterns[59088] = 29'b1_110011011010_000_1_110011011010;
      patterns[59089] = 29'b1_110011011010_001_1_011010110011;
      patterns[59090] = 29'b1_110011011010_010_1_100110110101;
      patterns[59091] = 29'b1_110011011010_011_1_001101101011;
      patterns[59092] = 29'b1_110011011010_100_0_111001101101;
      patterns[59093] = 29'b1_110011011010_101_1_011100110110;
      patterns[59094] = 29'b1_110011011010_110_1_110011011010;
      patterns[59095] = 29'b1_110011011010_111_1_110011011010;
      patterns[59096] = 29'b1_110011011011_000_1_110011011011;
      patterns[59097] = 29'b1_110011011011_001_1_011011110011;
      patterns[59098] = 29'b1_110011011011_010_1_100110110111;
      patterns[59099] = 29'b1_110011011011_011_1_001101101111;
      patterns[59100] = 29'b1_110011011011_100_1_111001101101;
      patterns[59101] = 29'b1_110011011011_101_1_111100110110;
      patterns[59102] = 29'b1_110011011011_110_1_110011011011;
      patterns[59103] = 29'b1_110011011011_111_1_110011011011;
      patterns[59104] = 29'b1_110011011100_000_1_110011011100;
      patterns[59105] = 29'b1_110011011100_001_1_011100110011;
      patterns[59106] = 29'b1_110011011100_010_1_100110111001;
      patterns[59107] = 29'b1_110011011100_011_1_001101110011;
      patterns[59108] = 29'b1_110011011100_100_0_111001101110;
      patterns[59109] = 29'b1_110011011100_101_0_011100110111;
      patterns[59110] = 29'b1_110011011100_110_1_110011011100;
      patterns[59111] = 29'b1_110011011100_111_1_110011011100;
      patterns[59112] = 29'b1_110011011101_000_1_110011011101;
      patterns[59113] = 29'b1_110011011101_001_1_011101110011;
      patterns[59114] = 29'b1_110011011101_010_1_100110111011;
      patterns[59115] = 29'b1_110011011101_011_1_001101110111;
      patterns[59116] = 29'b1_110011011101_100_1_111001101110;
      patterns[59117] = 29'b1_110011011101_101_0_111100110111;
      patterns[59118] = 29'b1_110011011101_110_1_110011011101;
      patterns[59119] = 29'b1_110011011101_111_1_110011011101;
      patterns[59120] = 29'b1_110011011110_000_1_110011011110;
      patterns[59121] = 29'b1_110011011110_001_1_011110110011;
      patterns[59122] = 29'b1_110011011110_010_1_100110111101;
      patterns[59123] = 29'b1_110011011110_011_1_001101111011;
      patterns[59124] = 29'b1_110011011110_100_0_111001101111;
      patterns[59125] = 29'b1_110011011110_101_1_011100110111;
      patterns[59126] = 29'b1_110011011110_110_1_110011011110;
      patterns[59127] = 29'b1_110011011110_111_1_110011011110;
      patterns[59128] = 29'b1_110011011111_000_1_110011011111;
      patterns[59129] = 29'b1_110011011111_001_1_011111110011;
      patterns[59130] = 29'b1_110011011111_010_1_100110111111;
      patterns[59131] = 29'b1_110011011111_011_1_001101111111;
      patterns[59132] = 29'b1_110011011111_100_1_111001101111;
      patterns[59133] = 29'b1_110011011111_101_1_111100110111;
      patterns[59134] = 29'b1_110011011111_110_1_110011011111;
      patterns[59135] = 29'b1_110011011111_111_1_110011011111;
      patterns[59136] = 29'b1_110011100000_000_1_110011100000;
      patterns[59137] = 29'b1_110011100000_001_1_100000110011;
      patterns[59138] = 29'b1_110011100000_010_1_100111000001;
      patterns[59139] = 29'b1_110011100000_011_1_001110000011;
      patterns[59140] = 29'b1_110011100000_100_0_111001110000;
      patterns[59141] = 29'b1_110011100000_101_0_011100111000;
      patterns[59142] = 29'b1_110011100000_110_1_110011100000;
      patterns[59143] = 29'b1_110011100000_111_1_110011100000;
      patterns[59144] = 29'b1_110011100001_000_1_110011100001;
      patterns[59145] = 29'b1_110011100001_001_1_100001110011;
      patterns[59146] = 29'b1_110011100001_010_1_100111000011;
      patterns[59147] = 29'b1_110011100001_011_1_001110000111;
      patterns[59148] = 29'b1_110011100001_100_1_111001110000;
      patterns[59149] = 29'b1_110011100001_101_0_111100111000;
      patterns[59150] = 29'b1_110011100001_110_1_110011100001;
      patterns[59151] = 29'b1_110011100001_111_1_110011100001;
      patterns[59152] = 29'b1_110011100010_000_1_110011100010;
      patterns[59153] = 29'b1_110011100010_001_1_100010110011;
      patterns[59154] = 29'b1_110011100010_010_1_100111000101;
      patterns[59155] = 29'b1_110011100010_011_1_001110001011;
      patterns[59156] = 29'b1_110011100010_100_0_111001110001;
      patterns[59157] = 29'b1_110011100010_101_1_011100111000;
      patterns[59158] = 29'b1_110011100010_110_1_110011100010;
      patterns[59159] = 29'b1_110011100010_111_1_110011100010;
      patterns[59160] = 29'b1_110011100011_000_1_110011100011;
      patterns[59161] = 29'b1_110011100011_001_1_100011110011;
      patterns[59162] = 29'b1_110011100011_010_1_100111000111;
      patterns[59163] = 29'b1_110011100011_011_1_001110001111;
      patterns[59164] = 29'b1_110011100011_100_1_111001110001;
      patterns[59165] = 29'b1_110011100011_101_1_111100111000;
      patterns[59166] = 29'b1_110011100011_110_1_110011100011;
      patterns[59167] = 29'b1_110011100011_111_1_110011100011;
      patterns[59168] = 29'b1_110011100100_000_1_110011100100;
      patterns[59169] = 29'b1_110011100100_001_1_100100110011;
      patterns[59170] = 29'b1_110011100100_010_1_100111001001;
      patterns[59171] = 29'b1_110011100100_011_1_001110010011;
      patterns[59172] = 29'b1_110011100100_100_0_111001110010;
      patterns[59173] = 29'b1_110011100100_101_0_011100111001;
      patterns[59174] = 29'b1_110011100100_110_1_110011100100;
      patterns[59175] = 29'b1_110011100100_111_1_110011100100;
      patterns[59176] = 29'b1_110011100101_000_1_110011100101;
      patterns[59177] = 29'b1_110011100101_001_1_100101110011;
      patterns[59178] = 29'b1_110011100101_010_1_100111001011;
      patterns[59179] = 29'b1_110011100101_011_1_001110010111;
      patterns[59180] = 29'b1_110011100101_100_1_111001110010;
      patterns[59181] = 29'b1_110011100101_101_0_111100111001;
      patterns[59182] = 29'b1_110011100101_110_1_110011100101;
      patterns[59183] = 29'b1_110011100101_111_1_110011100101;
      patterns[59184] = 29'b1_110011100110_000_1_110011100110;
      patterns[59185] = 29'b1_110011100110_001_1_100110110011;
      patterns[59186] = 29'b1_110011100110_010_1_100111001101;
      patterns[59187] = 29'b1_110011100110_011_1_001110011011;
      patterns[59188] = 29'b1_110011100110_100_0_111001110011;
      patterns[59189] = 29'b1_110011100110_101_1_011100111001;
      patterns[59190] = 29'b1_110011100110_110_1_110011100110;
      patterns[59191] = 29'b1_110011100110_111_1_110011100110;
      patterns[59192] = 29'b1_110011100111_000_1_110011100111;
      patterns[59193] = 29'b1_110011100111_001_1_100111110011;
      patterns[59194] = 29'b1_110011100111_010_1_100111001111;
      patterns[59195] = 29'b1_110011100111_011_1_001110011111;
      patterns[59196] = 29'b1_110011100111_100_1_111001110011;
      patterns[59197] = 29'b1_110011100111_101_1_111100111001;
      patterns[59198] = 29'b1_110011100111_110_1_110011100111;
      patterns[59199] = 29'b1_110011100111_111_1_110011100111;
      patterns[59200] = 29'b1_110011101000_000_1_110011101000;
      patterns[59201] = 29'b1_110011101000_001_1_101000110011;
      patterns[59202] = 29'b1_110011101000_010_1_100111010001;
      patterns[59203] = 29'b1_110011101000_011_1_001110100011;
      patterns[59204] = 29'b1_110011101000_100_0_111001110100;
      patterns[59205] = 29'b1_110011101000_101_0_011100111010;
      patterns[59206] = 29'b1_110011101000_110_1_110011101000;
      patterns[59207] = 29'b1_110011101000_111_1_110011101000;
      patterns[59208] = 29'b1_110011101001_000_1_110011101001;
      patterns[59209] = 29'b1_110011101001_001_1_101001110011;
      patterns[59210] = 29'b1_110011101001_010_1_100111010011;
      patterns[59211] = 29'b1_110011101001_011_1_001110100111;
      patterns[59212] = 29'b1_110011101001_100_1_111001110100;
      patterns[59213] = 29'b1_110011101001_101_0_111100111010;
      patterns[59214] = 29'b1_110011101001_110_1_110011101001;
      patterns[59215] = 29'b1_110011101001_111_1_110011101001;
      patterns[59216] = 29'b1_110011101010_000_1_110011101010;
      patterns[59217] = 29'b1_110011101010_001_1_101010110011;
      patterns[59218] = 29'b1_110011101010_010_1_100111010101;
      patterns[59219] = 29'b1_110011101010_011_1_001110101011;
      patterns[59220] = 29'b1_110011101010_100_0_111001110101;
      patterns[59221] = 29'b1_110011101010_101_1_011100111010;
      patterns[59222] = 29'b1_110011101010_110_1_110011101010;
      patterns[59223] = 29'b1_110011101010_111_1_110011101010;
      patterns[59224] = 29'b1_110011101011_000_1_110011101011;
      patterns[59225] = 29'b1_110011101011_001_1_101011110011;
      patterns[59226] = 29'b1_110011101011_010_1_100111010111;
      patterns[59227] = 29'b1_110011101011_011_1_001110101111;
      patterns[59228] = 29'b1_110011101011_100_1_111001110101;
      patterns[59229] = 29'b1_110011101011_101_1_111100111010;
      patterns[59230] = 29'b1_110011101011_110_1_110011101011;
      patterns[59231] = 29'b1_110011101011_111_1_110011101011;
      patterns[59232] = 29'b1_110011101100_000_1_110011101100;
      patterns[59233] = 29'b1_110011101100_001_1_101100110011;
      patterns[59234] = 29'b1_110011101100_010_1_100111011001;
      patterns[59235] = 29'b1_110011101100_011_1_001110110011;
      patterns[59236] = 29'b1_110011101100_100_0_111001110110;
      patterns[59237] = 29'b1_110011101100_101_0_011100111011;
      patterns[59238] = 29'b1_110011101100_110_1_110011101100;
      patterns[59239] = 29'b1_110011101100_111_1_110011101100;
      patterns[59240] = 29'b1_110011101101_000_1_110011101101;
      patterns[59241] = 29'b1_110011101101_001_1_101101110011;
      patterns[59242] = 29'b1_110011101101_010_1_100111011011;
      patterns[59243] = 29'b1_110011101101_011_1_001110110111;
      patterns[59244] = 29'b1_110011101101_100_1_111001110110;
      patterns[59245] = 29'b1_110011101101_101_0_111100111011;
      patterns[59246] = 29'b1_110011101101_110_1_110011101101;
      patterns[59247] = 29'b1_110011101101_111_1_110011101101;
      patterns[59248] = 29'b1_110011101110_000_1_110011101110;
      patterns[59249] = 29'b1_110011101110_001_1_101110110011;
      patterns[59250] = 29'b1_110011101110_010_1_100111011101;
      patterns[59251] = 29'b1_110011101110_011_1_001110111011;
      patterns[59252] = 29'b1_110011101110_100_0_111001110111;
      patterns[59253] = 29'b1_110011101110_101_1_011100111011;
      patterns[59254] = 29'b1_110011101110_110_1_110011101110;
      patterns[59255] = 29'b1_110011101110_111_1_110011101110;
      patterns[59256] = 29'b1_110011101111_000_1_110011101111;
      patterns[59257] = 29'b1_110011101111_001_1_101111110011;
      patterns[59258] = 29'b1_110011101111_010_1_100111011111;
      patterns[59259] = 29'b1_110011101111_011_1_001110111111;
      patterns[59260] = 29'b1_110011101111_100_1_111001110111;
      patterns[59261] = 29'b1_110011101111_101_1_111100111011;
      patterns[59262] = 29'b1_110011101111_110_1_110011101111;
      patterns[59263] = 29'b1_110011101111_111_1_110011101111;
      patterns[59264] = 29'b1_110011110000_000_1_110011110000;
      patterns[59265] = 29'b1_110011110000_001_1_110000110011;
      patterns[59266] = 29'b1_110011110000_010_1_100111100001;
      patterns[59267] = 29'b1_110011110000_011_1_001111000011;
      patterns[59268] = 29'b1_110011110000_100_0_111001111000;
      patterns[59269] = 29'b1_110011110000_101_0_011100111100;
      patterns[59270] = 29'b1_110011110000_110_1_110011110000;
      patterns[59271] = 29'b1_110011110000_111_1_110011110000;
      patterns[59272] = 29'b1_110011110001_000_1_110011110001;
      patterns[59273] = 29'b1_110011110001_001_1_110001110011;
      patterns[59274] = 29'b1_110011110001_010_1_100111100011;
      patterns[59275] = 29'b1_110011110001_011_1_001111000111;
      patterns[59276] = 29'b1_110011110001_100_1_111001111000;
      patterns[59277] = 29'b1_110011110001_101_0_111100111100;
      patterns[59278] = 29'b1_110011110001_110_1_110011110001;
      patterns[59279] = 29'b1_110011110001_111_1_110011110001;
      patterns[59280] = 29'b1_110011110010_000_1_110011110010;
      patterns[59281] = 29'b1_110011110010_001_1_110010110011;
      patterns[59282] = 29'b1_110011110010_010_1_100111100101;
      patterns[59283] = 29'b1_110011110010_011_1_001111001011;
      patterns[59284] = 29'b1_110011110010_100_0_111001111001;
      patterns[59285] = 29'b1_110011110010_101_1_011100111100;
      patterns[59286] = 29'b1_110011110010_110_1_110011110010;
      patterns[59287] = 29'b1_110011110010_111_1_110011110010;
      patterns[59288] = 29'b1_110011110011_000_1_110011110011;
      patterns[59289] = 29'b1_110011110011_001_1_110011110011;
      patterns[59290] = 29'b1_110011110011_010_1_100111100111;
      patterns[59291] = 29'b1_110011110011_011_1_001111001111;
      patterns[59292] = 29'b1_110011110011_100_1_111001111001;
      patterns[59293] = 29'b1_110011110011_101_1_111100111100;
      patterns[59294] = 29'b1_110011110011_110_1_110011110011;
      patterns[59295] = 29'b1_110011110011_111_1_110011110011;
      patterns[59296] = 29'b1_110011110100_000_1_110011110100;
      patterns[59297] = 29'b1_110011110100_001_1_110100110011;
      patterns[59298] = 29'b1_110011110100_010_1_100111101001;
      patterns[59299] = 29'b1_110011110100_011_1_001111010011;
      patterns[59300] = 29'b1_110011110100_100_0_111001111010;
      patterns[59301] = 29'b1_110011110100_101_0_011100111101;
      patterns[59302] = 29'b1_110011110100_110_1_110011110100;
      patterns[59303] = 29'b1_110011110100_111_1_110011110100;
      patterns[59304] = 29'b1_110011110101_000_1_110011110101;
      patterns[59305] = 29'b1_110011110101_001_1_110101110011;
      patterns[59306] = 29'b1_110011110101_010_1_100111101011;
      patterns[59307] = 29'b1_110011110101_011_1_001111010111;
      patterns[59308] = 29'b1_110011110101_100_1_111001111010;
      patterns[59309] = 29'b1_110011110101_101_0_111100111101;
      patterns[59310] = 29'b1_110011110101_110_1_110011110101;
      patterns[59311] = 29'b1_110011110101_111_1_110011110101;
      patterns[59312] = 29'b1_110011110110_000_1_110011110110;
      patterns[59313] = 29'b1_110011110110_001_1_110110110011;
      patterns[59314] = 29'b1_110011110110_010_1_100111101101;
      patterns[59315] = 29'b1_110011110110_011_1_001111011011;
      patterns[59316] = 29'b1_110011110110_100_0_111001111011;
      patterns[59317] = 29'b1_110011110110_101_1_011100111101;
      patterns[59318] = 29'b1_110011110110_110_1_110011110110;
      patterns[59319] = 29'b1_110011110110_111_1_110011110110;
      patterns[59320] = 29'b1_110011110111_000_1_110011110111;
      patterns[59321] = 29'b1_110011110111_001_1_110111110011;
      patterns[59322] = 29'b1_110011110111_010_1_100111101111;
      patterns[59323] = 29'b1_110011110111_011_1_001111011111;
      patterns[59324] = 29'b1_110011110111_100_1_111001111011;
      patterns[59325] = 29'b1_110011110111_101_1_111100111101;
      patterns[59326] = 29'b1_110011110111_110_1_110011110111;
      patterns[59327] = 29'b1_110011110111_111_1_110011110111;
      patterns[59328] = 29'b1_110011111000_000_1_110011111000;
      patterns[59329] = 29'b1_110011111000_001_1_111000110011;
      patterns[59330] = 29'b1_110011111000_010_1_100111110001;
      patterns[59331] = 29'b1_110011111000_011_1_001111100011;
      patterns[59332] = 29'b1_110011111000_100_0_111001111100;
      patterns[59333] = 29'b1_110011111000_101_0_011100111110;
      patterns[59334] = 29'b1_110011111000_110_1_110011111000;
      patterns[59335] = 29'b1_110011111000_111_1_110011111000;
      patterns[59336] = 29'b1_110011111001_000_1_110011111001;
      patterns[59337] = 29'b1_110011111001_001_1_111001110011;
      patterns[59338] = 29'b1_110011111001_010_1_100111110011;
      patterns[59339] = 29'b1_110011111001_011_1_001111100111;
      patterns[59340] = 29'b1_110011111001_100_1_111001111100;
      patterns[59341] = 29'b1_110011111001_101_0_111100111110;
      patterns[59342] = 29'b1_110011111001_110_1_110011111001;
      patterns[59343] = 29'b1_110011111001_111_1_110011111001;
      patterns[59344] = 29'b1_110011111010_000_1_110011111010;
      patterns[59345] = 29'b1_110011111010_001_1_111010110011;
      patterns[59346] = 29'b1_110011111010_010_1_100111110101;
      patterns[59347] = 29'b1_110011111010_011_1_001111101011;
      patterns[59348] = 29'b1_110011111010_100_0_111001111101;
      patterns[59349] = 29'b1_110011111010_101_1_011100111110;
      patterns[59350] = 29'b1_110011111010_110_1_110011111010;
      patterns[59351] = 29'b1_110011111010_111_1_110011111010;
      patterns[59352] = 29'b1_110011111011_000_1_110011111011;
      patterns[59353] = 29'b1_110011111011_001_1_111011110011;
      patterns[59354] = 29'b1_110011111011_010_1_100111110111;
      patterns[59355] = 29'b1_110011111011_011_1_001111101111;
      patterns[59356] = 29'b1_110011111011_100_1_111001111101;
      patterns[59357] = 29'b1_110011111011_101_1_111100111110;
      patterns[59358] = 29'b1_110011111011_110_1_110011111011;
      patterns[59359] = 29'b1_110011111011_111_1_110011111011;
      patterns[59360] = 29'b1_110011111100_000_1_110011111100;
      patterns[59361] = 29'b1_110011111100_001_1_111100110011;
      patterns[59362] = 29'b1_110011111100_010_1_100111111001;
      patterns[59363] = 29'b1_110011111100_011_1_001111110011;
      patterns[59364] = 29'b1_110011111100_100_0_111001111110;
      patterns[59365] = 29'b1_110011111100_101_0_011100111111;
      patterns[59366] = 29'b1_110011111100_110_1_110011111100;
      patterns[59367] = 29'b1_110011111100_111_1_110011111100;
      patterns[59368] = 29'b1_110011111101_000_1_110011111101;
      patterns[59369] = 29'b1_110011111101_001_1_111101110011;
      patterns[59370] = 29'b1_110011111101_010_1_100111111011;
      patterns[59371] = 29'b1_110011111101_011_1_001111110111;
      patterns[59372] = 29'b1_110011111101_100_1_111001111110;
      patterns[59373] = 29'b1_110011111101_101_0_111100111111;
      patterns[59374] = 29'b1_110011111101_110_1_110011111101;
      patterns[59375] = 29'b1_110011111101_111_1_110011111101;
      patterns[59376] = 29'b1_110011111110_000_1_110011111110;
      patterns[59377] = 29'b1_110011111110_001_1_111110110011;
      patterns[59378] = 29'b1_110011111110_010_1_100111111101;
      patterns[59379] = 29'b1_110011111110_011_1_001111111011;
      patterns[59380] = 29'b1_110011111110_100_0_111001111111;
      patterns[59381] = 29'b1_110011111110_101_1_011100111111;
      patterns[59382] = 29'b1_110011111110_110_1_110011111110;
      patterns[59383] = 29'b1_110011111110_111_1_110011111110;
      patterns[59384] = 29'b1_110011111111_000_1_110011111111;
      patterns[59385] = 29'b1_110011111111_001_1_111111110011;
      patterns[59386] = 29'b1_110011111111_010_1_100111111111;
      patterns[59387] = 29'b1_110011111111_011_1_001111111111;
      patterns[59388] = 29'b1_110011111111_100_1_111001111111;
      patterns[59389] = 29'b1_110011111111_101_1_111100111111;
      patterns[59390] = 29'b1_110011111111_110_1_110011111111;
      patterns[59391] = 29'b1_110011111111_111_1_110011111111;
      patterns[59392] = 29'b1_110100000000_000_1_110100000000;
      patterns[59393] = 29'b1_110100000000_001_1_000000110100;
      patterns[59394] = 29'b1_110100000000_010_1_101000000001;
      patterns[59395] = 29'b1_110100000000_011_1_010000000011;
      patterns[59396] = 29'b1_110100000000_100_0_111010000000;
      patterns[59397] = 29'b1_110100000000_101_0_011101000000;
      patterns[59398] = 29'b1_110100000000_110_1_110100000000;
      patterns[59399] = 29'b1_110100000000_111_1_110100000000;
      patterns[59400] = 29'b1_110100000001_000_1_110100000001;
      patterns[59401] = 29'b1_110100000001_001_1_000001110100;
      patterns[59402] = 29'b1_110100000001_010_1_101000000011;
      patterns[59403] = 29'b1_110100000001_011_1_010000000111;
      patterns[59404] = 29'b1_110100000001_100_1_111010000000;
      patterns[59405] = 29'b1_110100000001_101_0_111101000000;
      patterns[59406] = 29'b1_110100000001_110_1_110100000001;
      patterns[59407] = 29'b1_110100000001_111_1_110100000001;
      patterns[59408] = 29'b1_110100000010_000_1_110100000010;
      patterns[59409] = 29'b1_110100000010_001_1_000010110100;
      patterns[59410] = 29'b1_110100000010_010_1_101000000101;
      patterns[59411] = 29'b1_110100000010_011_1_010000001011;
      patterns[59412] = 29'b1_110100000010_100_0_111010000001;
      patterns[59413] = 29'b1_110100000010_101_1_011101000000;
      patterns[59414] = 29'b1_110100000010_110_1_110100000010;
      patterns[59415] = 29'b1_110100000010_111_1_110100000010;
      patterns[59416] = 29'b1_110100000011_000_1_110100000011;
      patterns[59417] = 29'b1_110100000011_001_1_000011110100;
      patterns[59418] = 29'b1_110100000011_010_1_101000000111;
      patterns[59419] = 29'b1_110100000011_011_1_010000001111;
      patterns[59420] = 29'b1_110100000011_100_1_111010000001;
      patterns[59421] = 29'b1_110100000011_101_1_111101000000;
      patterns[59422] = 29'b1_110100000011_110_1_110100000011;
      patterns[59423] = 29'b1_110100000011_111_1_110100000011;
      patterns[59424] = 29'b1_110100000100_000_1_110100000100;
      patterns[59425] = 29'b1_110100000100_001_1_000100110100;
      patterns[59426] = 29'b1_110100000100_010_1_101000001001;
      patterns[59427] = 29'b1_110100000100_011_1_010000010011;
      patterns[59428] = 29'b1_110100000100_100_0_111010000010;
      patterns[59429] = 29'b1_110100000100_101_0_011101000001;
      patterns[59430] = 29'b1_110100000100_110_1_110100000100;
      patterns[59431] = 29'b1_110100000100_111_1_110100000100;
      patterns[59432] = 29'b1_110100000101_000_1_110100000101;
      patterns[59433] = 29'b1_110100000101_001_1_000101110100;
      patterns[59434] = 29'b1_110100000101_010_1_101000001011;
      patterns[59435] = 29'b1_110100000101_011_1_010000010111;
      patterns[59436] = 29'b1_110100000101_100_1_111010000010;
      patterns[59437] = 29'b1_110100000101_101_0_111101000001;
      patterns[59438] = 29'b1_110100000101_110_1_110100000101;
      patterns[59439] = 29'b1_110100000101_111_1_110100000101;
      patterns[59440] = 29'b1_110100000110_000_1_110100000110;
      patterns[59441] = 29'b1_110100000110_001_1_000110110100;
      patterns[59442] = 29'b1_110100000110_010_1_101000001101;
      patterns[59443] = 29'b1_110100000110_011_1_010000011011;
      patterns[59444] = 29'b1_110100000110_100_0_111010000011;
      patterns[59445] = 29'b1_110100000110_101_1_011101000001;
      patterns[59446] = 29'b1_110100000110_110_1_110100000110;
      patterns[59447] = 29'b1_110100000110_111_1_110100000110;
      patterns[59448] = 29'b1_110100000111_000_1_110100000111;
      patterns[59449] = 29'b1_110100000111_001_1_000111110100;
      patterns[59450] = 29'b1_110100000111_010_1_101000001111;
      patterns[59451] = 29'b1_110100000111_011_1_010000011111;
      patterns[59452] = 29'b1_110100000111_100_1_111010000011;
      patterns[59453] = 29'b1_110100000111_101_1_111101000001;
      patterns[59454] = 29'b1_110100000111_110_1_110100000111;
      patterns[59455] = 29'b1_110100000111_111_1_110100000111;
      patterns[59456] = 29'b1_110100001000_000_1_110100001000;
      patterns[59457] = 29'b1_110100001000_001_1_001000110100;
      patterns[59458] = 29'b1_110100001000_010_1_101000010001;
      patterns[59459] = 29'b1_110100001000_011_1_010000100011;
      patterns[59460] = 29'b1_110100001000_100_0_111010000100;
      patterns[59461] = 29'b1_110100001000_101_0_011101000010;
      patterns[59462] = 29'b1_110100001000_110_1_110100001000;
      patterns[59463] = 29'b1_110100001000_111_1_110100001000;
      patterns[59464] = 29'b1_110100001001_000_1_110100001001;
      patterns[59465] = 29'b1_110100001001_001_1_001001110100;
      patterns[59466] = 29'b1_110100001001_010_1_101000010011;
      patterns[59467] = 29'b1_110100001001_011_1_010000100111;
      patterns[59468] = 29'b1_110100001001_100_1_111010000100;
      patterns[59469] = 29'b1_110100001001_101_0_111101000010;
      patterns[59470] = 29'b1_110100001001_110_1_110100001001;
      patterns[59471] = 29'b1_110100001001_111_1_110100001001;
      patterns[59472] = 29'b1_110100001010_000_1_110100001010;
      patterns[59473] = 29'b1_110100001010_001_1_001010110100;
      patterns[59474] = 29'b1_110100001010_010_1_101000010101;
      patterns[59475] = 29'b1_110100001010_011_1_010000101011;
      patterns[59476] = 29'b1_110100001010_100_0_111010000101;
      patterns[59477] = 29'b1_110100001010_101_1_011101000010;
      patterns[59478] = 29'b1_110100001010_110_1_110100001010;
      patterns[59479] = 29'b1_110100001010_111_1_110100001010;
      patterns[59480] = 29'b1_110100001011_000_1_110100001011;
      patterns[59481] = 29'b1_110100001011_001_1_001011110100;
      patterns[59482] = 29'b1_110100001011_010_1_101000010111;
      patterns[59483] = 29'b1_110100001011_011_1_010000101111;
      patterns[59484] = 29'b1_110100001011_100_1_111010000101;
      patterns[59485] = 29'b1_110100001011_101_1_111101000010;
      patterns[59486] = 29'b1_110100001011_110_1_110100001011;
      patterns[59487] = 29'b1_110100001011_111_1_110100001011;
      patterns[59488] = 29'b1_110100001100_000_1_110100001100;
      patterns[59489] = 29'b1_110100001100_001_1_001100110100;
      patterns[59490] = 29'b1_110100001100_010_1_101000011001;
      patterns[59491] = 29'b1_110100001100_011_1_010000110011;
      patterns[59492] = 29'b1_110100001100_100_0_111010000110;
      patterns[59493] = 29'b1_110100001100_101_0_011101000011;
      patterns[59494] = 29'b1_110100001100_110_1_110100001100;
      patterns[59495] = 29'b1_110100001100_111_1_110100001100;
      patterns[59496] = 29'b1_110100001101_000_1_110100001101;
      patterns[59497] = 29'b1_110100001101_001_1_001101110100;
      patterns[59498] = 29'b1_110100001101_010_1_101000011011;
      patterns[59499] = 29'b1_110100001101_011_1_010000110111;
      patterns[59500] = 29'b1_110100001101_100_1_111010000110;
      patterns[59501] = 29'b1_110100001101_101_0_111101000011;
      patterns[59502] = 29'b1_110100001101_110_1_110100001101;
      patterns[59503] = 29'b1_110100001101_111_1_110100001101;
      patterns[59504] = 29'b1_110100001110_000_1_110100001110;
      patterns[59505] = 29'b1_110100001110_001_1_001110110100;
      patterns[59506] = 29'b1_110100001110_010_1_101000011101;
      patterns[59507] = 29'b1_110100001110_011_1_010000111011;
      patterns[59508] = 29'b1_110100001110_100_0_111010000111;
      patterns[59509] = 29'b1_110100001110_101_1_011101000011;
      patterns[59510] = 29'b1_110100001110_110_1_110100001110;
      patterns[59511] = 29'b1_110100001110_111_1_110100001110;
      patterns[59512] = 29'b1_110100001111_000_1_110100001111;
      patterns[59513] = 29'b1_110100001111_001_1_001111110100;
      patterns[59514] = 29'b1_110100001111_010_1_101000011111;
      patterns[59515] = 29'b1_110100001111_011_1_010000111111;
      patterns[59516] = 29'b1_110100001111_100_1_111010000111;
      patterns[59517] = 29'b1_110100001111_101_1_111101000011;
      patterns[59518] = 29'b1_110100001111_110_1_110100001111;
      patterns[59519] = 29'b1_110100001111_111_1_110100001111;
      patterns[59520] = 29'b1_110100010000_000_1_110100010000;
      patterns[59521] = 29'b1_110100010000_001_1_010000110100;
      patterns[59522] = 29'b1_110100010000_010_1_101000100001;
      patterns[59523] = 29'b1_110100010000_011_1_010001000011;
      patterns[59524] = 29'b1_110100010000_100_0_111010001000;
      patterns[59525] = 29'b1_110100010000_101_0_011101000100;
      patterns[59526] = 29'b1_110100010000_110_1_110100010000;
      patterns[59527] = 29'b1_110100010000_111_1_110100010000;
      patterns[59528] = 29'b1_110100010001_000_1_110100010001;
      patterns[59529] = 29'b1_110100010001_001_1_010001110100;
      patterns[59530] = 29'b1_110100010001_010_1_101000100011;
      patterns[59531] = 29'b1_110100010001_011_1_010001000111;
      patterns[59532] = 29'b1_110100010001_100_1_111010001000;
      patterns[59533] = 29'b1_110100010001_101_0_111101000100;
      patterns[59534] = 29'b1_110100010001_110_1_110100010001;
      patterns[59535] = 29'b1_110100010001_111_1_110100010001;
      patterns[59536] = 29'b1_110100010010_000_1_110100010010;
      patterns[59537] = 29'b1_110100010010_001_1_010010110100;
      patterns[59538] = 29'b1_110100010010_010_1_101000100101;
      patterns[59539] = 29'b1_110100010010_011_1_010001001011;
      patterns[59540] = 29'b1_110100010010_100_0_111010001001;
      patterns[59541] = 29'b1_110100010010_101_1_011101000100;
      patterns[59542] = 29'b1_110100010010_110_1_110100010010;
      patterns[59543] = 29'b1_110100010010_111_1_110100010010;
      patterns[59544] = 29'b1_110100010011_000_1_110100010011;
      patterns[59545] = 29'b1_110100010011_001_1_010011110100;
      patterns[59546] = 29'b1_110100010011_010_1_101000100111;
      patterns[59547] = 29'b1_110100010011_011_1_010001001111;
      patterns[59548] = 29'b1_110100010011_100_1_111010001001;
      patterns[59549] = 29'b1_110100010011_101_1_111101000100;
      patterns[59550] = 29'b1_110100010011_110_1_110100010011;
      patterns[59551] = 29'b1_110100010011_111_1_110100010011;
      patterns[59552] = 29'b1_110100010100_000_1_110100010100;
      patterns[59553] = 29'b1_110100010100_001_1_010100110100;
      patterns[59554] = 29'b1_110100010100_010_1_101000101001;
      patterns[59555] = 29'b1_110100010100_011_1_010001010011;
      patterns[59556] = 29'b1_110100010100_100_0_111010001010;
      patterns[59557] = 29'b1_110100010100_101_0_011101000101;
      patterns[59558] = 29'b1_110100010100_110_1_110100010100;
      patterns[59559] = 29'b1_110100010100_111_1_110100010100;
      patterns[59560] = 29'b1_110100010101_000_1_110100010101;
      patterns[59561] = 29'b1_110100010101_001_1_010101110100;
      patterns[59562] = 29'b1_110100010101_010_1_101000101011;
      patterns[59563] = 29'b1_110100010101_011_1_010001010111;
      patterns[59564] = 29'b1_110100010101_100_1_111010001010;
      patterns[59565] = 29'b1_110100010101_101_0_111101000101;
      patterns[59566] = 29'b1_110100010101_110_1_110100010101;
      patterns[59567] = 29'b1_110100010101_111_1_110100010101;
      patterns[59568] = 29'b1_110100010110_000_1_110100010110;
      patterns[59569] = 29'b1_110100010110_001_1_010110110100;
      patterns[59570] = 29'b1_110100010110_010_1_101000101101;
      patterns[59571] = 29'b1_110100010110_011_1_010001011011;
      patterns[59572] = 29'b1_110100010110_100_0_111010001011;
      patterns[59573] = 29'b1_110100010110_101_1_011101000101;
      patterns[59574] = 29'b1_110100010110_110_1_110100010110;
      patterns[59575] = 29'b1_110100010110_111_1_110100010110;
      patterns[59576] = 29'b1_110100010111_000_1_110100010111;
      patterns[59577] = 29'b1_110100010111_001_1_010111110100;
      patterns[59578] = 29'b1_110100010111_010_1_101000101111;
      patterns[59579] = 29'b1_110100010111_011_1_010001011111;
      patterns[59580] = 29'b1_110100010111_100_1_111010001011;
      patterns[59581] = 29'b1_110100010111_101_1_111101000101;
      patterns[59582] = 29'b1_110100010111_110_1_110100010111;
      patterns[59583] = 29'b1_110100010111_111_1_110100010111;
      patterns[59584] = 29'b1_110100011000_000_1_110100011000;
      patterns[59585] = 29'b1_110100011000_001_1_011000110100;
      patterns[59586] = 29'b1_110100011000_010_1_101000110001;
      patterns[59587] = 29'b1_110100011000_011_1_010001100011;
      patterns[59588] = 29'b1_110100011000_100_0_111010001100;
      patterns[59589] = 29'b1_110100011000_101_0_011101000110;
      patterns[59590] = 29'b1_110100011000_110_1_110100011000;
      patterns[59591] = 29'b1_110100011000_111_1_110100011000;
      patterns[59592] = 29'b1_110100011001_000_1_110100011001;
      patterns[59593] = 29'b1_110100011001_001_1_011001110100;
      patterns[59594] = 29'b1_110100011001_010_1_101000110011;
      patterns[59595] = 29'b1_110100011001_011_1_010001100111;
      patterns[59596] = 29'b1_110100011001_100_1_111010001100;
      patterns[59597] = 29'b1_110100011001_101_0_111101000110;
      patterns[59598] = 29'b1_110100011001_110_1_110100011001;
      patterns[59599] = 29'b1_110100011001_111_1_110100011001;
      patterns[59600] = 29'b1_110100011010_000_1_110100011010;
      patterns[59601] = 29'b1_110100011010_001_1_011010110100;
      patterns[59602] = 29'b1_110100011010_010_1_101000110101;
      patterns[59603] = 29'b1_110100011010_011_1_010001101011;
      patterns[59604] = 29'b1_110100011010_100_0_111010001101;
      patterns[59605] = 29'b1_110100011010_101_1_011101000110;
      patterns[59606] = 29'b1_110100011010_110_1_110100011010;
      patterns[59607] = 29'b1_110100011010_111_1_110100011010;
      patterns[59608] = 29'b1_110100011011_000_1_110100011011;
      patterns[59609] = 29'b1_110100011011_001_1_011011110100;
      patterns[59610] = 29'b1_110100011011_010_1_101000110111;
      patterns[59611] = 29'b1_110100011011_011_1_010001101111;
      patterns[59612] = 29'b1_110100011011_100_1_111010001101;
      patterns[59613] = 29'b1_110100011011_101_1_111101000110;
      patterns[59614] = 29'b1_110100011011_110_1_110100011011;
      patterns[59615] = 29'b1_110100011011_111_1_110100011011;
      patterns[59616] = 29'b1_110100011100_000_1_110100011100;
      patterns[59617] = 29'b1_110100011100_001_1_011100110100;
      patterns[59618] = 29'b1_110100011100_010_1_101000111001;
      patterns[59619] = 29'b1_110100011100_011_1_010001110011;
      patterns[59620] = 29'b1_110100011100_100_0_111010001110;
      patterns[59621] = 29'b1_110100011100_101_0_011101000111;
      patterns[59622] = 29'b1_110100011100_110_1_110100011100;
      patterns[59623] = 29'b1_110100011100_111_1_110100011100;
      patterns[59624] = 29'b1_110100011101_000_1_110100011101;
      patterns[59625] = 29'b1_110100011101_001_1_011101110100;
      patterns[59626] = 29'b1_110100011101_010_1_101000111011;
      patterns[59627] = 29'b1_110100011101_011_1_010001110111;
      patterns[59628] = 29'b1_110100011101_100_1_111010001110;
      patterns[59629] = 29'b1_110100011101_101_0_111101000111;
      patterns[59630] = 29'b1_110100011101_110_1_110100011101;
      patterns[59631] = 29'b1_110100011101_111_1_110100011101;
      patterns[59632] = 29'b1_110100011110_000_1_110100011110;
      patterns[59633] = 29'b1_110100011110_001_1_011110110100;
      patterns[59634] = 29'b1_110100011110_010_1_101000111101;
      patterns[59635] = 29'b1_110100011110_011_1_010001111011;
      patterns[59636] = 29'b1_110100011110_100_0_111010001111;
      patterns[59637] = 29'b1_110100011110_101_1_011101000111;
      patterns[59638] = 29'b1_110100011110_110_1_110100011110;
      patterns[59639] = 29'b1_110100011110_111_1_110100011110;
      patterns[59640] = 29'b1_110100011111_000_1_110100011111;
      patterns[59641] = 29'b1_110100011111_001_1_011111110100;
      patterns[59642] = 29'b1_110100011111_010_1_101000111111;
      patterns[59643] = 29'b1_110100011111_011_1_010001111111;
      patterns[59644] = 29'b1_110100011111_100_1_111010001111;
      patterns[59645] = 29'b1_110100011111_101_1_111101000111;
      patterns[59646] = 29'b1_110100011111_110_1_110100011111;
      patterns[59647] = 29'b1_110100011111_111_1_110100011111;
      patterns[59648] = 29'b1_110100100000_000_1_110100100000;
      patterns[59649] = 29'b1_110100100000_001_1_100000110100;
      patterns[59650] = 29'b1_110100100000_010_1_101001000001;
      patterns[59651] = 29'b1_110100100000_011_1_010010000011;
      patterns[59652] = 29'b1_110100100000_100_0_111010010000;
      patterns[59653] = 29'b1_110100100000_101_0_011101001000;
      patterns[59654] = 29'b1_110100100000_110_1_110100100000;
      patterns[59655] = 29'b1_110100100000_111_1_110100100000;
      patterns[59656] = 29'b1_110100100001_000_1_110100100001;
      patterns[59657] = 29'b1_110100100001_001_1_100001110100;
      patterns[59658] = 29'b1_110100100001_010_1_101001000011;
      patterns[59659] = 29'b1_110100100001_011_1_010010000111;
      patterns[59660] = 29'b1_110100100001_100_1_111010010000;
      patterns[59661] = 29'b1_110100100001_101_0_111101001000;
      patterns[59662] = 29'b1_110100100001_110_1_110100100001;
      patterns[59663] = 29'b1_110100100001_111_1_110100100001;
      patterns[59664] = 29'b1_110100100010_000_1_110100100010;
      patterns[59665] = 29'b1_110100100010_001_1_100010110100;
      patterns[59666] = 29'b1_110100100010_010_1_101001000101;
      patterns[59667] = 29'b1_110100100010_011_1_010010001011;
      patterns[59668] = 29'b1_110100100010_100_0_111010010001;
      patterns[59669] = 29'b1_110100100010_101_1_011101001000;
      patterns[59670] = 29'b1_110100100010_110_1_110100100010;
      patterns[59671] = 29'b1_110100100010_111_1_110100100010;
      patterns[59672] = 29'b1_110100100011_000_1_110100100011;
      patterns[59673] = 29'b1_110100100011_001_1_100011110100;
      patterns[59674] = 29'b1_110100100011_010_1_101001000111;
      patterns[59675] = 29'b1_110100100011_011_1_010010001111;
      patterns[59676] = 29'b1_110100100011_100_1_111010010001;
      patterns[59677] = 29'b1_110100100011_101_1_111101001000;
      patterns[59678] = 29'b1_110100100011_110_1_110100100011;
      patterns[59679] = 29'b1_110100100011_111_1_110100100011;
      patterns[59680] = 29'b1_110100100100_000_1_110100100100;
      patterns[59681] = 29'b1_110100100100_001_1_100100110100;
      patterns[59682] = 29'b1_110100100100_010_1_101001001001;
      patterns[59683] = 29'b1_110100100100_011_1_010010010011;
      patterns[59684] = 29'b1_110100100100_100_0_111010010010;
      patterns[59685] = 29'b1_110100100100_101_0_011101001001;
      patterns[59686] = 29'b1_110100100100_110_1_110100100100;
      patterns[59687] = 29'b1_110100100100_111_1_110100100100;
      patterns[59688] = 29'b1_110100100101_000_1_110100100101;
      patterns[59689] = 29'b1_110100100101_001_1_100101110100;
      patterns[59690] = 29'b1_110100100101_010_1_101001001011;
      patterns[59691] = 29'b1_110100100101_011_1_010010010111;
      patterns[59692] = 29'b1_110100100101_100_1_111010010010;
      patterns[59693] = 29'b1_110100100101_101_0_111101001001;
      patterns[59694] = 29'b1_110100100101_110_1_110100100101;
      patterns[59695] = 29'b1_110100100101_111_1_110100100101;
      patterns[59696] = 29'b1_110100100110_000_1_110100100110;
      patterns[59697] = 29'b1_110100100110_001_1_100110110100;
      patterns[59698] = 29'b1_110100100110_010_1_101001001101;
      patterns[59699] = 29'b1_110100100110_011_1_010010011011;
      patterns[59700] = 29'b1_110100100110_100_0_111010010011;
      patterns[59701] = 29'b1_110100100110_101_1_011101001001;
      patterns[59702] = 29'b1_110100100110_110_1_110100100110;
      patterns[59703] = 29'b1_110100100110_111_1_110100100110;
      patterns[59704] = 29'b1_110100100111_000_1_110100100111;
      patterns[59705] = 29'b1_110100100111_001_1_100111110100;
      patterns[59706] = 29'b1_110100100111_010_1_101001001111;
      patterns[59707] = 29'b1_110100100111_011_1_010010011111;
      patterns[59708] = 29'b1_110100100111_100_1_111010010011;
      patterns[59709] = 29'b1_110100100111_101_1_111101001001;
      patterns[59710] = 29'b1_110100100111_110_1_110100100111;
      patterns[59711] = 29'b1_110100100111_111_1_110100100111;
      patterns[59712] = 29'b1_110100101000_000_1_110100101000;
      patterns[59713] = 29'b1_110100101000_001_1_101000110100;
      patterns[59714] = 29'b1_110100101000_010_1_101001010001;
      patterns[59715] = 29'b1_110100101000_011_1_010010100011;
      patterns[59716] = 29'b1_110100101000_100_0_111010010100;
      patterns[59717] = 29'b1_110100101000_101_0_011101001010;
      patterns[59718] = 29'b1_110100101000_110_1_110100101000;
      patterns[59719] = 29'b1_110100101000_111_1_110100101000;
      patterns[59720] = 29'b1_110100101001_000_1_110100101001;
      patterns[59721] = 29'b1_110100101001_001_1_101001110100;
      patterns[59722] = 29'b1_110100101001_010_1_101001010011;
      patterns[59723] = 29'b1_110100101001_011_1_010010100111;
      patterns[59724] = 29'b1_110100101001_100_1_111010010100;
      patterns[59725] = 29'b1_110100101001_101_0_111101001010;
      patterns[59726] = 29'b1_110100101001_110_1_110100101001;
      patterns[59727] = 29'b1_110100101001_111_1_110100101001;
      patterns[59728] = 29'b1_110100101010_000_1_110100101010;
      patterns[59729] = 29'b1_110100101010_001_1_101010110100;
      patterns[59730] = 29'b1_110100101010_010_1_101001010101;
      patterns[59731] = 29'b1_110100101010_011_1_010010101011;
      patterns[59732] = 29'b1_110100101010_100_0_111010010101;
      patterns[59733] = 29'b1_110100101010_101_1_011101001010;
      patterns[59734] = 29'b1_110100101010_110_1_110100101010;
      patterns[59735] = 29'b1_110100101010_111_1_110100101010;
      patterns[59736] = 29'b1_110100101011_000_1_110100101011;
      patterns[59737] = 29'b1_110100101011_001_1_101011110100;
      patterns[59738] = 29'b1_110100101011_010_1_101001010111;
      patterns[59739] = 29'b1_110100101011_011_1_010010101111;
      patterns[59740] = 29'b1_110100101011_100_1_111010010101;
      patterns[59741] = 29'b1_110100101011_101_1_111101001010;
      patterns[59742] = 29'b1_110100101011_110_1_110100101011;
      patterns[59743] = 29'b1_110100101011_111_1_110100101011;
      patterns[59744] = 29'b1_110100101100_000_1_110100101100;
      patterns[59745] = 29'b1_110100101100_001_1_101100110100;
      patterns[59746] = 29'b1_110100101100_010_1_101001011001;
      patterns[59747] = 29'b1_110100101100_011_1_010010110011;
      patterns[59748] = 29'b1_110100101100_100_0_111010010110;
      patterns[59749] = 29'b1_110100101100_101_0_011101001011;
      patterns[59750] = 29'b1_110100101100_110_1_110100101100;
      patterns[59751] = 29'b1_110100101100_111_1_110100101100;
      patterns[59752] = 29'b1_110100101101_000_1_110100101101;
      patterns[59753] = 29'b1_110100101101_001_1_101101110100;
      patterns[59754] = 29'b1_110100101101_010_1_101001011011;
      patterns[59755] = 29'b1_110100101101_011_1_010010110111;
      patterns[59756] = 29'b1_110100101101_100_1_111010010110;
      patterns[59757] = 29'b1_110100101101_101_0_111101001011;
      patterns[59758] = 29'b1_110100101101_110_1_110100101101;
      patterns[59759] = 29'b1_110100101101_111_1_110100101101;
      patterns[59760] = 29'b1_110100101110_000_1_110100101110;
      patterns[59761] = 29'b1_110100101110_001_1_101110110100;
      patterns[59762] = 29'b1_110100101110_010_1_101001011101;
      patterns[59763] = 29'b1_110100101110_011_1_010010111011;
      patterns[59764] = 29'b1_110100101110_100_0_111010010111;
      patterns[59765] = 29'b1_110100101110_101_1_011101001011;
      patterns[59766] = 29'b1_110100101110_110_1_110100101110;
      patterns[59767] = 29'b1_110100101110_111_1_110100101110;
      patterns[59768] = 29'b1_110100101111_000_1_110100101111;
      patterns[59769] = 29'b1_110100101111_001_1_101111110100;
      patterns[59770] = 29'b1_110100101111_010_1_101001011111;
      patterns[59771] = 29'b1_110100101111_011_1_010010111111;
      patterns[59772] = 29'b1_110100101111_100_1_111010010111;
      patterns[59773] = 29'b1_110100101111_101_1_111101001011;
      patterns[59774] = 29'b1_110100101111_110_1_110100101111;
      patterns[59775] = 29'b1_110100101111_111_1_110100101111;
      patterns[59776] = 29'b1_110100110000_000_1_110100110000;
      patterns[59777] = 29'b1_110100110000_001_1_110000110100;
      patterns[59778] = 29'b1_110100110000_010_1_101001100001;
      patterns[59779] = 29'b1_110100110000_011_1_010011000011;
      patterns[59780] = 29'b1_110100110000_100_0_111010011000;
      patterns[59781] = 29'b1_110100110000_101_0_011101001100;
      patterns[59782] = 29'b1_110100110000_110_1_110100110000;
      patterns[59783] = 29'b1_110100110000_111_1_110100110000;
      patterns[59784] = 29'b1_110100110001_000_1_110100110001;
      patterns[59785] = 29'b1_110100110001_001_1_110001110100;
      patterns[59786] = 29'b1_110100110001_010_1_101001100011;
      patterns[59787] = 29'b1_110100110001_011_1_010011000111;
      patterns[59788] = 29'b1_110100110001_100_1_111010011000;
      patterns[59789] = 29'b1_110100110001_101_0_111101001100;
      patterns[59790] = 29'b1_110100110001_110_1_110100110001;
      patterns[59791] = 29'b1_110100110001_111_1_110100110001;
      patterns[59792] = 29'b1_110100110010_000_1_110100110010;
      patterns[59793] = 29'b1_110100110010_001_1_110010110100;
      patterns[59794] = 29'b1_110100110010_010_1_101001100101;
      patterns[59795] = 29'b1_110100110010_011_1_010011001011;
      patterns[59796] = 29'b1_110100110010_100_0_111010011001;
      patterns[59797] = 29'b1_110100110010_101_1_011101001100;
      patterns[59798] = 29'b1_110100110010_110_1_110100110010;
      patterns[59799] = 29'b1_110100110010_111_1_110100110010;
      patterns[59800] = 29'b1_110100110011_000_1_110100110011;
      patterns[59801] = 29'b1_110100110011_001_1_110011110100;
      patterns[59802] = 29'b1_110100110011_010_1_101001100111;
      patterns[59803] = 29'b1_110100110011_011_1_010011001111;
      patterns[59804] = 29'b1_110100110011_100_1_111010011001;
      patterns[59805] = 29'b1_110100110011_101_1_111101001100;
      patterns[59806] = 29'b1_110100110011_110_1_110100110011;
      patterns[59807] = 29'b1_110100110011_111_1_110100110011;
      patterns[59808] = 29'b1_110100110100_000_1_110100110100;
      patterns[59809] = 29'b1_110100110100_001_1_110100110100;
      patterns[59810] = 29'b1_110100110100_010_1_101001101001;
      patterns[59811] = 29'b1_110100110100_011_1_010011010011;
      patterns[59812] = 29'b1_110100110100_100_0_111010011010;
      patterns[59813] = 29'b1_110100110100_101_0_011101001101;
      patterns[59814] = 29'b1_110100110100_110_1_110100110100;
      patterns[59815] = 29'b1_110100110100_111_1_110100110100;
      patterns[59816] = 29'b1_110100110101_000_1_110100110101;
      patterns[59817] = 29'b1_110100110101_001_1_110101110100;
      patterns[59818] = 29'b1_110100110101_010_1_101001101011;
      patterns[59819] = 29'b1_110100110101_011_1_010011010111;
      patterns[59820] = 29'b1_110100110101_100_1_111010011010;
      patterns[59821] = 29'b1_110100110101_101_0_111101001101;
      patterns[59822] = 29'b1_110100110101_110_1_110100110101;
      patterns[59823] = 29'b1_110100110101_111_1_110100110101;
      patterns[59824] = 29'b1_110100110110_000_1_110100110110;
      patterns[59825] = 29'b1_110100110110_001_1_110110110100;
      patterns[59826] = 29'b1_110100110110_010_1_101001101101;
      patterns[59827] = 29'b1_110100110110_011_1_010011011011;
      patterns[59828] = 29'b1_110100110110_100_0_111010011011;
      patterns[59829] = 29'b1_110100110110_101_1_011101001101;
      patterns[59830] = 29'b1_110100110110_110_1_110100110110;
      patterns[59831] = 29'b1_110100110110_111_1_110100110110;
      patterns[59832] = 29'b1_110100110111_000_1_110100110111;
      patterns[59833] = 29'b1_110100110111_001_1_110111110100;
      patterns[59834] = 29'b1_110100110111_010_1_101001101111;
      patterns[59835] = 29'b1_110100110111_011_1_010011011111;
      patterns[59836] = 29'b1_110100110111_100_1_111010011011;
      patterns[59837] = 29'b1_110100110111_101_1_111101001101;
      patterns[59838] = 29'b1_110100110111_110_1_110100110111;
      patterns[59839] = 29'b1_110100110111_111_1_110100110111;
      patterns[59840] = 29'b1_110100111000_000_1_110100111000;
      patterns[59841] = 29'b1_110100111000_001_1_111000110100;
      patterns[59842] = 29'b1_110100111000_010_1_101001110001;
      patterns[59843] = 29'b1_110100111000_011_1_010011100011;
      patterns[59844] = 29'b1_110100111000_100_0_111010011100;
      patterns[59845] = 29'b1_110100111000_101_0_011101001110;
      patterns[59846] = 29'b1_110100111000_110_1_110100111000;
      patterns[59847] = 29'b1_110100111000_111_1_110100111000;
      patterns[59848] = 29'b1_110100111001_000_1_110100111001;
      patterns[59849] = 29'b1_110100111001_001_1_111001110100;
      patterns[59850] = 29'b1_110100111001_010_1_101001110011;
      patterns[59851] = 29'b1_110100111001_011_1_010011100111;
      patterns[59852] = 29'b1_110100111001_100_1_111010011100;
      patterns[59853] = 29'b1_110100111001_101_0_111101001110;
      patterns[59854] = 29'b1_110100111001_110_1_110100111001;
      patterns[59855] = 29'b1_110100111001_111_1_110100111001;
      patterns[59856] = 29'b1_110100111010_000_1_110100111010;
      patterns[59857] = 29'b1_110100111010_001_1_111010110100;
      patterns[59858] = 29'b1_110100111010_010_1_101001110101;
      patterns[59859] = 29'b1_110100111010_011_1_010011101011;
      patterns[59860] = 29'b1_110100111010_100_0_111010011101;
      patterns[59861] = 29'b1_110100111010_101_1_011101001110;
      patterns[59862] = 29'b1_110100111010_110_1_110100111010;
      patterns[59863] = 29'b1_110100111010_111_1_110100111010;
      patterns[59864] = 29'b1_110100111011_000_1_110100111011;
      patterns[59865] = 29'b1_110100111011_001_1_111011110100;
      patterns[59866] = 29'b1_110100111011_010_1_101001110111;
      patterns[59867] = 29'b1_110100111011_011_1_010011101111;
      patterns[59868] = 29'b1_110100111011_100_1_111010011101;
      patterns[59869] = 29'b1_110100111011_101_1_111101001110;
      patterns[59870] = 29'b1_110100111011_110_1_110100111011;
      patterns[59871] = 29'b1_110100111011_111_1_110100111011;
      patterns[59872] = 29'b1_110100111100_000_1_110100111100;
      patterns[59873] = 29'b1_110100111100_001_1_111100110100;
      patterns[59874] = 29'b1_110100111100_010_1_101001111001;
      patterns[59875] = 29'b1_110100111100_011_1_010011110011;
      patterns[59876] = 29'b1_110100111100_100_0_111010011110;
      patterns[59877] = 29'b1_110100111100_101_0_011101001111;
      patterns[59878] = 29'b1_110100111100_110_1_110100111100;
      patterns[59879] = 29'b1_110100111100_111_1_110100111100;
      patterns[59880] = 29'b1_110100111101_000_1_110100111101;
      patterns[59881] = 29'b1_110100111101_001_1_111101110100;
      patterns[59882] = 29'b1_110100111101_010_1_101001111011;
      patterns[59883] = 29'b1_110100111101_011_1_010011110111;
      patterns[59884] = 29'b1_110100111101_100_1_111010011110;
      patterns[59885] = 29'b1_110100111101_101_0_111101001111;
      patterns[59886] = 29'b1_110100111101_110_1_110100111101;
      patterns[59887] = 29'b1_110100111101_111_1_110100111101;
      patterns[59888] = 29'b1_110100111110_000_1_110100111110;
      patterns[59889] = 29'b1_110100111110_001_1_111110110100;
      patterns[59890] = 29'b1_110100111110_010_1_101001111101;
      patterns[59891] = 29'b1_110100111110_011_1_010011111011;
      patterns[59892] = 29'b1_110100111110_100_0_111010011111;
      patterns[59893] = 29'b1_110100111110_101_1_011101001111;
      patterns[59894] = 29'b1_110100111110_110_1_110100111110;
      patterns[59895] = 29'b1_110100111110_111_1_110100111110;
      patterns[59896] = 29'b1_110100111111_000_1_110100111111;
      patterns[59897] = 29'b1_110100111111_001_1_111111110100;
      patterns[59898] = 29'b1_110100111111_010_1_101001111111;
      patterns[59899] = 29'b1_110100111111_011_1_010011111111;
      patterns[59900] = 29'b1_110100111111_100_1_111010011111;
      patterns[59901] = 29'b1_110100111111_101_1_111101001111;
      patterns[59902] = 29'b1_110100111111_110_1_110100111111;
      patterns[59903] = 29'b1_110100111111_111_1_110100111111;
      patterns[59904] = 29'b1_110101000000_000_1_110101000000;
      patterns[59905] = 29'b1_110101000000_001_1_000000110101;
      patterns[59906] = 29'b1_110101000000_010_1_101010000001;
      patterns[59907] = 29'b1_110101000000_011_1_010100000011;
      patterns[59908] = 29'b1_110101000000_100_0_111010100000;
      patterns[59909] = 29'b1_110101000000_101_0_011101010000;
      patterns[59910] = 29'b1_110101000000_110_1_110101000000;
      patterns[59911] = 29'b1_110101000000_111_1_110101000000;
      patterns[59912] = 29'b1_110101000001_000_1_110101000001;
      patterns[59913] = 29'b1_110101000001_001_1_000001110101;
      patterns[59914] = 29'b1_110101000001_010_1_101010000011;
      patterns[59915] = 29'b1_110101000001_011_1_010100000111;
      patterns[59916] = 29'b1_110101000001_100_1_111010100000;
      patterns[59917] = 29'b1_110101000001_101_0_111101010000;
      patterns[59918] = 29'b1_110101000001_110_1_110101000001;
      patterns[59919] = 29'b1_110101000001_111_1_110101000001;
      patterns[59920] = 29'b1_110101000010_000_1_110101000010;
      patterns[59921] = 29'b1_110101000010_001_1_000010110101;
      patterns[59922] = 29'b1_110101000010_010_1_101010000101;
      patterns[59923] = 29'b1_110101000010_011_1_010100001011;
      patterns[59924] = 29'b1_110101000010_100_0_111010100001;
      patterns[59925] = 29'b1_110101000010_101_1_011101010000;
      patterns[59926] = 29'b1_110101000010_110_1_110101000010;
      patterns[59927] = 29'b1_110101000010_111_1_110101000010;
      patterns[59928] = 29'b1_110101000011_000_1_110101000011;
      patterns[59929] = 29'b1_110101000011_001_1_000011110101;
      patterns[59930] = 29'b1_110101000011_010_1_101010000111;
      patterns[59931] = 29'b1_110101000011_011_1_010100001111;
      patterns[59932] = 29'b1_110101000011_100_1_111010100001;
      patterns[59933] = 29'b1_110101000011_101_1_111101010000;
      patterns[59934] = 29'b1_110101000011_110_1_110101000011;
      patterns[59935] = 29'b1_110101000011_111_1_110101000011;
      patterns[59936] = 29'b1_110101000100_000_1_110101000100;
      patterns[59937] = 29'b1_110101000100_001_1_000100110101;
      patterns[59938] = 29'b1_110101000100_010_1_101010001001;
      patterns[59939] = 29'b1_110101000100_011_1_010100010011;
      patterns[59940] = 29'b1_110101000100_100_0_111010100010;
      patterns[59941] = 29'b1_110101000100_101_0_011101010001;
      patterns[59942] = 29'b1_110101000100_110_1_110101000100;
      patterns[59943] = 29'b1_110101000100_111_1_110101000100;
      patterns[59944] = 29'b1_110101000101_000_1_110101000101;
      patterns[59945] = 29'b1_110101000101_001_1_000101110101;
      patterns[59946] = 29'b1_110101000101_010_1_101010001011;
      patterns[59947] = 29'b1_110101000101_011_1_010100010111;
      patterns[59948] = 29'b1_110101000101_100_1_111010100010;
      patterns[59949] = 29'b1_110101000101_101_0_111101010001;
      patterns[59950] = 29'b1_110101000101_110_1_110101000101;
      patterns[59951] = 29'b1_110101000101_111_1_110101000101;
      patterns[59952] = 29'b1_110101000110_000_1_110101000110;
      patterns[59953] = 29'b1_110101000110_001_1_000110110101;
      patterns[59954] = 29'b1_110101000110_010_1_101010001101;
      patterns[59955] = 29'b1_110101000110_011_1_010100011011;
      patterns[59956] = 29'b1_110101000110_100_0_111010100011;
      patterns[59957] = 29'b1_110101000110_101_1_011101010001;
      patterns[59958] = 29'b1_110101000110_110_1_110101000110;
      patterns[59959] = 29'b1_110101000110_111_1_110101000110;
      patterns[59960] = 29'b1_110101000111_000_1_110101000111;
      patterns[59961] = 29'b1_110101000111_001_1_000111110101;
      patterns[59962] = 29'b1_110101000111_010_1_101010001111;
      patterns[59963] = 29'b1_110101000111_011_1_010100011111;
      patterns[59964] = 29'b1_110101000111_100_1_111010100011;
      patterns[59965] = 29'b1_110101000111_101_1_111101010001;
      patterns[59966] = 29'b1_110101000111_110_1_110101000111;
      patterns[59967] = 29'b1_110101000111_111_1_110101000111;
      patterns[59968] = 29'b1_110101001000_000_1_110101001000;
      patterns[59969] = 29'b1_110101001000_001_1_001000110101;
      patterns[59970] = 29'b1_110101001000_010_1_101010010001;
      patterns[59971] = 29'b1_110101001000_011_1_010100100011;
      patterns[59972] = 29'b1_110101001000_100_0_111010100100;
      patterns[59973] = 29'b1_110101001000_101_0_011101010010;
      patterns[59974] = 29'b1_110101001000_110_1_110101001000;
      patterns[59975] = 29'b1_110101001000_111_1_110101001000;
      patterns[59976] = 29'b1_110101001001_000_1_110101001001;
      patterns[59977] = 29'b1_110101001001_001_1_001001110101;
      patterns[59978] = 29'b1_110101001001_010_1_101010010011;
      patterns[59979] = 29'b1_110101001001_011_1_010100100111;
      patterns[59980] = 29'b1_110101001001_100_1_111010100100;
      patterns[59981] = 29'b1_110101001001_101_0_111101010010;
      patterns[59982] = 29'b1_110101001001_110_1_110101001001;
      patterns[59983] = 29'b1_110101001001_111_1_110101001001;
      patterns[59984] = 29'b1_110101001010_000_1_110101001010;
      patterns[59985] = 29'b1_110101001010_001_1_001010110101;
      patterns[59986] = 29'b1_110101001010_010_1_101010010101;
      patterns[59987] = 29'b1_110101001010_011_1_010100101011;
      patterns[59988] = 29'b1_110101001010_100_0_111010100101;
      patterns[59989] = 29'b1_110101001010_101_1_011101010010;
      patterns[59990] = 29'b1_110101001010_110_1_110101001010;
      patterns[59991] = 29'b1_110101001010_111_1_110101001010;
      patterns[59992] = 29'b1_110101001011_000_1_110101001011;
      patterns[59993] = 29'b1_110101001011_001_1_001011110101;
      patterns[59994] = 29'b1_110101001011_010_1_101010010111;
      patterns[59995] = 29'b1_110101001011_011_1_010100101111;
      patterns[59996] = 29'b1_110101001011_100_1_111010100101;
      patterns[59997] = 29'b1_110101001011_101_1_111101010010;
      patterns[59998] = 29'b1_110101001011_110_1_110101001011;
      patterns[59999] = 29'b1_110101001011_111_1_110101001011;
      patterns[60000] = 29'b1_110101001100_000_1_110101001100;
      patterns[60001] = 29'b1_110101001100_001_1_001100110101;
      patterns[60002] = 29'b1_110101001100_010_1_101010011001;
      patterns[60003] = 29'b1_110101001100_011_1_010100110011;
      patterns[60004] = 29'b1_110101001100_100_0_111010100110;
      patterns[60005] = 29'b1_110101001100_101_0_011101010011;
      patterns[60006] = 29'b1_110101001100_110_1_110101001100;
      patterns[60007] = 29'b1_110101001100_111_1_110101001100;
      patterns[60008] = 29'b1_110101001101_000_1_110101001101;
      patterns[60009] = 29'b1_110101001101_001_1_001101110101;
      patterns[60010] = 29'b1_110101001101_010_1_101010011011;
      patterns[60011] = 29'b1_110101001101_011_1_010100110111;
      patterns[60012] = 29'b1_110101001101_100_1_111010100110;
      patterns[60013] = 29'b1_110101001101_101_0_111101010011;
      patterns[60014] = 29'b1_110101001101_110_1_110101001101;
      patterns[60015] = 29'b1_110101001101_111_1_110101001101;
      patterns[60016] = 29'b1_110101001110_000_1_110101001110;
      patterns[60017] = 29'b1_110101001110_001_1_001110110101;
      patterns[60018] = 29'b1_110101001110_010_1_101010011101;
      patterns[60019] = 29'b1_110101001110_011_1_010100111011;
      patterns[60020] = 29'b1_110101001110_100_0_111010100111;
      patterns[60021] = 29'b1_110101001110_101_1_011101010011;
      patterns[60022] = 29'b1_110101001110_110_1_110101001110;
      patterns[60023] = 29'b1_110101001110_111_1_110101001110;
      patterns[60024] = 29'b1_110101001111_000_1_110101001111;
      patterns[60025] = 29'b1_110101001111_001_1_001111110101;
      patterns[60026] = 29'b1_110101001111_010_1_101010011111;
      patterns[60027] = 29'b1_110101001111_011_1_010100111111;
      patterns[60028] = 29'b1_110101001111_100_1_111010100111;
      patterns[60029] = 29'b1_110101001111_101_1_111101010011;
      patterns[60030] = 29'b1_110101001111_110_1_110101001111;
      patterns[60031] = 29'b1_110101001111_111_1_110101001111;
      patterns[60032] = 29'b1_110101010000_000_1_110101010000;
      patterns[60033] = 29'b1_110101010000_001_1_010000110101;
      patterns[60034] = 29'b1_110101010000_010_1_101010100001;
      patterns[60035] = 29'b1_110101010000_011_1_010101000011;
      patterns[60036] = 29'b1_110101010000_100_0_111010101000;
      patterns[60037] = 29'b1_110101010000_101_0_011101010100;
      patterns[60038] = 29'b1_110101010000_110_1_110101010000;
      patterns[60039] = 29'b1_110101010000_111_1_110101010000;
      patterns[60040] = 29'b1_110101010001_000_1_110101010001;
      patterns[60041] = 29'b1_110101010001_001_1_010001110101;
      patterns[60042] = 29'b1_110101010001_010_1_101010100011;
      patterns[60043] = 29'b1_110101010001_011_1_010101000111;
      patterns[60044] = 29'b1_110101010001_100_1_111010101000;
      patterns[60045] = 29'b1_110101010001_101_0_111101010100;
      patterns[60046] = 29'b1_110101010001_110_1_110101010001;
      patterns[60047] = 29'b1_110101010001_111_1_110101010001;
      patterns[60048] = 29'b1_110101010010_000_1_110101010010;
      patterns[60049] = 29'b1_110101010010_001_1_010010110101;
      patterns[60050] = 29'b1_110101010010_010_1_101010100101;
      patterns[60051] = 29'b1_110101010010_011_1_010101001011;
      patterns[60052] = 29'b1_110101010010_100_0_111010101001;
      patterns[60053] = 29'b1_110101010010_101_1_011101010100;
      patterns[60054] = 29'b1_110101010010_110_1_110101010010;
      patterns[60055] = 29'b1_110101010010_111_1_110101010010;
      patterns[60056] = 29'b1_110101010011_000_1_110101010011;
      patterns[60057] = 29'b1_110101010011_001_1_010011110101;
      patterns[60058] = 29'b1_110101010011_010_1_101010100111;
      patterns[60059] = 29'b1_110101010011_011_1_010101001111;
      patterns[60060] = 29'b1_110101010011_100_1_111010101001;
      patterns[60061] = 29'b1_110101010011_101_1_111101010100;
      patterns[60062] = 29'b1_110101010011_110_1_110101010011;
      patterns[60063] = 29'b1_110101010011_111_1_110101010011;
      patterns[60064] = 29'b1_110101010100_000_1_110101010100;
      patterns[60065] = 29'b1_110101010100_001_1_010100110101;
      patterns[60066] = 29'b1_110101010100_010_1_101010101001;
      patterns[60067] = 29'b1_110101010100_011_1_010101010011;
      patterns[60068] = 29'b1_110101010100_100_0_111010101010;
      patterns[60069] = 29'b1_110101010100_101_0_011101010101;
      patterns[60070] = 29'b1_110101010100_110_1_110101010100;
      patterns[60071] = 29'b1_110101010100_111_1_110101010100;
      patterns[60072] = 29'b1_110101010101_000_1_110101010101;
      patterns[60073] = 29'b1_110101010101_001_1_010101110101;
      patterns[60074] = 29'b1_110101010101_010_1_101010101011;
      patterns[60075] = 29'b1_110101010101_011_1_010101010111;
      patterns[60076] = 29'b1_110101010101_100_1_111010101010;
      patterns[60077] = 29'b1_110101010101_101_0_111101010101;
      patterns[60078] = 29'b1_110101010101_110_1_110101010101;
      patterns[60079] = 29'b1_110101010101_111_1_110101010101;
      patterns[60080] = 29'b1_110101010110_000_1_110101010110;
      patterns[60081] = 29'b1_110101010110_001_1_010110110101;
      patterns[60082] = 29'b1_110101010110_010_1_101010101101;
      patterns[60083] = 29'b1_110101010110_011_1_010101011011;
      patterns[60084] = 29'b1_110101010110_100_0_111010101011;
      patterns[60085] = 29'b1_110101010110_101_1_011101010101;
      patterns[60086] = 29'b1_110101010110_110_1_110101010110;
      patterns[60087] = 29'b1_110101010110_111_1_110101010110;
      patterns[60088] = 29'b1_110101010111_000_1_110101010111;
      patterns[60089] = 29'b1_110101010111_001_1_010111110101;
      patterns[60090] = 29'b1_110101010111_010_1_101010101111;
      patterns[60091] = 29'b1_110101010111_011_1_010101011111;
      patterns[60092] = 29'b1_110101010111_100_1_111010101011;
      patterns[60093] = 29'b1_110101010111_101_1_111101010101;
      patterns[60094] = 29'b1_110101010111_110_1_110101010111;
      patterns[60095] = 29'b1_110101010111_111_1_110101010111;
      patterns[60096] = 29'b1_110101011000_000_1_110101011000;
      patterns[60097] = 29'b1_110101011000_001_1_011000110101;
      patterns[60098] = 29'b1_110101011000_010_1_101010110001;
      patterns[60099] = 29'b1_110101011000_011_1_010101100011;
      patterns[60100] = 29'b1_110101011000_100_0_111010101100;
      patterns[60101] = 29'b1_110101011000_101_0_011101010110;
      patterns[60102] = 29'b1_110101011000_110_1_110101011000;
      patterns[60103] = 29'b1_110101011000_111_1_110101011000;
      patterns[60104] = 29'b1_110101011001_000_1_110101011001;
      patterns[60105] = 29'b1_110101011001_001_1_011001110101;
      patterns[60106] = 29'b1_110101011001_010_1_101010110011;
      patterns[60107] = 29'b1_110101011001_011_1_010101100111;
      patterns[60108] = 29'b1_110101011001_100_1_111010101100;
      patterns[60109] = 29'b1_110101011001_101_0_111101010110;
      patterns[60110] = 29'b1_110101011001_110_1_110101011001;
      patterns[60111] = 29'b1_110101011001_111_1_110101011001;
      patterns[60112] = 29'b1_110101011010_000_1_110101011010;
      patterns[60113] = 29'b1_110101011010_001_1_011010110101;
      patterns[60114] = 29'b1_110101011010_010_1_101010110101;
      patterns[60115] = 29'b1_110101011010_011_1_010101101011;
      patterns[60116] = 29'b1_110101011010_100_0_111010101101;
      patterns[60117] = 29'b1_110101011010_101_1_011101010110;
      patterns[60118] = 29'b1_110101011010_110_1_110101011010;
      patterns[60119] = 29'b1_110101011010_111_1_110101011010;
      patterns[60120] = 29'b1_110101011011_000_1_110101011011;
      patterns[60121] = 29'b1_110101011011_001_1_011011110101;
      patterns[60122] = 29'b1_110101011011_010_1_101010110111;
      patterns[60123] = 29'b1_110101011011_011_1_010101101111;
      patterns[60124] = 29'b1_110101011011_100_1_111010101101;
      patterns[60125] = 29'b1_110101011011_101_1_111101010110;
      patterns[60126] = 29'b1_110101011011_110_1_110101011011;
      patterns[60127] = 29'b1_110101011011_111_1_110101011011;
      patterns[60128] = 29'b1_110101011100_000_1_110101011100;
      patterns[60129] = 29'b1_110101011100_001_1_011100110101;
      patterns[60130] = 29'b1_110101011100_010_1_101010111001;
      patterns[60131] = 29'b1_110101011100_011_1_010101110011;
      patterns[60132] = 29'b1_110101011100_100_0_111010101110;
      patterns[60133] = 29'b1_110101011100_101_0_011101010111;
      patterns[60134] = 29'b1_110101011100_110_1_110101011100;
      patterns[60135] = 29'b1_110101011100_111_1_110101011100;
      patterns[60136] = 29'b1_110101011101_000_1_110101011101;
      patterns[60137] = 29'b1_110101011101_001_1_011101110101;
      patterns[60138] = 29'b1_110101011101_010_1_101010111011;
      patterns[60139] = 29'b1_110101011101_011_1_010101110111;
      patterns[60140] = 29'b1_110101011101_100_1_111010101110;
      patterns[60141] = 29'b1_110101011101_101_0_111101010111;
      patterns[60142] = 29'b1_110101011101_110_1_110101011101;
      patterns[60143] = 29'b1_110101011101_111_1_110101011101;
      patterns[60144] = 29'b1_110101011110_000_1_110101011110;
      patterns[60145] = 29'b1_110101011110_001_1_011110110101;
      patterns[60146] = 29'b1_110101011110_010_1_101010111101;
      patterns[60147] = 29'b1_110101011110_011_1_010101111011;
      patterns[60148] = 29'b1_110101011110_100_0_111010101111;
      patterns[60149] = 29'b1_110101011110_101_1_011101010111;
      patterns[60150] = 29'b1_110101011110_110_1_110101011110;
      patterns[60151] = 29'b1_110101011110_111_1_110101011110;
      patterns[60152] = 29'b1_110101011111_000_1_110101011111;
      patterns[60153] = 29'b1_110101011111_001_1_011111110101;
      patterns[60154] = 29'b1_110101011111_010_1_101010111111;
      patterns[60155] = 29'b1_110101011111_011_1_010101111111;
      patterns[60156] = 29'b1_110101011111_100_1_111010101111;
      patterns[60157] = 29'b1_110101011111_101_1_111101010111;
      patterns[60158] = 29'b1_110101011111_110_1_110101011111;
      patterns[60159] = 29'b1_110101011111_111_1_110101011111;
      patterns[60160] = 29'b1_110101100000_000_1_110101100000;
      patterns[60161] = 29'b1_110101100000_001_1_100000110101;
      patterns[60162] = 29'b1_110101100000_010_1_101011000001;
      patterns[60163] = 29'b1_110101100000_011_1_010110000011;
      patterns[60164] = 29'b1_110101100000_100_0_111010110000;
      patterns[60165] = 29'b1_110101100000_101_0_011101011000;
      patterns[60166] = 29'b1_110101100000_110_1_110101100000;
      patterns[60167] = 29'b1_110101100000_111_1_110101100000;
      patterns[60168] = 29'b1_110101100001_000_1_110101100001;
      patterns[60169] = 29'b1_110101100001_001_1_100001110101;
      patterns[60170] = 29'b1_110101100001_010_1_101011000011;
      patterns[60171] = 29'b1_110101100001_011_1_010110000111;
      patterns[60172] = 29'b1_110101100001_100_1_111010110000;
      patterns[60173] = 29'b1_110101100001_101_0_111101011000;
      patterns[60174] = 29'b1_110101100001_110_1_110101100001;
      patterns[60175] = 29'b1_110101100001_111_1_110101100001;
      patterns[60176] = 29'b1_110101100010_000_1_110101100010;
      patterns[60177] = 29'b1_110101100010_001_1_100010110101;
      patterns[60178] = 29'b1_110101100010_010_1_101011000101;
      patterns[60179] = 29'b1_110101100010_011_1_010110001011;
      patterns[60180] = 29'b1_110101100010_100_0_111010110001;
      patterns[60181] = 29'b1_110101100010_101_1_011101011000;
      patterns[60182] = 29'b1_110101100010_110_1_110101100010;
      patterns[60183] = 29'b1_110101100010_111_1_110101100010;
      patterns[60184] = 29'b1_110101100011_000_1_110101100011;
      patterns[60185] = 29'b1_110101100011_001_1_100011110101;
      patterns[60186] = 29'b1_110101100011_010_1_101011000111;
      patterns[60187] = 29'b1_110101100011_011_1_010110001111;
      patterns[60188] = 29'b1_110101100011_100_1_111010110001;
      patterns[60189] = 29'b1_110101100011_101_1_111101011000;
      patterns[60190] = 29'b1_110101100011_110_1_110101100011;
      patterns[60191] = 29'b1_110101100011_111_1_110101100011;
      patterns[60192] = 29'b1_110101100100_000_1_110101100100;
      patterns[60193] = 29'b1_110101100100_001_1_100100110101;
      patterns[60194] = 29'b1_110101100100_010_1_101011001001;
      patterns[60195] = 29'b1_110101100100_011_1_010110010011;
      patterns[60196] = 29'b1_110101100100_100_0_111010110010;
      patterns[60197] = 29'b1_110101100100_101_0_011101011001;
      patterns[60198] = 29'b1_110101100100_110_1_110101100100;
      patterns[60199] = 29'b1_110101100100_111_1_110101100100;
      patterns[60200] = 29'b1_110101100101_000_1_110101100101;
      patterns[60201] = 29'b1_110101100101_001_1_100101110101;
      patterns[60202] = 29'b1_110101100101_010_1_101011001011;
      patterns[60203] = 29'b1_110101100101_011_1_010110010111;
      patterns[60204] = 29'b1_110101100101_100_1_111010110010;
      patterns[60205] = 29'b1_110101100101_101_0_111101011001;
      patterns[60206] = 29'b1_110101100101_110_1_110101100101;
      patterns[60207] = 29'b1_110101100101_111_1_110101100101;
      patterns[60208] = 29'b1_110101100110_000_1_110101100110;
      patterns[60209] = 29'b1_110101100110_001_1_100110110101;
      patterns[60210] = 29'b1_110101100110_010_1_101011001101;
      patterns[60211] = 29'b1_110101100110_011_1_010110011011;
      patterns[60212] = 29'b1_110101100110_100_0_111010110011;
      patterns[60213] = 29'b1_110101100110_101_1_011101011001;
      patterns[60214] = 29'b1_110101100110_110_1_110101100110;
      patterns[60215] = 29'b1_110101100110_111_1_110101100110;
      patterns[60216] = 29'b1_110101100111_000_1_110101100111;
      patterns[60217] = 29'b1_110101100111_001_1_100111110101;
      patterns[60218] = 29'b1_110101100111_010_1_101011001111;
      patterns[60219] = 29'b1_110101100111_011_1_010110011111;
      patterns[60220] = 29'b1_110101100111_100_1_111010110011;
      patterns[60221] = 29'b1_110101100111_101_1_111101011001;
      patterns[60222] = 29'b1_110101100111_110_1_110101100111;
      patterns[60223] = 29'b1_110101100111_111_1_110101100111;
      patterns[60224] = 29'b1_110101101000_000_1_110101101000;
      patterns[60225] = 29'b1_110101101000_001_1_101000110101;
      patterns[60226] = 29'b1_110101101000_010_1_101011010001;
      patterns[60227] = 29'b1_110101101000_011_1_010110100011;
      patterns[60228] = 29'b1_110101101000_100_0_111010110100;
      patterns[60229] = 29'b1_110101101000_101_0_011101011010;
      patterns[60230] = 29'b1_110101101000_110_1_110101101000;
      patterns[60231] = 29'b1_110101101000_111_1_110101101000;
      patterns[60232] = 29'b1_110101101001_000_1_110101101001;
      patterns[60233] = 29'b1_110101101001_001_1_101001110101;
      patterns[60234] = 29'b1_110101101001_010_1_101011010011;
      patterns[60235] = 29'b1_110101101001_011_1_010110100111;
      patterns[60236] = 29'b1_110101101001_100_1_111010110100;
      patterns[60237] = 29'b1_110101101001_101_0_111101011010;
      patterns[60238] = 29'b1_110101101001_110_1_110101101001;
      patterns[60239] = 29'b1_110101101001_111_1_110101101001;
      patterns[60240] = 29'b1_110101101010_000_1_110101101010;
      patterns[60241] = 29'b1_110101101010_001_1_101010110101;
      patterns[60242] = 29'b1_110101101010_010_1_101011010101;
      patterns[60243] = 29'b1_110101101010_011_1_010110101011;
      patterns[60244] = 29'b1_110101101010_100_0_111010110101;
      patterns[60245] = 29'b1_110101101010_101_1_011101011010;
      patterns[60246] = 29'b1_110101101010_110_1_110101101010;
      patterns[60247] = 29'b1_110101101010_111_1_110101101010;
      patterns[60248] = 29'b1_110101101011_000_1_110101101011;
      patterns[60249] = 29'b1_110101101011_001_1_101011110101;
      patterns[60250] = 29'b1_110101101011_010_1_101011010111;
      patterns[60251] = 29'b1_110101101011_011_1_010110101111;
      patterns[60252] = 29'b1_110101101011_100_1_111010110101;
      patterns[60253] = 29'b1_110101101011_101_1_111101011010;
      patterns[60254] = 29'b1_110101101011_110_1_110101101011;
      patterns[60255] = 29'b1_110101101011_111_1_110101101011;
      patterns[60256] = 29'b1_110101101100_000_1_110101101100;
      patterns[60257] = 29'b1_110101101100_001_1_101100110101;
      patterns[60258] = 29'b1_110101101100_010_1_101011011001;
      patterns[60259] = 29'b1_110101101100_011_1_010110110011;
      patterns[60260] = 29'b1_110101101100_100_0_111010110110;
      patterns[60261] = 29'b1_110101101100_101_0_011101011011;
      patterns[60262] = 29'b1_110101101100_110_1_110101101100;
      patterns[60263] = 29'b1_110101101100_111_1_110101101100;
      patterns[60264] = 29'b1_110101101101_000_1_110101101101;
      patterns[60265] = 29'b1_110101101101_001_1_101101110101;
      patterns[60266] = 29'b1_110101101101_010_1_101011011011;
      patterns[60267] = 29'b1_110101101101_011_1_010110110111;
      patterns[60268] = 29'b1_110101101101_100_1_111010110110;
      patterns[60269] = 29'b1_110101101101_101_0_111101011011;
      patterns[60270] = 29'b1_110101101101_110_1_110101101101;
      patterns[60271] = 29'b1_110101101101_111_1_110101101101;
      patterns[60272] = 29'b1_110101101110_000_1_110101101110;
      patterns[60273] = 29'b1_110101101110_001_1_101110110101;
      patterns[60274] = 29'b1_110101101110_010_1_101011011101;
      patterns[60275] = 29'b1_110101101110_011_1_010110111011;
      patterns[60276] = 29'b1_110101101110_100_0_111010110111;
      patterns[60277] = 29'b1_110101101110_101_1_011101011011;
      patterns[60278] = 29'b1_110101101110_110_1_110101101110;
      patterns[60279] = 29'b1_110101101110_111_1_110101101110;
      patterns[60280] = 29'b1_110101101111_000_1_110101101111;
      patterns[60281] = 29'b1_110101101111_001_1_101111110101;
      patterns[60282] = 29'b1_110101101111_010_1_101011011111;
      patterns[60283] = 29'b1_110101101111_011_1_010110111111;
      patterns[60284] = 29'b1_110101101111_100_1_111010110111;
      patterns[60285] = 29'b1_110101101111_101_1_111101011011;
      patterns[60286] = 29'b1_110101101111_110_1_110101101111;
      patterns[60287] = 29'b1_110101101111_111_1_110101101111;
      patterns[60288] = 29'b1_110101110000_000_1_110101110000;
      patterns[60289] = 29'b1_110101110000_001_1_110000110101;
      patterns[60290] = 29'b1_110101110000_010_1_101011100001;
      patterns[60291] = 29'b1_110101110000_011_1_010111000011;
      patterns[60292] = 29'b1_110101110000_100_0_111010111000;
      patterns[60293] = 29'b1_110101110000_101_0_011101011100;
      patterns[60294] = 29'b1_110101110000_110_1_110101110000;
      patterns[60295] = 29'b1_110101110000_111_1_110101110000;
      patterns[60296] = 29'b1_110101110001_000_1_110101110001;
      patterns[60297] = 29'b1_110101110001_001_1_110001110101;
      patterns[60298] = 29'b1_110101110001_010_1_101011100011;
      patterns[60299] = 29'b1_110101110001_011_1_010111000111;
      patterns[60300] = 29'b1_110101110001_100_1_111010111000;
      patterns[60301] = 29'b1_110101110001_101_0_111101011100;
      patterns[60302] = 29'b1_110101110001_110_1_110101110001;
      patterns[60303] = 29'b1_110101110001_111_1_110101110001;
      patterns[60304] = 29'b1_110101110010_000_1_110101110010;
      patterns[60305] = 29'b1_110101110010_001_1_110010110101;
      patterns[60306] = 29'b1_110101110010_010_1_101011100101;
      patterns[60307] = 29'b1_110101110010_011_1_010111001011;
      patterns[60308] = 29'b1_110101110010_100_0_111010111001;
      patterns[60309] = 29'b1_110101110010_101_1_011101011100;
      patterns[60310] = 29'b1_110101110010_110_1_110101110010;
      patterns[60311] = 29'b1_110101110010_111_1_110101110010;
      patterns[60312] = 29'b1_110101110011_000_1_110101110011;
      patterns[60313] = 29'b1_110101110011_001_1_110011110101;
      patterns[60314] = 29'b1_110101110011_010_1_101011100111;
      patterns[60315] = 29'b1_110101110011_011_1_010111001111;
      patterns[60316] = 29'b1_110101110011_100_1_111010111001;
      patterns[60317] = 29'b1_110101110011_101_1_111101011100;
      patterns[60318] = 29'b1_110101110011_110_1_110101110011;
      patterns[60319] = 29'b1_110101110011_111_1_110101110011;
      patterns[60320] = 29'b1_110101110100_000_1_110101110100;
      patterns[60321] = 29'b1_110101110100_001_1_110100110101;
      patterns[60322] = 29'b1_110101110100_010_1_101011101001;
      patterns[60323] = 29'b1_110101110100_011_1_010111010011;
      patterns[60324] = 29'b1_110101110100_100_0_111010111010;
      patterns[60325] = 29'b1_110101110100_101_0_011101011101;
      patterns[60326] = 29'b1_110101110100_110_1_110101110100;
      patterns[60327] = 29'b1_110101110100_111_1_110101110100;
      patterns[60328] = 29'b1_110101110101_000_1_110101110101;
      patterns[60329] = 29'b1_110101110101_001_1_110101110101;
      patterns[60330] = 29'b1_110101110101_010_1_101011101011;
      patterns[60331] = 29'b1_110101110101_011_1_010111010111;
      patterns[60332] = 29'b1_110101110101_100_1_111010111010;
      patterns[60333] = 29'b1_110101110101_101_0_111101011101;
      patterns[60334] = 29'b1_110101110101_110_1_110101110101;
      patterns[60335] = 29'b1_110101110101_111_1_110101110101;
      patterns[60336] = 29'b1_110101110110_000_1_110101110110;
      patterns[60337] = 29'b1_110101110110_001_1_110110110101;
      patterns[60338] = 29'b1_110101110110_010_1_101011101101;
      patterns[60339] = 29'b1_110101110110_011_1_010111011011;
      patterns[60340] = 29'b1_110101110110_100_0_111010111011;
      patterns[60341] = 29'b1_110101110110_101_1_011101011101;
      patterns[60342] = 29'b1_110101110110_110_1_110101110110;
      patterns[60343] = 29'b1_110101110110_111_1_110101110110;
      patterns[60344] = 29'b1_110101110111_000_1_110101110111;
      patterns[60345] = 29'b1_110101110111_001_1_110111110101;
      patterns[60346] = 29'b1_110101110111_010_1_101011101111;
      patterns[60347] = 29'b1_110101110111_011_1_010111011111;
      patterns[60348] = 29'b1_110101110111_100_1_111010111011;
      patterns[60349] = 29'b1_110101110111_101_1_111101011101;
      patterns[60350] = 29'b1_110101110111_110_1_110101110111;
      patterns[60351] = 29'b1_110101110111_111_1_110101110111;
      patterns[60352] = 29'b1_110101111000_000_1_110101111000;
      patterns[60353] = 29'b1_110101111000_001_1_111000110101;
      patterns[60354] = 29'b1_110101111000_010_1_101011110001;
      patterns[60355] = 29'b1_110101111000_011_1_010111100011;
      patterns[60356] = 29'b1_110101111000_100_0_111010111100;
      patterns[60357] = 29'b1_110101111000_101_0_011101011110;
      patterns[60358] = 29'b1_110101111000_110_1_110101111000;
      patterns[60359] = 29'b1_110101111000_111_1_110101111000;
      patterns[60360] = 29'b1_110101111001_000_1_110101111001;
      patterns[60361] = 29'b1_110101111001_001_1_111001110101;
      patterns[60362] = 29'b1_110101111001_010_1_101011110011;
      patterns[60363] = 29'b1_110101111001_011_1_010111100111;
      patterns[60364] = 29'b1_110101111001_100_1_111010111100;
      patterns[60365] = 29'b1_110101111001_101_0_111101011110;
      patterns[60366] = 29'b1_110101111001_110_1_110101111001;
      patterns[60367] = 29'b1_110101111001_111_1_110101111001;
      patterns[60368] = 29'b1_110101111010_000_1_110101111010;
      patterns[60369] = 29'b1_110101111010_001_1_111010110101;
      patterns[60370] = 29'b1_110101111010_010_1_101011110101;
      patterns[60371] = 29'b1_110101111010_011_1_010111101011;
      patterns[60372] = 29'b1_110101111010_100_0_111010111101;
      patterns[60373] = 29'b1_110101111010_101_1_011101011110;
      patterns[60374] = 29'b1_110101111010_110_1_110101111010;
      patterns[60375] = 29'b1_110101111010_111_1_110101111010;
      patterns[60376] = 29'b1_110101111011_000_1_110101111011;
      patterns[60377] = 29'b1_110101111011_001_1_111011110101;
      patterns[60378] = 29'b1_110101111011_010_1_101011110111;
      patterns[60379] = 29'b1_110101111011_011_1_010111101111;
      patterns[60380] = 29'b1_110101111011_100_1_111010111101;
      patterns[60381] = 29'b1_110101111011_101_1_111101011110;
      patterns[60382] = 29'b1_110101111011_110_1_110101111011;
      patterns[60383] = 29'b1_110101111011_111_1_110101111011;
      patterns[60384] = 29'b1_110101111100_000_1_110101111100;
      patterns[60385] = 29'b1_110101111100_001_1_111100110101;
      patterns[60386] = 29'b1_110101111100_010_1_101011111001;
      patterns[60387] = 29'b1_110101111100_011_1_010111110011;
      patterns[60388] = 29'b1_110101111100_100_0_111010111110;
      patterns[60389] = 29'b1_110101111100_101_0_011101011111;
      patterns[60390] = 29'b1_110101111100_110_1_110101111100;
      patterns[60391] = 29'b1_110101111100_111_1_110101111100;
      patterns[60392] = 29'b1_110101111101_000_1_110101111101;
      patterns[60393] = 29'b1_110101111101_001_1_111101110101;
      patterns[60394] = 29'b1_110101111101_010_1_101011111011;
      patterns[60395] = 29'b1_110101111101_011_1_010111110111;
      patterns[60396] = 29'b1_110101111101_100_1_111010111110;
      patterns[60397] = 29'b1_110101111101_101_0_111101011111;
      patterns[60398] = 29'b1_110101111101_110_1_110101111101;
      patterns[60399] = 29'b1_110101111101_111_1_110101111101;
      patterns[60400] = 29'b1_110101111110_000_1_110101111110;
      patterns[60401] = 29'b1_110101111110_001_1_111110110101;
      patterns[60402] = 29'b1_110101111110_010_1_101011111101;
      patterns[60403] = 29'b1_110101111110_011_1_010111111011;
      patterns[60404] = 29'b1_110101111110_100_0_111010111111;
      patterns[60405] = 29'b1_110101111110_101_1_011101011111;
      patterns[60406] = 29'b1_110101111110_110_1_110101111110;
      patterns[60407] = 29'b1_110101111110_111_1_110101111110;
      patterns[60408] = 29'b1_110101111111_000_1_110101111111;
      patterns[60409] = 29'b1_110101111111_001_1_111111110101;
      patterns[60410] = 29'b1_110101111111_010_1_101011111111;
      patterns[60411] = 29'b1_110101111111_011_1_010111111111;
      patterns[60412] = 29'b1_110101111111_100_1_111010111111;
      patterns[60413] = 29'b1_110101111111_101_1_111101011111;
      patterns[60414] = 29'b1_110101111111_110_1_110101111111;
      patterns[60415] = 29'b1_110101111111_111_1_110101111111;
      patterns[60416] = 29'b1_110110000000_000_1_110110000000;
      patterns[60417] = 29'b1_110110000000_001_1_000000110110;
      patterns[60418] = 29'b1_110110000000_010_1_101100000001;
      patterns[60419] = 29'b1_110110000000_011_1_011000000011;
      patterns[60420] = 29'b1_110110000000_100_0_111011000000;
      patterns[60421] = 29'b1_110110000000_101_0_011101100000;
      patterns[60422] = 29'b1_110110000000_110_1_110110000000;
      patterns[60423] = 29'b1_110110000000_111_1_110110000000;
      patterns[60424] = 29'b1_110110000001_000_1_110110000001;
      patterns[60425] = 29'b1_110110000001_001_1_000001110110;
      patterns[60426] = 29'b1_110110000001_010_1_101100000011;
      patterns[60427] = 29'b1_110110000001_011_1_011000000111;
      patterns[60428] = 29'b1_110110000001_100_1_111011000000;
      patterns[60429] = 29'b1_110110000001_101_0_111101100000;
      patterns[60430] = 29'b1_110110000001_110_1_110110000001;
      patterns[60431] = 29'b1_110110000001_111_1_110110000001;
      patterns[60432] = 29'b1_110110000010_000_1_110110000010;
      patterns[60433] = 29'b1_110110000010_001_1_000010110110;
      patterns[60434] = 29'b1_110110000010_010_1_101100000101;
      patterns[60435] = 29'b1_110110000010_011_1_011000001011;
      patterns[60436] = 29'b1_110110000010_100_0_111011000001;
      patterns[60437] = 29'b1_110110000010_101_1_011101100000;
      patterns[60438] = 29'b1_110110000010_110_1_110110000010;
      patterns[60439] = 29'b1_110110000010_111_1_110110000010;
      patterns[60440] = 29'b1_110110000011_000_1_110110000011;
      patterns[60441] = 29'b1_110110000011_001_1_000011110110;
      patterns[60442] = 29'b1_110110000011_010_1_101100000111;
      patterns[60443] = 29'b1_110110000011_011_1_011000001111;
      patterns[60444] = 29'b1_110110000011_100_1_111011000001;
      patterns[60445] = 29'b1_110110000011_101_1_111101100000;
      patterns[60446] = 29'b1_110110000011_110_1_110110000011;
      patterns[60447] = 29'b1_110110000011_111_1_110110000011;
      patterns[60448] = 29'b1_110110000100_000_1_110110000100;
      patterns[60449] = 29'b1_110110000100_001_1_000100110110;
      patterns[60450] = 29'b1_110110000100_010_1_101100001001;
      patterns[60451] = 29'b1_110110000100_011_1_011000010011;
      patterns[60452] = 29'b1_110110000100_100_0_111011000010;
      patterns[60453] = 29'b1_110110000100_101_0_011101100001;
      patterns[60454] = 29'b1_110110000100_110_1_110110000100;
      patterns[60455] = 29'b1_110110000100_111_1_110110000100;
      patterns[60456] = 29'b1_110110000101_000_1_110110000101;
      patterns[60457] = 29'b1_110110000101_001_1_000101110110;
      patterns[60458] = 29'b1_110110000101_010_1_101100001011;
      patterns[60459] = 29'b1_110110000101_011_1_011000010111;
      patterns[60460] = 29'b1_110110000101_100_1_111011000010;
      patterns[60461] = 29'b1_110110000101_101_0_111101100001;
      patterns[60462] = 29'b1_110110000101_110_1_110110000101;
      patterns[60463] = 29'b1_110110000101_111_1_110110000101;
      patterns[60464] = 29'b1_110110000110_000_1_110110000110;
      patterns[60465] = 29'b1_110110000110_001_1_000110110110;
      patterns[60466] = 29'b1_110110000110_010_1_101100001101;
      patterns[60467] = 29'b1_110110000110_011_1_011000011011;
      patterns[60468] = 29'b1_110110000110_100_0_111011000011;
      patterns[60469] = 29'b1_110110000110_101_1_011101100001;
      patterns[60470] = 29'b1_110110000110_110_1_110110000110;
      patterns[60471] = 29'b1_110110000110_111_1_110110000110;
      patterns[60472] = 29'b1_110110000111_000_1_110110000111;
      patterns[60473] = 29'b1_110110000111_001_1_000111110110;
      patterns[60474] = 29'b1_110110000111_010_1_101100001111;
      patterns[60475] = 29'b1_110110000111_011_1_011000011111;
      patterns[60476] = 29'b1_110110000111_100_1_111011000011;
      patterns[60477] = 29'b1_110110000111_101_1_111101100001;
      patterns[60478] = 29'b1_110110000111_110_1_110110000111;
      patterns[60479] = 29'b1_110110000111_111_1_110110000111;
      patterns[60480] = 29'b1_110110001000_000_1_110110001000;
      patterns[60481] = 29'b1_110110001000_001_1_001000110110;
      patterns[60482] = 29'b1_110110001000_010_1_101100010001;
      patterns[60483] = 29'b1_110110001000_011_1_011000100011;
      patterns[60484] = 29'b1_110110001000_100_0_111011000100;
      patterns[60485] = 29'b1_110110001000_101_0_011101100010;
      patterns[60486] = 29'b1_110110001000_110_1_110110001000;
      patterns[60487] = 29'b1_110110001000_111_1_110110001000;
      patterns[60488] = 29'b1_110110001001_000_1_110110001001;
      patterns[60489] = 29'b1_110110001001_001_1_001001110110;
      patterns[60490] = 29'b1_110110001001_010_1_101100010011;
      patterns[60491] = 29'b1_110110001001_011_1_011000100111;
      patterns[60492] = 29'b1_110110001001_100_1_111011000100;
      patterns[60493] = 29'b1_110110001001_101_0_111101100010;
      patterns[60494] = 29'b1_110110001001_110_1_110110001001;
      patterns[60495] = 29'b1_110110001001_111_1_110110001001;
      patterns[60496] = 29'b1_110110001010_000_1_110110001010;
      patterns[60497] = 29'b1_110110001010_001_1_001010110110;
      patterns[60498] = 29'b1_110110001010_010_1_101100010101;
      patterns[60499] = 29'b1_110110001010_011_1_011000101011;
      patterns[60500] = 29'b1_110110001010_100_0_111011000101;
      patterns[60501] = 29'b1_110110001010_101_1_011101100010;
      patterns[60502] = 29'b1_110110001010_110_1_110110001010;
      patterns[60503] = 29'b1_110110001010_111_1_110110001010;
      patterns[60504] = 29'b1_110110001011_000_1_110110001011;
      patterns[60505] = 29'b1_110110001011_001_1_001011110110;
      patterns[60506] = 29'b1_110110001011_010_1_101100010111;
      patterns[60507] = 29'b1_110110001011_011_1_011000101111;
      patterns[60508] = 29'b1_110110001011_100_1_111011000101;
      patterns[60509] = 29'b1_110110001011_101_1_111101100010;
      patterns[60510] = 29'b1_110110001011_110_1_110110001011;
      patterns[60511] = 29'b1_110110001011_111_1_110110001011;
      patterns[60512] = 29'b1_110110001100_000_1_110110001100;
      patterns[60513] = 29'b1_110110001100_001_1_001100110110;
      patterns[60514] = 29'b1_110110001100_010_1_101100011001;
      patterns[60515] = 29'b1_110110001100_011_1_011000110011;
      patterns[60516] = 29'b1_110110001100_100_0_111011000110;
      patterns[60517] = 29'b1_110110001100_101_0_011101100011;
      patterns[60518] = 29'b1_110110001100_110_1_110110001100;
      patterns[60519] = 29'b1_110110001100_111_1_110110001100;
      patterns[60520] = 29'b1_110110001101_000_1_110110001101;
      patterns[60521] = 29'b1_110110001101_001_1_001101110110;
      patterns[60522] = 29'b1_110110001101_010_1_101100011011;
      patterns[60523] = 29'b1_110110001101_011_1_011000110111;
      patterns[60524] = 29'b1_110110001101_100_1_111011000110;
      patterns[60525] = 29'b1_110110001101_101_0_111101100011;
      patterns[60526] = 29'b1_110110001101_110_1_110110001101;
      patterns[60527] = 29'b1_110110001101_111_1_110110001101;
      patterns[60528] = 29'b1_110110001110_000_1_110110001110;
      patterns[60529] = 29'b1_110110001110_001_1_001110110110;
      patterns[60530] = 29'b1_110110001110_010_1_101100011101;
      patterns[60531] = 29'b1_110110001110_011_1_011000111011;
      patterns[60532] = 29'b1_110110001110_100_0_111011000111;
      patterns[60533] = 29'b1_110110001110_101_1_011101100011;
      patterns[60534] = 29'b1_110110001110_110_1_110110001110;
      patterns[60535] = 29'b1_110110001110_111_1_110110001110;
      patterns[60536] = 29'b1_110110001111_000_1_110110001111;
      patterns[60537] = 29'b1_110110001111_001_1_001111110110;
      patterns[60538] = 29'b1_110110001111_010_1_101100011111;
      patterns[60539] = 29'b1_110110001111_011_1_011000111111;
      patterns[60540] = 29'b1_110110001111_100_1_111011000111;
      patterns[60541] = 29'b1_110110001111_101_1_111101100011;
      patterns[60542] = 29'b1_110110001111_110_1_110110001111;
      patterns[60543] = 29'b1_110110001111_111_1_110110001111;
      patterns[60544] = 29'b1_110110010000_000_1_110110010000;
      patterns[60545] = 29'b1_110110010000_001_1_010000110110;
      patterns[60546] = 29'b1_110110010000_010_1_101100100001;
      patterns[60547] = 29'b1_110110010000_011_1_011001000011;
      patterns[60548] = 29'b1_110110010000_100_0_111011001000;
      patterns[60549] = 29'b1_110110010000_101_0_011101100100;
      patterns[60550] = 29'b1_110110010000_110_1_110110010000;
      patterns[60551] = 29'b1_110110010000_111_1_110110010000;
      patterns[60552] = 29'b1_110110010001_000_1_110110010001;
      patterns[60553] = 29'b1_110110010001_001_1_010001110110;
      patterns[60554] = 29'b1_110110010001_010_1_101100100011;
      patterns[60555] = 29'b1_110110010001_011_1_011001000111;
      patterns[60556] = 29'b1_110110010001_100_1_111011001000;
      patterns[60557] = 29'b1_110110010001_101_0_111101100100;
      patterns[60558] = 29'b1_110110010001_110_1_110110010001;
      patterns[60559] = 29'b1_110110010001_111_1_110110010001;
      patterns[60560] = 29'b1_110110010010_000_1_110110010010;
      patterns[60561] = 29'b1_110110010010_001_1_010010110110;
      patterns[60562] = 29'b1_110110010010_010_1_101100100101;
      patterns[60563] = 29'b1_110110010010_011_1_011001001011;
      patterns[60564] = 29'b1_110110010010_100_0_111011001001;
      patterns[60565] = 29'b1_110110010010_101_1_011101100100;
      patterns[60566] = 29'b1_110110010010_110_1_110110010010;
      patterns[60567] = 29'b1_110110010010_111_1_110110010010;
      patterns[60568] = 29'b1_110110010011_000_1_110110010011;
      patterns[60569] = 29'b1_110110010011_001_1_010011110110;
      patterns[60570] = 29'b1_110110010011_010_1_101100100111;
      patterns[60571] = 29'b1_110110010011_011_1_011001001111;
      patterns[60572] = 29'b1_110110010011_100_1_111011001001;
      patterns[60573] = 29'b1_110110010011_101_1_111101100100;
      patterns[60574] = 29'b1_110110010011_110_1_110110010011;
      patterns[60575] = 29'b1_110110010011_111_1_110110010011;
      patterns[60576] = 29'b1_110110010100_000_1_110110010100;
      patterns[60577] = 29'b1_110110010100_001_1_010100110110;
      patterns[60578] = 29'b1_110110010100_010_1_101100101001;
      patterns[60579] = 29'b1_110110010100_011_1_011001010011;
      patterns[60580] = 29'b1_110110010100_100_0_111011001010;
      patterns[60581] = 29'b1_110110010100_101_0_011101100101;
      patterns[60582] = 29'b1_110110010100_110_1_110110010100;
      patterns[60583] = 29'b1_110110010100_111_1_110110010100;
      patterns[60584] = 29'b1_110110010101_000_1_110110010101;
      patterns[60585] = 29'b1_110110010101_001_1_010101110110;
      patterns[60586] = 29'b1_110110010101_010_1_101100101011;
      patterns[60587] = 29'b1_110110010101_011_1_011001010111;
      patterns[60588] = 29'b1_110110010101_100_1_111011001010;
      patterns[60589] = 29'b1_110110010101_101_0_111101100101;
      patterns[60590] = 29'b1_110110010101_110_1_110110010101;
      patterns[60591] = 29'b1_110110010101_111_1_110110010101;
      patterns[60592] = 29'b1_110110010110_000_1_110110010110;
      patterns[60593] = 29'b1_110110010110_001_1_010110110110;
      patterns[60594] = 29'b1_110110010110_010_1_101100101101;
      patterns[60595] = 29'b1_110110010110_011_1_011001011011;
      patterns[60596] = 29'b1_110110010110_100_0_111011001011;
      patterns[60597] = 29'b1_110110010110_101_1_011101100101;
      patterns[60598] = 29'b1_110110010110_110_1_110110010110;
      patterns[60599] = 29'b1_110110010110_111_1_110110010110;
      patterns[60600] = 29'b1_110110010111_000_1_110110010111;
      patterns[60601] = 29'b1_110110010111_001_1_010111110110;
      patterns[60602] = 29'b1_110110010111_010_1_101100101111;
      patterns[60603] = 29'b1_110110010111_011_1_011001011111;
      patterns[60604] = 29'b1_110110010111_100_1_111011001011;
      patterns[60605] = 29'b1_110110010111_101_1_111101100101;
      patterns[60606] = 29'b1_110110010111_110_1_110110010111;
      patterns[60607] = 29'b1_110110010111_111_1_110110010111;
      patterns[60608] = 29'b1_110110011000_000_1_110110011000;
      patterns[60609] = 29'b1_110110011000_001_1_011000110110;
      patterns[60610] = 29'b1_110110011000_010_1_101100110001;
      patterns[60611] = 29'b1_110110011000_011_1_011001100011;
      patterns[60612] = 29'b1_110110011000_100_0_111011001100;
      patterns[60613] = 29'b1_110110011000_101_0_011101100110;
      patterns[60614] = 29'b1_110110011000_110_1_110110011000;
      patterns[60615] = 29'b1_110110011000_111_1_110110011000;
      patterns[60616] = 29'b1_110110011001_000_1_110110011001;
      patterns[60617] = 29'b1_110110011001_001_1_011001110110;
      patterns[60618] = 29'b1_110110011001_010_1_101100110011;
      patterns[60619] = 29'b1_110110011001_011_1_011001100111;
      patterns[60620] = 29'b1_110110011001_100_1_111011001100;
      patterns[60621] = 29'b1_110110011001_101_0_111101100110;
      patterns[60622] = 29'b1_110110011001_110_1_110110011001;
      patterns[60623] = 29'b1_110110011001_111_1_110110011001;
      patterns[60624] = 29'b1_110110011010_000_1_110110011010;
      patterns[60625] = 29'b1_110110011010_001_1_011010110110;
      patterns[60626] = 29'b1_110110011010_010_1_101100110101;
      patterns[60627] = 29'b1_110110011010_011_1_011001101011;
      patterns[60628] = 29'b1_110110011010_100_0_111011001101;
      patterns[60629] = 29'b1_110110011010_101_1_011101100110;
      patterns[60630] = 29'b1_110110011010_110_1_110110011010;
      patterns[60631] = 29'b1_110110011010_111_1_110110011010;
      patterns[60632] = 29'b1_110110011011_000_1_110110011011;
      patterns[60633] = 29'b1_110110011011_001_1_011011110110;
      patterns[60634] = 29'b1_110110011011_010_1_101100110111;
      patterns[60635] = 29'b1_110110011011_011_1_011001101111;
      patterns[60636] = 29'b1_110110011011_100_1_111011001101;
      patterns[60637] = 29'b1_110110011011_101_1_111101100110;
      patterns[60638] = 29'b1_110110011011_110_1_110110011011;
      patterns[60639] = 29'b1_110110011011_111_1_110110011011;
      patterns[60640] = 29'b1_110110011100_000_1_110110011100;
      patterns[60641] = 29'b1_110110011100_001_1_011100110110;
      patterns[60642] = 29'b1_110110011100_010_1_101100111001;
      patterns[60643] = 29'b1_110110011100_011_1_011001110011;
      patterns[60644] = 29'b1_110110011100_100_0_111011001110;
      patterns[60645] = 29'b1_110110011100_101_0_011101100111;
      patterns[60646] = 29'b1_110110011100_110_1_110110011100;
      patterns[60647] = 29'b1_110110011100_111_1_110110011100;
      patterns[60648] = 29'b1_110110011101_000_1_110110011101;
      patterns[60649] = 29'b1_110110011101_001_1_011101110110;
      patterns[60650] = 29'b1_110110011101_010_1_101100111011;
      patterns[60651] = 29'b1_110110011101_011_1_011001110111;
      patterns[60652] = 29'b1_110110011101_100_1_111011001110;
      patterns[60653] = 29'b1_110110011101_101_0_111101100111;
      patterns[60654] = 29'b1_110110011101_110_1_110110011101;
      patterns[60655] = 29'b1_110110011101_111_1_110110011101;
      patterns[60656] = 29'b1_110110011110_000_1_110110011110;
      patterns[60657] = 29'b1_110110011110_001_1_011110110110;
      patterns[60658] = 29'b1_110110011110_010_1_101100111101;
      patterns[60659] = 29'b1_110110011110_011_1_011001111011;
      patterns[60660] = 29'b1_110110011110_100_0_111011001111;
      patterns[60661] = 29'b1_110110011110_101_1_011101100111;
      patterns[60662] = 29'b1_110110011110_110_1_110110011110;
      patterns[60663] = 29'b1_110110011110_111_1_110110011110;
      patterns[60664] = 29'b1_110110011111_000_1_110110011111;
      patterns[60665] = 29'b1_110110011111_001_1_011111110110;
      patterns[60666] = 29'b1_110110011111_010_1_101100111111;
      patterns[60667] = 29'b1_110110011111_011_1_011001111111;
      patterns[60668] = 29'b1_110110011111_100_1_111011001111;
      patterns[60669] = 29'b1_110110011111_101_1_111101100111;
      patterns[60670] = 29'b1_110110011111_110_1_110110011111;
      patterns[60671] = 29'b1_110110011111_111_1_110110011111;
      patterns[60672] = 29'b1_110110100000_000_1_110110100000;
      patterns[60673] = 29'b1_110110100000_001_1_100000110110;
      patterns[60674] = 29'b1_110110100000_010_1_101101000001;
      patterns[60675] = 29'b1_110110100000_011_1_011010000011;
      patterns[60676] = 29'b1_110110100000_100_0_111011010000;
      patterns[60677] = 29'b1_110110100000_101_0_011101101000;
      patterns[60678] = 29'b1_110110100000_110_1_110110100000;
      patterns[60679] = 29'b1_110110100000_111_1_110110100000;
      patterns[60680] = 29'b1_110110100001_000_1_110110100001;
      patterns[60681] = 29'b1_110110100001_001_1_100001110110;
      patterns[60682] = 29'b1_110110100001_010_1_101101000011;
      patterns[60683] = 29'b1_110110100001_011_1_011010000111;
      patterns[60684] = 29'b1_110110100001_100_1_111011010000;
      patterns[60685] = 29'b1_110110100001_101_0_111101101000;
      patterns[60686] = 29'b1_110110100001_110_1_110110100001;
      patterns[60687] = 29'b1_110110100001_111_1_110110100001;
      patterns[60688] = 29'b1_110110100010_000_1_110110100010;
      patterns[60689] = 29'b1_110110100010_001_1_100010110110;
      patterns[60690] = 29'b1_110110100010_010_1_101101000101;
      patterns[60691] = 29'b1_110110100010_011_1_011010001011;
      patterns[60692] = 29'b1_110110100010_100_0_111011010001;
      patterns[60693] = 29'b1_110110100010_101_1_011101101000;
      patterns[60694] = 29'b1_110110100010_110_1_110110100010;
      patterns[60695] = 29'b1_110110100010_111_1_110110100010;
      patterns[60696] = 29'b1_110110100011_000_1_110110100011;
      patterns[60697] = 29'b1_110110100011_001_1_100011110110;
      patterns[60698] = 29'b1_110110100011_010_1_101101000111;
      patterns[60699] = 29'b1_110110100011_011_1_011010001111;
      patterns[60700] = 29'b1_110110100011_100_1_111011010001;
      patterns[60701] = 29'b1_110110100011_101_1_111101101000;
      patterns[60702] = 29'b1_110110100011_110_1_110110100011;
      patterns[60703] = 29'b1_110110100011_111_1_110110100011;
      patterns[60704] = 29'b1_110110100100_000_1_110110100100;
      patterns[60705] = 29'b1_110110100100_001_1_100100110110;
      patterns[60706] = 29'b1_110110100100_010_1_101101001001;
      patterns[60707] = 29'b1_110110100100_011_1_011010010011;
      patterns[60708] = 29'b1_110110100100_100_0_111011010010;
      patterns[60709] = 29'b1_110110100100_101_0_011101101001;
      patterns[60710] = 29'b1_110110100100_110_1_110110100100;
      patterns[60711] = 29'b1_110110100100_111_1_110110100100;
      patterns[60712] = 29'b1_110110100101_000_1_110110100101;
      patterns[60713] = 29'b1_110110100101_001_1_100101110110;
      patterns[60714] = 29'b1_110110100101_010_1_101101001011;
      patterns[60715] = 29'b1_110110100101_011_1_011010010111;
      patterns[60716] = 29'b1_110110100101_100_1_111011010010;
      patterns[60717] = 29'b1_110110100101_101_0_111101101001;
      patterns[60718] = 29'b1_110110100101_110_1_110110100101;
      patterns[60719] = 29'b1_110110100101_111_1_110110100101;
      patterns[60720] = 29'b1_110110100110_000_1_110110100110;
      patterns[60721] = 29'b1_110110100110_001_1_100110110110;
      patterns[60722] = 29'b1_110110100110_010_1_101101001101;
      patterns[60723] = 29'b1_110110100110_011_1_011010011011;
      patterns[60724] = 29'b1_110110100110_100_0_111011010011;
      patterns[60725] = 29'b1_110110100110_101_1_011101101001;
      patterns[60726] = 29'b1_110110100110_110_1_110110100110;
      patterns[60727] = 29'b1_110110100110_111_1_110110100110;
      patterns[60728] = 29'b1_110110100111_000_1_110110100111;
      patterns[60729] = 29'b1_110110100111_001_1_100111110110;
      patterns[60730] = 29'b1_110110100111_010_1_101101001111;
      patterns[60731] = 29'b1_110110100111_011_1_011010011111;
      patterns[60732] = 29'b1_110110100111_100_1_111011010011;
      patterns[60733] = 29'b1_110110100111_101_1_111101101001;
      patterns[60734] = 29'b1_110110100111_110_1_110110100111;
      patterns[60735] = 29'b1_110110100111_111_1_110110100111;
      patterns[60736] = 29'b1_110110101000_000_1_110110101000;
      patterns[60737] = 29'b1_110110101000_001_1_101000110110;
      patterns[60738] = 29'b1_110110101000_010_1_101101010001;
      patterns[60739] = 29'b1_110110101000_011_1_011010100011;
      patterns[60740] = 29'b1_110110101000_100_0_111011010100;
      patterns[60741] = 29'b1_110110101000_101_0_011101101010;
      patterns[60742] = 29'b1_110110101000_110_1_110110101000;
      patterns[60743] = 29'b1_110110101000_111_1_110110101000;
      patterns[60744] = 29'b1_110110101001_000_1_110110101001;
      patterns[60745] = 29'b1_110110101001_001_1_101001110110;
      patterns[60746] = 29'b1_110110101001_010_1_101101010011;
      patterns[60747] = 29'b1_110110101001_011_1_011010100111;
      patterns[60748] = 29'b1_110110101001_100_1_111011010100;
      patterns[60749] = 29'b1_110110101001_101_0_111101101010;
      patterns[60750] = 29'b1_110110101001_110_1_110110101001;
      patterns[60751] = 29'b1_110110101001_111_1_110110101001;
      patterns[60752] = 29'b1_110110101010_000_1_110110101010;
      patterns[60753] = 29'b1_110110101010_001_1_101010110110;
      patterns[60754] = 29'b1_110110101010_010_1_101101010101;
      patterns[60755] = 29'b1_110110101010_011_1_011010101011;
      patterns[60756] = 29'b1_110110101010_100_0_111011010101;
      patterns[60757] = 29'b1_110110101010_101_1_011101101010;
      patterns[60758] = 29'b1_110110101010_110_1_110110101010;
      patterns[60759] = 29'b1_110110101010_111_1_110110101010;
      patterns[60760] = 29'b1_110110101011_000_1_110110101011;
      patterns[60761] = 29'b1_110110101011_001_1_101011110110;
      patterns[60762] = 29'b1_110110101011_010_1_101101010111;
      patterns[60763] = 29'b1_110110101011_011_1_011010101111;
      patterns[60764] = 29'b1_110110101011_100_1_111011010101;
      patterns[60765] = 29'b1_110110101011_101_1_111101101010;
      patterns[60766] = 29'b1_110110101011_110_1_110110101011;
      patterns[60767] = 29'b1_110110101011_111_1_110110101011;
      patterns[60768] = 29'b1_110110101100_000_1_110110101100;
      patterns[60769] = 29'b1_110110101100_001_1_101100110110;
      patterns[60770] = 29'b1_110110101100_010_1_101101011001;
      patterns[60771] = 29'b1_110110101100_011_1_011010110011;
      patterns[60772] = 29'b1_110110101100_100_0_111011010110;
      patterns[60773] = 29'b1_110110101100_101_0_011101101011;
      patterns[60774] = 29'b1_110110101100_110_1_110110101100;
      patterns[60775] = 29'b1_110110101100_111_1_110110101100;
      patterns[60776] = 29'b1_110110101101_000_1_110110101101;
      patterns[60777] = 29'b1_110110101101_001_1_101101110110;
      patterns[60778] = 29'b1_110110101101_010_1_101101011011;
      patterns[60779] = 29'b1_110110101101_011_1_011010110111;
      patterns[60780] = 29'b1_110110101101_100_1_111011010110;
      patterns[60781] = 29'b1_110110101101_101_0_111101101011;
      patterns[60782] = 29'b1_110110101101_110_1_110110101101;
      patterns[60783] = 29'b1_110110101101_111_1_110110101101;
      patterns[60784] = 29'b1_110110101110_000_1_110110101110;
      patterns[60785] = 29'b1_110110101110_001_1_101110110110;
      patterns[60786] = 29'b1_110110101110_010_1_101101011101;
      patterns[60787] = 29'b1_110110101110_011_1_011010111011;
      patterns[60788] = 29'b1_110110101110_100_0_111011010111;
      patterns[60789] = 29'b1_110110101110_101_1_011101101011;
      patterns[60790] = 29'b1_110110101110_110_1_110110101110;
      patterns[60791] = 29'b1_110110101110_111_1_110110101110;
      patterns[60792] = 29'b1_110110101111_000_1_110110101111;
      patterns[60793] = 29'b1_110110101111_001_1_101111110110;
      patterns[60794] = 29'b1_110110101111_010_1_101101011111;
      patterns[60795] = 29'b1_110110101111_011_1_011010111111;
      patterns[60796] = 29'b1_110110101111_100_1_111011010111;
      patterns[60797] = 29'b1_110110101111_101_1_111101101011;
      patterns[60798] = 29'b1_110110101111_110_1_110110101111;
      patterns[60799] = 29'b1_110110101111_111_1_110110101111;
      patterns[60800] = 29'b1_110110110000_000_1_110110110000;
      patterns[60801] = 29'b1_110110110000_001_1_110000110110;
      patterns[60802] = 29'b1_110110110000_010_1_101101100001;
      patterns[60803] = 29'b1_110110110000_011_1_011011000011;
      patterns[60804] = 29'b1_110110110000_100_0_111011011000;
      patterns[60805] = 29'b1_110110110000_101_0_011101101100;
      patterns[60806] = 29'b1_110110110000_110_1_110110110000;
      patterns[60807] = 29'b1_110110110000_111_1_110110110000;
      patterns[60808] = 29'b1_110110110001_000_1_110110110001;
      patterns[60809] = 29'b1_110110110001_001_1_110001110110;
      patterns[60810] = 29'b1_110110110001_010_1_101101100011;
      patterns[60811] = 29'b1_110110110001_011_1_011011000111;
      patterns[60812] = 29'b1_110110110001_100_1_111011011000;
      patterns[60813] = 29'b1_110110110001_101_0_111101101100;
      patterns[60814] = 29'b1_110110110001_110_1_110110110001;
      patterns[60815] = 29'b1_110110110001_111_1_110110110001;
      patterns[60816] = 29'b1_110110110010_000_1_110110110010;
      patterns[60817] = 29'b1_110110110010_001_1_110010110110;
      patterns[60818] = 29'b1_110110110010_010_1_101101100101;
      patterns[60819] = 29'b1_110110110010_011_1_011011001011;
      patterns[60820] = 29'b1_110110110010_100_0_111011011001;
      patterns[60821] = 29'b1_110110110010_101_1_011101101100;
      patterns[60822] = 29'b1_110110110010_110_1_110110110010;
      patterns[60823] = 29'b1_110110110010_111_1_110110110010;
      patterns[60824] = 29'b1_110110110011_000_1_110110110011;
      patterns[60825] = 29'b1_110110110011_001_1_110011110110;
      patterns[60826] = 29'b1_110110110011_010_1_101101100111;
      patterns[60827] = 29'b1_110110110011_011_1_011011001111;
      patterns[60828] = 29'b1_110110110011_100_1_111011011001;
      patterns[60829] = 29'b1_110110110011_101_1_111101101100;
      patterns[60830] = 29'b1_110110110011_110_1_110110110011;
      patterns[60831] = 29'b1_110110110011_111_1_110110110011;
      patterns[60832] = 29'b1_110110110100_000_1_110110110100;
      patterns[60833] = 29'b1_110110110100_001_1_110100110110;
      patterns[60834] = 29'b1_110110110100_010_1_101101101001;
      patterns[60835] = 29'b1_110110110100_011_1_011011010011;
      patterns[60836] = 29'b1_110110110100_100_0_111011011010;
      patterns[60837] = 29'b1_110110110100_101_0_011101101101;
      patterns[60838] = 29'b1_110110110100_110_1_110110110100;
      patterns[60839] = 29'b1_110110110100_111_1_110110110100;
      patterns[60840] = 29'b1_110110110101_000_1_110110110101;
      patterns[60841] = 29'b1_110110110101_001_1_110101110110;
      patterns[60842] = 29'b1_110110110101_010_1_101101101011;
      patterns[60843] = 29'b1_110110110101_011_1_011011010111;
      patterns[60844] = 29'b1_110110110101_100_1_111011011010;
      patterns[60845] = 29'b1_110110110101_101_0_111101101101;
      patterns[60846] = 29'b1_110110110101_110_1_110110110101;
      patterns[60847] = 29'b1_110110110101_111_1_110110110101;
      patterns[60848] = 29'b1_110110110110_000_1_110110110110;
      patterns[60849] = 29'b1_110110110110_001_1_110110110110;
      patterns[60850] = 29'b1_110110110110_010_1_101101101101;
      patterns[60851] = 29'b1_110110110110_011_1_011011011011;
      patterns[60852] = 29'b1_110110110110_100_0_111011011011;
      patterns[60853] = 29'b1_110110110110_101_1_011101101101;
      patterns[60854] = 29'b1_110110110110_110_1_110110110110;
      patterns[60855] = 29'b1_110110110110_111_1_110110110110;
      patterns[60856] = 29'b1_110110110111_000_1_110110110111;
      patterns[60857] = 29'b1_110110110111_001_1_110111110110;
      patterns[60858] = 29'b1_110110110111_010_1_101101101111;
      patterns[60859] = 29'b1_110110110111_011_1_011011011111;
      patterns[60860] = 29'b1_110110110111_100_1_111011011011;
      patterns[60861] = 29'b1_110110110111_101_1_111101101101;
      patterns[60862] = 29'b1_110110110111_110_1_110110110111;
      patterns[60863] = 29'b1_110110110111_111_1_110110110111;
      patterns[60864] = 29'b1_110110111000_000_1_110110111000;
      patterns[60865] = 29'b1_110110111000_001_1_111000110110;
      patterns[60866] = 29'b1_110110111000_010_1_101101110001;
      patterns[60867] = 29'b1_110110111000_011_1_011011100011;
      patterns[60868] = 29'b1_110110111000_100_0_111011011100;
      patterns[60869] = 29'b1_110110111000_101_0_011101101110;
      patterns[60870] = 29'b1_110110111000_110_1_110110111000;
      patterns[60871] = 29'b1_110110111000_111_1_110110111000;
      patterns[60872] = 29'b1_110110111001_000_1_110110111001;
      patterns[60873] = 29'b1_110110111001_001_1_111001110110;
      patterns[60874] = 29'b1_110110111001_010_1_101101110011;
      patterns[60875] = 29'b1_110110111001_011_1_011011100111;
      patterns[60876] = 29'b1_110110111001_100_1_111011011100;
      patterns[60877] = 29'b1_110110111001_101_0_111101101110;
      patterns[60878] = 29'b1_110110111001_110_1_110110111001;
      patterns[60879] = 29'b1_110110111001_111_1_110110111001;
      patterns[60880] = 29'b1_110110111010_000_1_110110111010;
      patterns[60881] = 29'b1_110110111010_001_1_111010110110;
      patterns[60882] = 29'b1_110110111010_010_1_101101110101;
      patterns[60883] = 29'b1_110110111010_011_1_011011101011;
      patterns[60884] = 29'b1_110110111010_100_0_111011011101;
      patterns[60885] = 29'b1_110110111010_101_1_011101101110;
      patterns[60886] = 29'b1_110110111010_110_1_110110111010;
      patterns[60887] = 29'b1_110110111010_111_1_110110111010;
      patterns[60888] = 29'b1_110110111011_000_1_110110111011;
      patterns[60889] = 29'b1_110110111011_001_1_111011110110;
      patterns[60890] = 29'b1_110110111011_010_1_101101110111;
      patterns[60891] = 29'b1_110110111011_011_1_011011101111;
      patterns[60892] = 29'b1_110110111011_100_1_111011011101;
      patterns[60893] = 29'b1_110110111011_101_1_111101101110;
      patterns[60894] = 29'b1_110110111011_110_1_110110111011;
      patterns[60895] = 29'b1_110110111011_111_1_110110111011;
      patterns[60896] = 29'b1_110110111100_000_1_110110111100;
      patterns[60897] = 29'b1_110110111100_001_1_111100110110;
      patterns[60898] = 29'b1_110110111100_010_1_101101111001;
      patterns[60899] = 29'b1_110110111100_011_1_011011110011;
      patterns[60900] = 29'b1_110110111100_100_0_111011011110;
      patterns[60901] = 29'b1_110110111100_101_0_011101101111;
      patterns[60902] = 29'b1_110110111100_110_1_110110111100;
      patterns[60903] = 29'b1_110110111100_111_1_110110111100;
      patterns[60904] = 29'b1_110110111101_000_1_110110111101;
      patterns[60905] = 29'b1_110110111101_001_1_111101110110;
      patterns[60906] = 29'b1_110110111101_010_1_101101111011;
      patterns[60907] = 29'b1_110110111101_011_1_011011110111;
      patterns[60908] = 29'b1_110110111101_100_1_111011011110;
      patterns[60909] = 29'b1_110110111101_101_0_111101101111;
      patterns[60910] = 29'b1_110110111101_110_1_110110111101;
      patterns[60911] = 29'b1_110110111101_111_1_110110111101;
      patterns[60912] = 29'b1_110110111110_000_1_110110111110;
      patterns[60913] = 29'b1_110110111110_001_1_111110110110;
      patterns[60914] = 29'b1_110110111110_010_1_101101111101;
      patterns[60915] = 29'b1_110110111110_011_1_011011111011;
      patterns[60916] = 29'b1_110110111110_100_0_111011011111;
      patterns[60917] = 29'b1_110110111110_101_1_011101101111;
      patterns[60918] = 29'b1_110110111110_110_1_110110111110;
      patterns[60919] = 29'b1_110110111110_111_1_110110111110;
      patterns[60920] = 29'b1_110110111111_000_1_110110111111;
      patterns[60921] = 29'b1_110110111111_001_1_111111110110;
      patterns[60922] = 29'b1_110110111111_010_1_101101111111;
      patterns[60923] = 29'b1_110110111111_011_1_011011111111;
      patterns[60924] = 29'b1_110110111111_100_1_111011011111;
      patterns[60925] = 29'b1_110110111111_101_1_111101101111;
      patterns[60926] = 29'b1_110110111111_110_1_110110111111;
      patterns[60927] = 29'b1_110110111111_111_1_110110111111;
      patterns[60928] = 29'b1_110111000000_000_1_110111000000;
      patterns[60929] = 29'b1_110111000000_001_1_000000110111;
      patterns[60930] = 29'b1_110111000000_010_1_101110000001;
      patterns[60931] = 29'b1_110111000000_011_1_011100000011;
      patterns[60932] = 29'b1_110111000000_100_0_111011100000;
      patterns[60933] = 29'b1_110111000000_101_0_011101110000;
      patterns[60934] = 29'b1_110111000000_110_1_110111000000;
      patterns[60935] = 29'b1_110111000000_111_1_110111000000;
      patterns[60936] = 29'b1_110111000001_000_1_110111000001;
      patterns[60937] = 29'b1_110111000001_001_1_000001110111;
      patterns[60938] = 29'b1_110111000001_010_1_101110000011;
      patterns[60939] = 29'b1_110111000001_011_1_011100000111;
      patterns[60940] = 29'b1_110111000001_100_1_111011100000;
      patterns[60941] = 29'b1_110111000001_101_0_111101110000;
      patterns[60942] = 29'b1_110111000001_110_1_110111000001;
      patterns[60943] = 29'b1_110111000001_111_1_110111000001;
      patterns[60944] = 29'b1_110111000010_000_1_110111000010;
      patterns[60945] = 29'b1_110111000010_001_1_000010110111;
      patterns[60946] = 29'b1_110111000010_010_1_101110000101;
      patterns[60947] = 29'b1_110111000010_011_1_011100001011;
      patterns[60948] = 29'b1_110111000010_100_0_111011100001;
      patterns[60949] = 29'b1_110111000010_101_1_011101110000;
      patterns[60950] = 29'b1_110111000010_110_1_110111000010;
      patterns[60951] = 29'b1_110111000010_111_1_110111000010;
      patterns[60952] = 29'b1_110111000011_000_1_110111000011;
      patterns[60953] = 29'b1_110111000011_001_1_000011110111;
      patterns[60954] = 29'b1_110111000011_010_1_101110000111;
      patterns[60955] = 29'b1_110111000011_011_1_011100001111;
      patterns[60956] = 29'b1_110111000011_100_1_111011100001;
      patterns[60957] = 29'b1_110111000011_101_1_111101110000;
      patterns[60958] = 29'b1_110111000011_110_1_110111000011;
      patterns[60959] = 29'b1_110111000011_111_1_110111000011;
      patterns[60960] = 29'b1_110111000100_000_1_110111000100;
      patterns[60961] = 29'b1_110111000100_001_1_000100110111;
      patterns[60962] = 29'b1_110111000100_010_1_101110001001;
      patterns[60963] = 29'b1_110111000100_011_1_011100010011;
      patterns[60964] = 29'b1_110111000100_100_0_111011100010;
      patterns[60965] = 29'b1_110111000100_101_0_011101110001;
      patterns[60966] = 29'b1_110111000100_110_1_110111000100;
      patterns[60967] = 29'b1_110111000100_111_1_110111000100;
      patterns[60968] = 29'b1_110111000101_000_1_110111000101;
      patterns[60969] = 29'b1_110111000101_001_1_000101110111;
      patterns[60970] = 29'b1_110111000101_010_1_101110001011;
      patterns[60971] = 29'b1_110111000101_011_1_011100010111;
      patterns[60972] = 29'b1_110111000101_100_1_111011100010;
      patterns[60973] = 29'b1_110111000101_101_0_111101110001;
      patterns[60974] = 29'b1_110111000101_110_1_110111000101;
      patterns[60975] = 29'b1_110111000101_111_1_110111000101;
      patterns[60976] = 29'b1_110111000110_000_1_110111000110;
      patterns[60977] = 29'b1_110111000110_001_1_000110110111;
      patterns[60978] = 29'b1_110111000110_010_1_101110001101;
      patterns[60979] = 29'b1_110111000110_011_1_011100011011;
      patterns[60980] = 29'b1_110111000110_100_0_111011100011;
      patterns[60981] = 29'b1_110111000110_101_1_011101110001;
      patterns[60982] = 29'b1_110111000110_110_1_110111000110;
      patterns[60983] = 29'b1_110111000110_111_1_110111000110;
      patterns[60984] = 29'b1_110111000111_000_1_110111000111;
      patterns[60985] = 29'b1_110111000111_001_1_000111110111;
      patterns[60986] = 29'b1_110111000111_010_1_101110001111;
      patterns[60987] = 29'b1_110111000111_011_1_011100011111;
      patterns[60988] = 29'b1_110111000111_100_1_111011100011;
      patterns[60989] = 29'b1_110111000111_101_1_111101110001;
      patterns[60990] = 29'b1_110111000111_110_1_110111000111;
      patterns[60991] = 29'b1_110111000111_111_1_110111000111;
      patterns[60992] = 29'b1_110111001000_000_1_110111001000;
      patterns[60993] = 29'b1_110111001000_001_1_001000110111;
      patterns[60994] = 29'b1_110111001000_010_1_101110010001;
      patterns[60995] = 29'b1_110111001000_011_1_011100100011;
      patterns[60996] = 29'b1_110111001000_100_0_111011100100;
      patterns[60997] = 29'b1_110111001000_101_0_011101110010;
      patterns[60998] = 29'b1_110111001000_110_1_110111001000;
      patterns[60999] = 29'b1_110111001000_111_1_110111001000;
      patterns[61000] = 29'b1_110111001001_000_1_110111001001;
      patterns[61001] = 29'b1_110111001001_001_1_001001110111;
      patterns[61002] = 29'b1_110111001001_010_1_101110010011;
      patterns[61003] = 29'b1_110111001001_011_1_011100100111;
      patterns[61004] = 29'b1_110111001001_100_1_111011100100;
      patterns[61005] = 29'b1_110111001001_101_0_111101110010;
      patterns[61006] = 29'b1_110111001001_110_1_110111001001;
      patterns[61007] = 29'b1_110111001001_111_1_110111001001;
      patterns[61008] = 29'b1_110111001010_000_1_110111001010;
      patterns[61009] = 29'b1_110111001010_001_1_001010110111;
      patterns[61010] = 29'b1_110111001010_010_1_101110010101;
      patterns[61011] = 29'b1_110111001010_011_1_011100101011;
      patterns[61012] = 29'b1_110111001010_100_0_111011100101;
      patterns[61013] = 29'b1_110111001010_101_1_011101110010;
      patterns[61014] = 29'b1_110111001010_110_1_110111001010;
      patterns[61015] = 29'b1_110111001010_111_1_110111001010;
      patterns[61016] = 29'b1_110111001011_000_1_110111001011;
      patterns[61017] = 29'b1_110111001011_001_1_001011110111;
      patterns[61018] = 29'b1_110111001011_010_1_101110010111;
      patterns[61019] = 29'b1_110111001011_011_1_011100101111;
      patterns[61020] = 29'b1_110111001011_100_1_111011100101;
      patterns[61021] = 29'b1_110111001011_101_1_111101110010;
      patterns[61022] = 29'b1_110111001011_110_1_110111001011;
      patterns[61023] = 29'b1_110111001011_111_1_110111001011;
      patterns[61024] = 29'b1_110111001100_000_1_110111001100;
      patterns[61025] = 29'b1_110111001100_001_1_001100110111;
      patterns[61026] = 29'b1_110111001100_010_1_101110011001;
      patterns[61027] = 29'b1_110111001100_011_1_011100110011;
      patterns[61028] = 29'b1_110111001100_100_0_111011100110;
      patterns[61029] = 29'b1_110111001100_101_0_011101110011;
      patterns[61030] = 29'b1_110111001100_110_1_110111001100;
      patterns[61031] = 29'b1_110111001100_111_1_110111001100;
      patterns[61032] = 29'b1_110111001101_000_1_110111001101;
      patterns[61033] = 29'b1_110111001101_001_1_001101110111;
      patterns[61034] = 29'b1_110111001101_010_1_101110011011;
      patterns[61035] = 29'b1_110111001101_011_1_011100110111;
      patterns[61036] = 29'b1_110111001101_100_1_111011100110;
      patterns[61037] = 29'b1_110111001101_101_0_111101110011;
      patterns[61038] = 29'b1_110111001101_110_1_110111001101;
      patterns[61039] = 29'b1_110111001101_111_1_110111001101;
      patterns[61040] = 29'b1_110111001110_000_1_110111001110;
      patterns[61041] = 29'b1_110111001110_001_1_001110110111;
      patterns[61042] = 29'b1_110111001110_010_1_101110011101;
      patterns[61043] = 29'b1_110111001110_011_1_011100111011;
      patterns[61044] = 29'b1_110111001110_100_0_111011100111;
      patterns[61045] = 29'b1_110111001110_101_1_011101110011;
      patterns[61046] = 29'b1_110111001110_110_1_110111001110;
      patterns[61047] = 29'b1_110111001110_111_1_110111001110;
      patterns[61048] = 29'b1_110111001111_000_1_110111001111;
      patterns[61049] = 29'b1_110111001111_001_1_001111110111;
      patterns[61050] = 29'b1_110111001111_010_1_101110011111;
      patterns[61051] = 29'b1_110111001111_011_1_011100111111;
      patterns[61052] = 29'b1_110111001111_100_1_111011100111;
      patterns[61053] = 29'b1_110111001111_101_1_111101110011;
      patterns[61054] = 29'b1_110111001111_110_1_110111001111;
      patterns[61055] = 29'b1_110111001111_111_1_110111001111;
      patterns[61056] = 29'b1_110111010000_000_1_110111010000;
      patterns[61057] = 29'b1_110111010000_001_1_010000110111;
      patterns[61058] = 29'b1_110111010000_010_1_101110100001;
      patterns[61059] = 29'b1_110111010000_011_1_011101000011;
      patterns[61060] = 29'b1_110111010000_100_0_111011101000;
      patterns[61061] = 29'b1_110111010000_101_0_011101110100;
      patterns[61062] = 29'b1_110111010000_110_1_110111010000;
      patterns[61063] = 29'b1_110111010000_111_1_110111010000;
      patterns[61064] = 29'b1_110111010001_000_1_110111010001;
      patterns[61065] = 29'b1_110111010001_001_1_010001110111;
      patterns[61066] = 29'b1_110111010001_010_1_101110100011;
      patterns[61067] = 29'b1_110111010001_011_1_011101000111;
      patterns[61068] = 29'b1_110111010001_100_1_111011101000;
      patterns[61069] = 29'b1_110111010001_101_0_111101110100;
      patterns[61070] = 29'b1_110111010001_110_1_110111010001;
      patterns[61071] = 29'b1_110111010001_111_1_110111010001;
      patterns[61072] = 29'b1_110111010010_000_1_110111010010;
      patterns[61073] = 29'b1_110111010010_001_1_010010110111;
      patterns[61074] = 29'b1_110111010010_010_1_101110100101;
      patterns[61075] = 29'b1_110111010010_011_1_011101001011;
      patterns[61076] = 29'b1_110111010010_100_0_111011101001;
      patterns[61077] = 29'b1_110111010010_101_1_011101110100;
      patterns[61078] = 29'b1_110111010010_110_1_110111010010;
      patterns[61079] = 29'b1_110111010010_111_1_110111010010;
      patterns[61080] = 29'b1_110111010011_000_1_110111010011;
      patterns[61081] = 29'b1_110111010011_001_1_010011110111;
      patterns[61082] = 29'b1_110111010011_010_1_101110100111;
      patterns[61083] = 29'b1_110111010011_011_1_011101001111;
      patterns[61084] = 29'b1_110111010011_100_1_111011101001;
      patterns[61085] = 29'b1_110111010011_101_1_111101110100;
      patterns[61086] = 29'b1_110111010011_110_1_110111010011;
      patterns[61087] = 29'b1_110111010011_111_1_110111010011;
      patterns[61088] = 29'b1_110111010100_000_1_110111010100;
      patterns[61089] = 29'b1_110111010100_001_1_010100110111;
      patterns[61090] = 29'b1_110111010100_010_1_101110101001;
      patterns[61091] = 29'b1_110111010100_011_1_011101010011;
      patterns[61092] = 29'b1_110111010100_100_0_111011101010;
      patterns[61093] = 29'b1_110111010100_101_0_011101110101;
      patterns[61094] = 29'b1_110111010100_110_1_110111010100;
      patterns[61095] = 29'b1_110111010100_111_1_110111010100;
      patterns[61096] = 29'b1_110111010101_000_1_110111010101;
      patterns[61097] = 29'b1_110111010101_001_1_010101110111;
      patterns[61098] = 29'b1_110111010101_010_1_101110101011;
      patterns[61099] = 29'b1_110111010101_011_1_011101010111;
      patterns[61100] = 29'b1_110111010101_100_1_111011101010;
      patterns[61101] = 29'b1_110111010101_101_0_111101110101;
      patterns[61102] = 29'b1_110111010101_110_1_110111010101;
      patterns[61103] = 29'b1_110111010101_111_1_110111010101;
      patterns[61104] = 29'b1_110111010110_000_1_110111010110;
      patterns[61105] = 29'b1_110111010110_001_1_010110110111;
      patterns[61106] = 29'b1_110111010110_010_1_101110101101;
      patterns[61107] = 29'b1_110111010110_011_1_011101011011;
      patterns[61108] = 29'b1_110111010110_100_0_111011101011;
      patterns[61109] = 29'b1_110111010110_101_1_011101110101;
      patterns[61110] = 29'b1_110111010110_110_1_110111010110;
      patterns[61111] = 29'b1_110111010110_111_1_110111010110;
      patterns[61112] = 29'b1_110111010111_000_1_110111010111;
      patterns[61113] = 29'b1_110111010111_001_1_010111110111;
      patterns[61114] = 29'b1_110111010111_010_1_101110101111;
      patterns[61115] = 29'b1_110111010111_011_1_011101011111;
      patterns[61116] = 29'b1_110111010111_100_1_111011101011;
      patterns[61117] = 29'b1_110111010111_101_1_111101110101;
      patterns[61118] = 29'b1_110111010111_110_1_110111010111;
      patterns[61119] = 29'b1_110111010111_111_1_110111010111;
      patterns[61120] = 29'b1_110111011000_000_1_110111011000;
      patterns[61121] = 29'b1_110111011000_001_1_011000110111;
      patterns[61122] = 29'b1_110111011000_010_1_101110110001;
      patterns[61123] = 29'b1_110111011000_011_1_011101100011;
      patterns[61124] = 29'b1_110111011000_100_0_111011101100;
      patterns[61125] = 29'b1_110111011000_101_0_011101110110;
      patterns[61126] = 29'b1_110111011000_110_1_110111011000;
      patterns[61127] = 29'b1_110111011000_111_1_110111011000;
      patterns[61128] = 29'b1_110111011001_000_1_110111011001;
      patterns[61129] = 29'b1_110111011001_001_1_011001110111;
      patterns[61130] = 29'b1_110111011001_010_1_101110110011;
      patterns[61131] = 29'b1_110111011001_011_1_011101100111;
      patterns[61132] = 29'b1_110111011001_100_1_111011101100;
      patterns[61133] = 29'b1_110111011001_101_0_111101110110;
      patterns[61134] = 29'b1_110111011001_110_1_110111011001;
      patterns[61135] = 29'b1_110111011001_111_1_110111011001;
      patterns[61136] = 29'b1_110111011010_000_1_110111011010;
      patterns[61137] = 29'b1_110111011010_001_1_011010110111;
      patterns[61138] = 29'b1_110111011010_010_1_101110110101;
      patterns[61139] = 29'b1_110111011010_011_1_011101101011;
      patterns[61140] = 29'b1_110111011010_100_0_111011101101;
      patterns[61141] = 29'b1_110111011010_101_1_011101110110;
      patterns[61142] = 29'b1_110111011010_110_1_110111011010;
      patterns[61143] = 29'b1_110111011010_111_1_110111011010;
      patterns[61144] = 29'b1_110111011011_000_1_110111011011;
      patterns[61145] = 29'b1_110111011011_001_1_011011110111;
      patterns[61146] = 29'b1_110111011011_010_1_101110110111;
      patterns[61147] = 29'b1_110111011011_011_1_011101101111;
      patterns[61148] = 29'b1_110111011011_100_1_111011101101;
      patterns[61149] = 29'b1_110111011011_101_1_111101110110;
      patterns[61150] = 29'b1_110111011011_110_1_110111011011;
      patterns[61151] = 29'b1_110111011011_111_1_110111011011;
      patterns[61152] = 29'b1_110111011100_000_1_110111011100;
      patterns[61153] = 29'b1_110111011100_001_1_011100110111;
      patterns[61154] = 29'b1_110111011100_010_1_101110111001;
      patterns[61155] = 29'b1_110111011100_011_1_011101110011;
      patterns[61156] = 29'b1_110111011100_100_0_111011101110;
      patterns[61157] = 29'b1_110111011100_101_0_011101110111;
      patterns[61158] = 29'b1_110111011100_110_1_110111011100;
      patterns[61159] = 29'b1_110111011100_111_1_110111011100;
      patterns[61160] = 29'b1_110111011101_000_1_110111011101;
      patterns[61161] = 29'b1_110111011101_001_1_011101110111;
      patterns[61162] = 29'b1_110111011101_010_1_101110111011;
      patterns[61163] = 29'b1_110111011101_011_1_011101110111;
      patterns[61164] = 29'b1_110111011101_100_1_111011101110;
      patterns[61165] = 29'b1_110111011101_101_0_111101110111;
      patterns[61166] = 29'b1_110111011101_110_1_110111011101;
      patterns[61167] = 29'b1_110111011101_111_1_110111011101;
      patterns[61168] = 29'b1_110111011110_000_1_110111011110;
      patterns[61169] = 29'b1_110111011110_001_1_011110110111;
      patterns[61170] = 29'b1_110111011110_010_1_101110111101;
      patterns[61171] = 29'b1_110111011110_011_1_011101111011;
      patterns[61172] = 29'b1_110111011110_100_0_111011101111;
      patterns[61173] = 29'b1_110111011110_101_1_011101110111;
      patterns[61174] = 29'b1_110111011110_110_1_110111011110;
      patterns[61175] = 29'b1_110111011110_111_1_110111011110;
      patterns[61176] = 29'b1_110111011111_000_1_110111011111;
      patterns[61177] = 29'b1_110111011111_001_1_011111110111;
      patterns[61178] = 29'b1_110111011111_010_1_101110111111;
      patterns[61179] = 29'b1_110111011111_011_1_011101111111;
      patterns[61180] = 29'b1_110111011111_100_1_111011101111;
      patterns[61181] = 29'b1_110111011111_101_1_111101110111;
      patterns[61182] = 29'b1_110111011111_110_1_110111011111;
      patterns[61183] = 29'b1_110111011111_111_1_110111011111;
      patterns[61184] = 29'b1_110111100000_000_1_110111100000;
      patterns[61185] = 29'b1_110111100000_001_1_100000110111;
      patterns[61186] = 29'b1_110111100000_010_1_101111000001;
      patterns[61187] = 29'b1_110111100000_011_1_011110000011;
      patterns[61188] = 29'b1_110111100000_100_0_111011110000;
      patterns[61189] = 29'b1_110111100000_101_0_011101111000;
      patterns[61190] = 29'b1_110111100000_110_1_110111100000;
      patterns[61191] = 29'b1_110111100000_111_1_110111100000;
      patterns[61192] = 29'b1_110111100001_000_1_110111100001;
      patterns[61193] = 29'b1_110111100001_001_1_100001110111;
      patterns[61194] = 29'b1_110111100001_010_1_101111000011;
      patterns[61195] = 29'b1_110111100001_011_1_011110000111;
      patterns[61196] = 29'b1_110111100001_100_1_111011110000;
      patterns[61197] = 29'b1_110111100001_101_0_111101111000;
      patterns[61198] = 29'b1_110111100001_110_1_110111100001;
      patterns[61199] = 29'b1_110111100001_111_1_110111100001;
      patterns[61200] = 29'b1_110111100010_000_1_110111100010;
      patterns[61201] = 29'b1_110111100010_001_1_100010110111;
      patterns[61202] = 29'b1_110111100010_010_1_101111000101;
      patterns[61203] = 29'b1_110111100010_011_1_011110001011;
      patterns[61204] = 29'b1_110111100010_100_0_111011110001;
      patterns[61205] = 29'b1_110111100010_101_1_011101111000;
      patterns[61206] = 29'b1_110111100010_110_1_110111100010;
      patterns[61207] = 29'b1_110111100010_111_1_110111100010;
      patterns[61208] = 29'b1_110111100011_000_1_110111100011;
      patterns[61209] = 29'b1_110111100011_001_1_100011110111;
      patterns[61210] = 29'b1_110111100011_010_1_101111000111;
      patterns[61211] = 29'b1_110111100011_011_1_011110001111;
      patterns[61212] = 29'b1_110111100011_100_1_111011110001;
      patterns[61213] = 29'b1_110111100011_101_1_111101111000;
      patterns[61214] = 29'b1_110111100011_110_1_110111100011;
      patterns[61215] = 29'b1_110111100011_111_1_110111100011;
      patterns[61216] = 29'b1_110111100100_000_1_110111100100;
      patterns[61217] = 29'b1_110111100100_001_1_100100110111;
      patterns[61218] = 29'b1_110111100100_010_1_101111001001;
      patterns[61219] = 29'b1_110111100100_011_1_011110010011;
      patterns[61220] = 29'b1_110111100100_100_0_111011110010;
      patterns[61221] = 29'b1_110111100100_101_0_011101111001;
      patterns[61222] = 29'b1_110111100100_110_1_110111100100;
      patterns[61223] = 29'b1_110111100100_111_1_110111100100;
      patterns[61224] = 29'b1_110111100101_000_1_110111100101;
      patterns[61225] = 29'b1_110111100101_001_1_100101110111;
      patterns[61226] = 29'b1_110111100101_010_1_101111001011;
      patterns[61227] = 29'b1_110111100101_011_1_011110010111;
      patterns[61228] = 29'b1_110111100101_100_1_111011110010;
      patterns[61229] = 29'b1_110111100101_101_0_111101111001;
      patterns[61230] = 29'b1_110111100101_110_1_110111100101;
      patterns[61231] = 29'b1_110111100101_111_1_110111100101;
      patterns[61232] = 29'b1_110111100110_000_1_110111100110;
      patterns[61233] = 29'b1_110111100110_001_1_100110110111;
      patterns[61234] = 29'b1_110111100110_010_1_101111001101;
      patterns[61235] = 29'b1_110111100110_011_1_011110011011;
      patterns[61236] = 29'b1_110111100110_100_0_111011110011;
      patterns[61237] = 29'b1_110111100110_101_1_011101111001;
      patterns[61238] = 29'b1_110111100110_110_1_110111100110;
      patterns[61239] = 29'b1_110111100110_111_1_110111100110;
      patterns[61240] = 29'b1_110111100111_000_1_110111100111;
      patterns[61241] = 29'b1_110111100111_001_1_100111110111;
      patterns[61242] = 29'b1_110111100111_010_1_101111001111;
      patterns[61243] = 29'b1_110111100111_011_1_011110011111;
      patterns[61244] = 29'b1_110111100111_100_1_111011110011;
      patterns[61245] = 29'b1_110111100111_101_1_111101111001;
      patterns[61246] = 29'b1_110111100111_110_1_110111100111;
      patterns[61247] = 29'b1_110111100111_111_1_110111100111;
      patterns[61248] = 29'b1_110111101000_000_1_110111101000;
      patterns[61249] = 29'b1_110111101000_001_1_101000110111;
      patterns[61250] = 29'b1_110111101000_010_1_101111010001;
      patterns[61251] = 29'b1_110111101000_011_1_011110100011;
      patterns[61252] = 29'b1_110111101000_100_0_111011110100;
      patterns[61253] = 29'b1_110111101000_101_0_011101111010;
      patterns[61254] = 29'b1_110111101000_110_1_110111101000;
      patterns[61255] = 29'b1_110111101000_111_1_110111101000;
      patterns[61256] = 29'b1_110111101001_000_1_110111101001;
      patterns[61257] = 29'b1_110111101001_001_1_101001110111;
      patterns[61258] = 29'b1_110111101001_010_1_101111010011;
      patterns[61259] = 29'b1_110111101001_011_1_011110100111;
      patterns[61260] = 29'b1_110111101001_100_1_111011110100;
      patterns[61261] = 29'b1_110111101001_101_0_111101111010;
      patterns[61262] = 29'b1_110111101001_110_1_110111101001;
      patterns[61263] = 29'b1_110111101001_111_1_110111101001;
      patterns[61264] = 29'b1_110111101010_000_1_110111101010;
      patterns[61265] = 29'b1_110111101010_001_1_101010110111;
      patterns[61266] = 29'b1_110111101010_010_1_101111010101;
      patterns[61267] = 29'b1_110111101010_011_1_011110101011;
      patterns[61268] = 29'b1_110111101010_100_0_111011110101;
      patterns[61269] = 29'b1_110111101010_101_1_011101111010;
      patterns[61270] = 29'b1_110111101010_110_1_110111101010;
      patterns[61271] = 29'b1_110111101010_111_1_110111101010;
      patterns[61272] = 29'b1_110111101011_000_1_110111101011;
      patterns[61273] = 29'b1_110111101011_001_1_101011110111;
      patterns[61274] = 29'b1_110111101011_010_1_101111010111;
      patterns[61275] = 29'b1_110111101011_011_1_011110101111;
      patterns[61276] = 29'b1_110111101011_100_1_111011110101;
      patterns[61277] = 29'b1_110111101011_101_1_111101111010;
      patterns[61278] = 29'b1_110111101011_110_1_110111101011;
      patterns[61279] = 29'b1_110111101011_111_1_110111101011;
      patterns[61280] = 29'b1_110111101100_000_1_110111101100;
      patterns[61281] = 29'b1_110111101100_001_1_101100110111;
      patterns[61282] = 29'b1_110111101100_010_1_101111011001;
      patterns[61283] = 29'b1_110111101100_011_1_011110110011;
      patterns[61284] = 29'b1_110111101100_100_0_111011110110;
      patterns[61285] = 29'b1_110111101100_101_0_011101111011;
      patterns[61286] = 29'b1_110111101100_110_1_110111101100;
      patterns[61287] = 29'b1_110111101100_111_1_110111101100;
      patterns[61288] = 29'b1_110111101101_000_1_110111101101;
      patterns[61289] = 29'b1_110111101101_001_1_101101110111;
      patterns[61290] = 29'b1_110111101101_010_1_101111011011;
      patterns[61291] = 29'b1_110111101101_011_1_011110110111;
      patterns[61292] = 29'b1_110111101101_100_1_111011110110;
      patterns[61293] = 29'b1_110111101101_101_0_111101111011;
      patterns[61294] = 29'b1_110111101101_110_1_110111101101;
      patterns[61295] = 29'b1_110111101101_111_1_110111101101;
      patterns[61296] = 29'b1_110111101110_000_1_110111101110;
      patterns[61297] = 29'b1_110111101110_001_1_101110110111;
      patterns[61298] = 29'b1_110111101110_010_1_101111011101;
      patterns[61299] = 29'b1_110111101110_011_1_011110111011;
      patterns[61300] = 29'b1_110111101110_100_0_111011110111;
      patterns[61301] = 29'b1_110111101110_101_1_011101111011;
      patterns[61302] = 29'b1_110111101110_110_1_110111101110;
      patterns[61303] = 29'b1_110111101110_111_1_110111101110;
      patterns[61304] = 29'b1_110111101111_000_1_110111101111;
      patterns[61305] = 29'b1_110111101111_001_1_101111110111;
      patterns[61306] = 29'b1_110111101111_010_1_101111011111;
      patterns[61307] = 29'b1_110111101111_011_1_011110111111;
      patterns[61308] = 29'b1_110111101111_100_1_111011110111;
      patterns[61309] = 29'b1_110111101111_101_1_111101111011;
      patterns[61310] = 29'b1_110111101111_110_1_110111101111;
      patterns[61311] = 29'b1_110111101111_111_1_110111101111;
      patterns[61312] = 29'b1_110111110000_000_1_110111110000;
      patterns[61313] = 29'b1_110111110000_001_1_110000110111;
      patterns[61314] = 29'b1_110111110000_010_1_101111100001;
      patterns[61315] = 29'b1_110111110000_011_1_011111000011;
      patterns[61316] = 29'b1_110111110000_100_0_111011111000;
      patterns[61317] = 29'b1_110111110000_101_0_011101111100;
      patterns[61318] = 29'b1_110111110000_110_1_110111110000;
      patterns[61319] = 29'b1_110111110000_111_1_110111110000;
      patterns[61320] = 29'b1_110111110001_000_1_110111110001;
      patterns[61321] = 29'b1_110111110001_001_1_110001110111;
      patterns[61322] = 29'b1_110111110001_010_1_101111100011;
      patterns[61323] = 29'b1_110111110001_011_1_011111000111;
      patterns[61324] = 29'b1_110111110001_100_1_111011111000;
      patterns[61325] = 29'b1_110111110001_101_0_111101111100;
      patterns[61326] = 29'b1_110111110001_110_1_110111110001;
      patterns[61327] = 29'b1_110111110001_111_1_110111110001;
      patterns[61328] = 29'b1_110111110010_000_1_110111110010;
      patterns[61329] = 29'b1_110111110010_001_1_110010110111;
      patterns[61330] = 29'b1_110111110010_010_1_101111100101;
      patterns[61331] = 29'b1_110111110010_011_1_011111001011;
      patterns[61332] = 29'b1_110111110010_100_0_111011111001;
      patterns[61333] = 29'b1_110111110010_101_1_011101111100;
      patterns[61334] = 29'b1_110111110010_110_1_110111110010;
      patterns[61335] = 29'b1_110111110010_111_1_110111110010;
      patterns[61336] = 29'b1_110111110011_000_1_110111110011;
      patterns[61337] = 29'b1_110111110011_001_1_110011110111;
      patterns[61338] = 29'b1_110111110011_010_1_101111100111;
      patterns[61339] = 29'b1_110111110011_011_1_011111001111;
      patterns[61340] = 29'b1_110111110011_100_1_111011111001;
      patterns[61341] = 29'b1_110111110011_101_1_111101111100;
      patterns[61342] = 29'b1_110111110011_110_1_110111110011;
      patterns[61343] = 29'b1_110111110011_111_1_110111110011;
      patterns[61344] = 29'b1_110111110100_000_1_110111110100;
      patterns[61345] = 29'b1_110111110100_001_1_110100110111;
      patterns[61346] = 29'b1_110111110100_010_1_101111101001;
      patterns[61347] = 29'b1_110111110100_011_1_011111010011;
      patterns[61348] = 29'b1_110111110100_100_0_111011111010;
      patterns[61349] = 29'b1_110111110100_101_0_011101111101;
      patterns[61350] = 29'b1_110111110100_110_1_110111110100;
      patterns[61351] = 29'b1_110111110100_111_1_110111110100;
      patterns[61352] = 29'b1_110111110101_000_1_110111110101;
      patterns[61353] = 29'b1_110111110101_001_1_110101110111;
      patterns[61354] = 29'b1_110111110101_010_1_101111101011;
      patterns[61355] = 29'b1_110111110101_011_1_011111010111;
      patterns[61356] = 29'b1_110111110101_100_1_111011111010;
      patterns[61357] = 29'b1_110111110101_101_0_111101111101;
      patterns[61358] = 29'b1_110111110101_110_1_110111110101;
      patterns[61359] = 29'b1_110111110101_111_1_110111110101;
      patterns[61360] = 29'b1_110111110110_000_1_110111110110;
      patterns[61361] = 29'b1_110111110110_001_1_110110110111;
      patterns[61362] = 29'b1_110111110110_010_1_101111101101;
      patterns[61363] = 29'b1_110111110110_011_1_011111011011;
      patterns[61364] = 29'b1_110111110110_100_0_111011111011;
      patterns[61365] = 29'b1_110111110110_101_1_011101111101;
      patterns[61366] = 29'b1_110111110110_110_1_110111110110;
      patterns[61367] = 29'b1_110111110110_111_1_110111110110;
      patterns[61368] = 29'b1_110111110111_000_1_110111110111;
      patterns[61369] = 29'b1_110111110111_001_1_110111110111;
      patterns[61370] = 29'b1_110111110111_010_1_101111101111;
      patterns[61371] = 29'b1_110111110111_011_1_011111011111;
      patterns[61372] = 29'b1_110111110111_100_1_111011111011;
      patterns[61373] = 29'b1_110111110111_101_1_111101111101;
      patterns[61374] = 29'b1_110111110111_110_1_110111110111;
      patterns[61375] = 29'b1_110111110111_111_1_110111110111;
      patterns[61376] = 29'b1_110111111000_000_1_110111111000;
      patterns[61377] = 29'b1_110111111000_001_1_111000110111;
      patterns[61378] = 29'b1_110111111000_010_1_101111110001;
      patterns[61379] = 29'b1_110111111000_011_1_011111100011;
      patterns[61380] = 29'b1_110111111000_100_0_111011111100;
      patterns[61381] = 29'b1_110111111000_101_0_011101111110;
      patterns[61382] = 29'b1_110111111000_110_1_110111111000;
      patterns[61383] = 29'b1_110111111000_111_1_110111111000;
      patterns[61384] = 29'b1_110111111001_000_1_110111111001;
      patterns[61385] = 29'b1_110111111001_001_1_111001110111;
      patterns[61386] = 29'b1_110111111001_010_1_101111110011;
      patterns[61387] = 29'b1_110111111001_011_1_011111100111;
      patterns[61388] = 29'b1_110111111001_100_1_111011111100;
      patterns[61389] = 29'b1_110111111001_101_0_111101111110;
      patterns[61390] = 29'b1_110111111001_110_1_110111111001;
      patterns[61391] = 29'b1_110111111001_111_1_110111111001;
      patterns[61392] = 29'b1_110111111010_000_1_110111111010;
      patterns[61393] = 29'b1_110111111010_001_1_111010110111;
      patterns[61394] = 29'b1_110111111010_010_1_101111110101;
      patterns[61395] = 29'b1_110111111010_011_1_011111101011;
      patterns[61396] = 29'b1_110111111010_100_0_111011111101;
      patterns[61397] = 29'b1_110111111010_101_1_011101111110;
      patterns[61398] = 29'b1_110111111010_110_1_110111111010;
      patterns[61399] = 29'b1_110111111010_111_1_110111111010;
      patterns[61400] = 29'b1_110111111011_000_1_110111111011;
      patterns[61401] = 29'b1_110111111011_001_1_111011110111;
      patterns[61402] = 29'b1_110111111011_010_1_101111110111;
      patterns[61403] = 29'b1_110111111011_011_1_011111101111;
      patterns[61404] = 29'b1_110111111011_100_1_111011111101;
      patterns[61405] = 29'b1_110111111011_101_1_111101111110;
      patterns[61406] = 29'b1_110111111011_110_1_110111111011;
      patterns[61407] = 29'b1_110111111011_111_1_110111111011;
      patterns[61408] = 29'b1_110111111100_000_1_110111111100;
      patterns[61409] = 29'b1_110111111100_001_1_111100110111;
      patterns[61410] = 29'b1_110111111100_010_1_101111111001;
      patterns[61411] = 29'b1_110111111100_011_1_011111110011;
      patterns[61412] = 29'b1_110111111100_100_0_111011111110;
      patterns[61413] = 29'b1_110111111100_101_0_011101111111;
      patterns[61414] = 29'b1_110111111100_110_1_110111111100;
      patterns[61415] = 29'b1_110111111100_111_1_110111111100;
      patterns[61416] = 29'b1_110111111101_000_1_110111111101;
      patterns[61417] = 29'b1_110111111101_001_1_111101110111;
      patterns[61418] = 29'b1_110111111101_010_1_101111111011;
      patterns[61419] = 29'b1_110111111101_011_1_011111110111;
      patterns[61420] = 29'b1_110111111101_100_1_111011111110;
      patterns[61421] = 29'b1_110111111101_101_0_111101111111;
      patterns[61422] = 29'b1_110111111101_110_1_110111111101;
      patterns[61423] = 29'b1_110111111101_111_1_110111111101;
      patterns[61424] = 29'b1_110111111110_000_1_110111111110;
      patterns[61425] = 29'b1_110111111110_001_1_111110110111;
      patterns[61426] = 29'b1_110111111110_010_1_101111111101;
      patterns[61427] = 29'b1_110111111110_011_1_011111111011;
      patterns[61428] = 29'b1_110111111110_100_0_111011111111;
      patterns[61429] = 29'b1_110111111110_101_1_011101111111;
      patterns[61430] = 29'b1_110111111110_110_1_110111111110;
      patterns[61431] = 29'b1_110111111110_111_1_110111111110;
      patterns[61432] = 29'b1_110111111111_000_1_110111111111;
      patterns[61433] = 29'b1_110111111111_001_1_111111110111;
      patterns[61434] = 29'b1_110111111111_010_1_101111111111;
      patterns[61435] = 29'b1_110111111111_011_1_011111111111;
      patterns[61436] = 29'b1_110111111111_100_1_111011111111;
      patterns[61437] = 29'b1_110111111111_101_1_111101111111;
      patterns[61438] = 29'b1_110111111111_110_1_110111111111;
      patterns[61439] = 29'b1_110111111111_111_1_110111111111;
      patterns[61440] = 29'b1_111000000000_000_1_111000000000;
      patterns[61441] = 29'b1_111000000000_001_1_000000111000;
      patterns[61442] = 29'b1_111000000000_010_1_110000000001;
      patterns[61443] = 29'b1_111000000000_011_1_100000000011;
      patterns[61444] = 29'b1_111000000000_100_0_111100000000;
      patterns[61445] = 29'b1_111000000000_101_0_011110000000;
      patterns[61446] = 29'b1_111000000000_110_1_111000000000;
      patterns[61447] = 29'b1_111000000000_111_1_111000000000;
      patterns[61448] = 29'b1_111000000001_000_1_111000000001;
      patterns[61449] = 29'b1_111000000001_001_1_000001111000;
      patterns[61450] = 29'b1_111000000001_010_1_110000000011;
      patterns[61451] = 29'b1_111000000001_011_1_100000000111;
      patterns[61452] = 29'b1_111000000001_100_1_111100000000;
      patterns[61453] = 29'b1_111000000001_101_0_111110000000;
      patterns[61454] = 29'b1_111000000001_110_1_111000000001;
      patterns[61455] = 29'b1_111000000001_111_1_111000000001;
      patterns[61456] = 29'b1_111000000010_000_1_111000000010;
      patterns[61457] = 29'b1_111000000010_001_1_000010111000;
      patterns[61458] = 29'b1_111000000010_010_1_110000000101;
      patterns[61459] = 29'b1_111000000010_011_1_100000001011;
      patterns[61460] = 29'b1_111000000010_100_0_111100000001;
      patterns[61461] = 29'b1_111000000010_101_1_011110000000;
      patterns[61462] = 29'b1_111000000010_110_1_111000000010;
      patterns[61463] = 29'b1_111000000010_111_1_111000000010;
      patterns[61464] = 29'b1_111000000011_000_1_111000000011;
      patterns[61465] = 29'b1_111000000011_001_1_000011111000;
      patterns[61466] = 29'b1_111000000011_010_1_110000000111;
      patterns[61467] = 29'b1_111000000011_011_1_100000001111;
      patterns[61468] = 29'b1_111000000011_100_1_111100000001;
      patterns[61469] = 29'b1_111000000011_101_1_111110000000;
      patterns[61470] = 29'b1_111000000011_110_1_111000000011;
      patterns[61471] = 29'b1_111000000011_111_1_111000000011;
      patterns[61472] = 29'b1_111000000100_000_1_111000000100;
      patterns[61473] = 29'b1_111000000100_001_1_000100111000;
      patterns[61474] = 29'b1_111000000100_010_1_110000001001;
      patterns[61475] = 29'b1_111000000100_011_1_100000010011;
      patterns[61476] = 29'b1_111000000100_100_0_111100000010;
      patterns[61477] = 29'b1_111000000100_101_0_011110000001;
      patterns[61478] = 29'b1_111000000100_110_1_111000000100;
      patterns[61479] = 29'b1_111000000100_111_1_111000000100;
      patterns[61480] = 29'b1_111000000101_000_1_111000000101;
      patterns[61481] = 29'b1_111000000101_001_1_000101111000;
      patterns[61482] = 29'b1_111000000101_010_1_110000001011;
      patterns[61483] = 29'b1_111000000101_011_1_100000010111;
      patterns[61484] = 29'b1_111000000101_100_1_111100000010;
      patterns[61485] = 29'b1_111000000101_101_0_111110000001;
      patterns[61486] = 29'b1_111000000101_110_1_111000000101;
      patterns[61487] = 29'b1_111000000101_111_1_111000000101;
      patterns[61488] = 29'b1_111000000110_000_1_111000000110;
      patterns[61489] = 29'b1_111000000110_001_1_000110111000;
      patterns[61490] = 29'b1_111000000110_010_1_110000001101;
      patterns[61491] = 29'b1_111000000110_011_1_100000011011;
      patterns[61492] = 29'b1_111000000110_100_0_111100000011;
      patterns[61493] = 29'b1_111000000110_101_1_011110000001;
      patterns[61494] = 29'b1_111000000110_110_1_111000000110;
      patterns[61495] = 29'b1_111000000110_111_1_111000000110;
      patterns[61496] = 29'b1_111000000111_000_1_111000000111;
      patterns[61497] = 29'b1_111000000111_001_1_000111111000;
      patterns[61498] = 29'b1_111000000111_010_1_110000001111;
      patterns[61499] = 29'b1_111000000111_011_1_100000011111;
      patterns[61500] = 29'b1_111000000111_100_1_111100000011;
      patterns[61501] = 29'b1_111000000111_101_1_111110000001;
      patterns[61502] = 29'b1_111000000111_110_1_111000000111;
      patterns[61503] = 29'b1_111000000111_111_1_111000000111;
      patterns[61504] = 29'b1_111000001000_000_1_111000001000;
      patterns[61505] = 29'b1_111000001000_001_1_001000111000;
      patterns[61506] = 29'b1_111000001000_010_1_110000010001;
      patterns[61507] = 29'b1_111000001000_011_1_100000100011;
      patterns[61508] = 29'b1_111000001000_100_0_111100000100;
      patterns[61509] = 29'b1_111000001000_101_0_011110000010;
      patterns[61510] = 29'b1_111000001000_110_1_111000001000;
      patterns[61511] = 29'b1_111000001000_111_1_111000001000;
      patterns[61512] = 29'b1_111000001001_000_1_111000001001;
      patterns[61513] = 29'b1_111000001001_001_1_001001111000;
      patterns[61514] = 29'b1_111000001001_010_1_110000010011;
      patterns[61515] = 29'b1_111000001001_011_1_100000100111;
      patterns[61516] = 29'b1_111000001001_100_1_111100000100;
      patterns[61517] = 29'b1_111000001001_101_0_111110000010;
      patterns[61518] = 29'b1_111000001001_110_1_111000001001;
      patterns[61519] = 29'b1_111000001001_111_1_111000001001;
      patterns[61520] = 29'b1_111000001010_000_1_111000001010;
      patterns[61521] = 29'b1_111000001010_001_1_001010111000;
      patterns[61522] = 29'b1_111000001010_010_1_110000010101;
      patterns[61523] = 29'b1_111000001010_011_1_100000101011;
      patterns[61524] = 29'b1_111000001010_100_0_111100000101;
      patterns[61525] = 29'b1_111000001010_101_1_011110000010;
      patterns[61526] = 29'b1_111000001010_110_1_111000001010;
      patterns[61527] = 29'b1_111000001010_111_1_111000001010;
      patterns[61528] = 29'b1_111000001011_000_1_111000001011;
      patterns[61529] = 29'b1_111000001011_001_1_001011111000;
      patterns[61530] = 29'b1_111000001011_010_1_110000010111;
      patterns[61531] = 29'b1_111000001011_011_1_100000101111;
      patterns[61532] = 29'b1_111000001011_100_1_111100000101;
      patterns[61533] = 29'b1_111000001011_101_1_111110000010;
      patterns[61534] = 29'b1_111000001011_110_1_111000001011;
      patterns[61535] = 29'b1_111000001011_111_1_111000001011;
      patterns[61536] = 29'b1_111000001100_000_1_111000001100;
      patterns[61537] = 29'b1_111000001100_001_1_001100111000;
      patterns[61538] = 29'b1_111000001100_010_1_110000011001;
      patterns[61539] = 29'b1_111000001100_011_1_100000110011;
      patterns[61540] = 29'b1_111000001100_100_0_111100000110;
      patterns[61541] = 29'b1_111000001100_101_0_011110000011;
      patterns[61542] = 29'b1_111000001100_110_1_111000001100;
      patterns[61543] = 29'b1_111000001100_111_1_111000001100;
      patterns[61544] = 29'b1_111000001101_000_1_111000001101;
      patterns[61545] = 29'b1_111000001101_001_1_001101111000;
      patterns[61546] = 29'b1_111000001101_010_1_110000011011;
      patterns[61547] = 29'b1_111000001101_011_1_100000110111;
      patterns[61548] = 29'b1_111000001101_100_1_111100000110;
      patterns[61549] = 29'b1_111000001101_101_0_111110000011;
      patterns[61550] = 29'b1_111000001101_110_1_111000001101;
      patterns[61551] = 29'b1_111000001101_111_1_111000001101;
      patterns[61552] = 29'b1_111000001110_000_1_111000001110;
      patterns[61553] = 29'b1_111000001110_001_1_001110111000;
      patterns[61554] = 29'b1_111000001110_010_1_110000011101;
      patterns[61555] = 29'b1_111000001110_011_1_100000111011;
      patterns[61556] = 29'b1_111000001110_100_0_111100000111;
      patterns[61557] = 29'b1_111000001110_101_1_011110000011;
      patterns[61558] = 29'b1_111000001110_110_1_111000001110;
      patterns[61559] = 29'b1_111000001110_111_1_111000001110;
      patterns[61560] = 29'b1_111000001111_000_1_111000001111;
      patterns[61561] = 29'b1_111000001111_001_1_001111111000;
      patterns[61562] = 29'b1_111000001111_010_1_110000011111;
      patterns[61563] = 29'b1_111000001111_011_1_100000111111;
      patterns[61564] = 29'b1_111000001111_100_1_111100000111;
      patterns[61565] = 29'b1_111000001111_101_1_111110000011;
      patterns[61566] = 29'b1_111000001111_110_1_111000001111;
      patterns[61567] = 29'b1_111000001111_111_1_111000001111;
      patterns[61568] = 29'b1_111000010000_000_1_111000010000;
      patterns[61569] = 29'b1_111000010000_001_1_010000111000;
      patterns[61570] = 29'b1_111000010000_010_1_110000100001;
      patterns[61571] = 29'b1_111000010000_011_1_100001000011;
      patterns[61572] = 29'b1_111000010000_100_0_111100001000;
      patterns[61573] = 29'b1_111000010000_101_0_011110000100;
      patterns[61574] = 29'b1_111000010000_110_1_111000010000;
      patterns[61575] = 29'b1_111000010000_111_1_111000010000;
      patterns[61576] = 29'b1_111000010001_000_1_111000010001;
      patterns[61577] = 29'b1_111000010001_001_1_010001111000;
      patterns[61578] = 29'b1_111000010001_010_1_110000100011;
      patterns[61579] = 29'b1_111000010001_011_1_100001000111;
      patterns[61580] = 29'b1_111000010001_100_1_111100001000;
      patterns[61581] = 29'b1_111000010001_101_0_111110000100;
      patterns[61582] = 29'b1_111000010001_110_1_111000010001;
      patterns[61583] = 29'b1_111000010001_111_1_111000010001;
      patterns[61584] = 29'b1_111000010010_000_1_111000010010;
      patterns[61585] = 29'b1_111000010010_001_1_010010111000;
      patterns[61586] = 29'b1_111000010010_010_1_110000100101;
      patterns[61587] = 29'b1_111000010010_011_1_100001001011;
      patterns[61588] = 29'b1_111000010010_100_0_111100001001;
      patterns[61589] = 29'b1_111000010010_101_1_011110000100;
      patterns[61590] = 29'b1_111000010010_110_1_111000010010;
      patterns[61591] = 29'b1_111000010010_111_1_111000010010;
      patterns[61592] = 29'b1_111000010011_000_1_111000010011;
      patterns[61593] = 29'b1_111000010011_001_1_010011111000;
      patterns[61594] = 29'b1_111000010011_010_1_110000100111;
      patterns[61595] = 29'b1_111000010011_011_1_100001001111;
      patterns[61596] = 29'b1_111000010011_100_1_111100001001;
      patterns[61597] = 29'b1_111000010011_101_1_111110000100;
      patterns[61598] = 29'b1_111000010011_110_1_111000010011;
      patterns[61599] = 29'b1_111000010011_111_1_111000010011;
      patterns[61600] = 29'b1_111000010100_000_1_111000010100;
      patterns[61601] = 29'b1_111000010100_001_1_010100111000;
      patterns[61602] = 29'b1_111000010100_010_1_110000101001;
      patterns[61603] = 29'b1_111000010100_011_1_100001010011;
      patterns[61604] = 29'b1_111000010100_100_0_111100001010;
      patterns[61605] = 29'b1_111000010100_101_0_011110000101;
      patterns[61606] = 29'b1_111000010100_110_1_111000010100;
      patterns[61607] = 29'b1_111000010100_111_1_111000010100;
      patterns[61608] = 29'b1_111000010101_000_1_111000010101;
      patterns[61609] = 29'b1_111000010101_001_1_010101111000;
      patterns[61610] = 29'b1_111000010101_010_1_110000101011;
      patterns[61611] = 29'b1_111000010101_011_1_100001010111;
      patterns[61612] = 29'b1_111000010101_100_1_111100001010;
      patterns[61613] = 29'b1_111000010101_101_0_111110000101;
      patterns[61614] = 29'b1_111000010101_110_1_111000010101;
      patterns[61615] = 29'b1_111000010101_111_1_111000010101;
      patterns[61616] = 29'b1_111000010110_000_1_111000010110;
      patterns[61617] = 29'b1_111000010110_001_1_010110111000;
      patterns[61618] = 29'b1_111000010110_010_1_110000101101;
      patterns[61619] = 29'b1_111000010110_011_1_100001011011;
      patterns[61620] = 29'b1_111000010110_100_0_111100001011;
      patterns[61621] = 29'b1_111000010110_101_1_011110000101;
      patterns[61622] = 29'b1_111000010110_110_1_111000010110;
      patterns[61623] = 29'b1_111000010110_111_1_111000010110;
      patterns[61624] = 29'b1_111000010111_000_1_111000010111;
      patterns[61625] = 29'b1_111000010111_001_1_010111111000;
      patterns[61626] = 29'b1_111000010111_010_1_110000101111;
      patterns[61627] = 29'b1_111000010111_011_1_100001011111;
      patterns[61628] = 29'b1_111000010111_100_1_111100001011;
      patterns[61629] = 29'b1_111000010111_101_1_111110000101;
      patterns[61630] = 29'b1_111000010111_110_1_111000010111;
      patterns[61631] = 29'b1_111000010111_111_1_111000010111;
      patterns[61632] = 29'b1_111000011000_000_1_111000011000;
      patterns[61633] = 29'b1_111000011000_001_1_011000111000;
      patterns[61634] = 29'b1_111000011000_010_1_110000110001;
      patterns[61635] = 29'b1_111000011000_011_1_100001100011;
      patterns[61636] = 29'b1_111000011000_100_0_111100001100;
      patterns[61637] = 29'b1_111000011000_101_0_011110000110;
      patterns[61638] = 29'b1_111000011000_110_1_111000011000;
      patterns[61639] = 29'b1_111000011000_111_1_111000011000;
      patterns[61640] = 29'b1_111000011001_000_1_111000011001;
      patterns[61641] = 29'b1_111000011001_001_1_011001111000;
      patterns[61642] = 29'b1_111000011001_010_1_110000110011;
      patterns[61643] = 29'b1_111000011001_011_1_100001100111;
      patterns[61644] = 29'b1_111000011001_100_1_111100001100;
      patterns[61645] = 29'b1_111000011001_101_0_111110000110;
      patterns[61646] = 29'b1_111000011001_110_1_111000011001;
      patterns[61647] = 29'b1_111000011001_111_1_111000011001;
      patterns[61648] = 29'b1_111000011010_000_1_111000011010;
      patterns[61649] = 29'b1_111000011010_001_1_011010111000;
      patterns[61650] = 29'b1_111000011010_010_1_110000110101;
      patterns[61651] = 29'b1_111000011010_011_1_100001101011;
      patterns[61652] = 29'b1_111000011010_100_0_111100001101;
      patterns[61653] = 29'b1_111000011010_101_1_011110000110;
      patterns[61654] = 29'b1_111000011010_110_1_111000011010;
      patterns[61655] = 29'b1_111000011010_111_1_111000011010;
      patterns[61656] = 29'b1_111000011011_000_1_111000011011;
      patterns[61657] = 29'b1_111000011011_001_1_011011111000;
      patterns[61658] = 29'b1_111000011011_010_1_110000110111;
      patterns[61659] = 29'b1_111000011011_011_1_100001101111;
      patterns[61660] = 29'b1_111000011011_100_1_111100001101;
      patterns[61661] = 29'b1_111000011011_101_1_111110000110;
      patterns[61662] = 29'b1_111000011011_110_1_111000011011;
      patterns[61663] = 29'b1_111000011011_111_1_111000011011;
      patterns[61664] = 29'b1_111000011100_000_1_111000011100;
      patterns[61665] = 29'b1_111000011100_001_1_011100111000;
      patterns[61666] = 29'b1_111000011100_010_1_110000111001;
      patterns[61667] = 29'b1_111000011100_011_1_100001110011;
      patterns[61668] = 29'b1_111000011100_100_0_111100001110;
      patterns[61669] = 29'b1_111000011100_101_0_011110000111;
      patterns[61670] = 29'b1_111000011100_110_1_111000011100;
      patterns[61671] = 29'b1_111000011100_111_1_111000011100;
      patterns[61672] = 29'b1_111000011101_000_1_111000011101;
      patterns[61673] = 29'b1_111000011101_001_1_011101111000;
      patterns[61674] = 29'b1_111000011101_010_1_110000111011;
      patterns[61675] = 29'b1_111000011101_011_1_100001110111;
      patterns[61676] = 29'b1_111000011101_100_1_111100001110;
      patterns[61677] = 29'b1_111000011101_101_0_111110000111;
      patterns[61678] = 29'b1_111000011101_110_1_111000011101;
      patterns[61679] = 29'b1_111000011101_111_1_111000011101;
      patterns[61680] = 29'b1_111000011110_000_1_111000011110;
      patterns[61681] = 29'b1_111000011110_001_1_011110111000;
      patterns[61682] = 29'b1_111000011110_010_1_110000111101;
      patterns[61683] = 29'b1_111000011110_011_1_100001111011;
      patterns[61684] = 29'b1_111000011110_100_0_111100001111;
      patterns[61685] = 29'b1_111000011110_101_1_011110000111;
      patterns[61686] = 29'b1_111000011110_110_1_111000011110;
      patterns[61687] = 29'b1_111000011110_111_1_111000011110;
      patterns[61688] = 29'b1_111000011111_000_1_111000011111;
      patterns[61689] = 29'b1_111000011111_001_1_011111111000;
      patterns[61690] = 29'b1_111000011111_010_1_110000111111;
      patterns[61691] = 29'b1_111000011111_011_1_100001111111;
      patterns[61692] = 29'b1_111000011111_100_1_111100001111;
      patterns[61693] = 29'b1_111000011111_101_1_111110000111;
      patterns[61694] = 29'b1_111000011111_110_1_111000011111;
      patterns[61695] = 29'b1_111000011111_111_1_111000011111;
      patterns[61696] = 29'b1_111000100000_000_1_111000100000;
      patterns[61697] = 29'b1_111000100000_001_1_100000111000;
      patterns[61698] = 29'b1_111000100000_010_1_110001000001;
      patterns[61699] = 29'b1_111000100000_011_1_100010000011;
      patterns[61700] = 29'b1_111000100000_100_0_111100010000;
      patterns[61701] = 29'b1_111000100000_101_0_011110001000;
      patterns[61702] = 29'b1_111000100000_110_1_111000100000;
      patterns[61703] = 29'b1_111000100000_111_1_111000100000;
      patterns[61704] = 29'b1_111000100001_000_1_111000100001;
      patterns[61705] = 29'b1_111000100001_001_1_100001111000;
      patterns[61706] = 29'b1_111000100001_010_1_110001000011;
      patterns[61707] = 29'b1_111000100001_011_1_100010000111;
      patterns[61708] = 29'b1_111000100001_100_1_111100010000;
      patterns[61709] = 29'b1_111000100001_101_0_111110001000;
      patterns[61710] = 29'b1_111000100001_110_1_111000100001;
      patterns[61711] = 29'b1_111000100001_111_1_111000100001;
      patterns[61712] = 29'b1_111000100010_000_1_111000100010;
      patterns[61713] = 29'b1_111000100010_001_1_100010111000;
      patterns[61714] = 29'b1_111000100010_010_1_110001000101;
      patterns[61715] = 29'b1_111000100010_011_1_100010001011;
      patterns[61716] = 29'b1_111000100010_100_0_111100010001;
      patterns[61717] = 29'b1_111000100010_101_1_011110001000;
      patterns[61718] = 29'b1_111000100010_110_1_111000100010;
      patterns[61719] = 29'b1_111000100010_111_1_111000100010;
      patterns[61720] = 29'b1_111000100011_000_1_111000100011;
      patterns[61721] = 29'b1_111000100011_001_1_100011111000;
      patterns[61722] = 29'b1_111000100011_010_1_110001000111;
      patterns[61723] = 29'b1_111000100011_011_1_100010001111;
      patterns[61724] = 29'b1_111000100011_100_1_111100010001;
      patterns[61725] = 29'b1_111000100011_101_1_111110001000;
      patterns[61726] = 29'b1_111000100011_110_1_111000100011;
      patterns[61727] = 29'b1_111000100011_111_1_111000100011;
      patterns[61728] = 29'b1_111000100100_000_1_111000100100;
      patterns[61729] = 29'b1_111000100100_001_1_100100111000;
      patterns[61730] = 29'b1_111000100100_010_1_110001001001;
      patterns[61731] = 29'b1_111000100100_011_1_100010010011;
      patterns[61732] = 29'b1_111000100100_100_0_111100010010;
      patterns[61733] = 29'b1_111000100100_101_0_011110001001;
      patterns[61734] = 29'b1_111000100100_110_1_111000100100;
      patterns[61735] = 29'b1_111000100100_111_1_111000100100;
      patterns[61736] = 29'b1_111000100101_000_1_111000100101;
      patterns[61737] = 29'b1_111000100101_001_1_100101111000;
      patterns[61738] = 29'b1_111000100101_010_1_110001001011;
      patterns[61739] = 29'b1_111000100101_011_1_100010010111;
      patterns[61740] = 29'b1_111000100101_100_1_111100010010;
      patterns[61741] = 29'b1_111000100101_101_0_111110001001;
      patterns[61742] = 29'b1_111000100101_110_1_111000100101;
      patterns[61743] = 29'b1_111000100101_111_1_111000100101;
      patterns[61744] = 29'b1_111000100110_000_1_111000100110;
      patterns[61745] = 29'b1_111000100110_001_1_100110111000;
      patterns[61746] = 29'b1_111000100110_010_1_110001001101;
      patterns[61747] = 29'b1_111000100110_011_1_100010011011;
      patterns[61748] = 29'b1_111000100110_100_0_111100010011;
      patterns[61749] = 29'b1_111000100110_101_1_011110001001;
      patterns[61750] = 29'b1_111000100110_110_1_111000100110;
      patterns[61751] = 29'b1_111000100110_111_1_111000100110;
      patterns[61752] = 29'b1_111000100111_000_1_111000100111;
      patterns[61753] = 29'b1_111000100111_001_1_100111111000;
      patterns[61754] = 29'b1_111000100111_010_1_110001001111;
      patterns[61755] = 29'b1_111000100111_011_1_100010011111;
      patterns[61756] = 29'b1_111000100111_100_1_111100010011;
      patterns[61757] = 29'b1_111000100111_101_1_111110001001;
      patterns[61758] = 29'b1_111000100111_110_1_111000100111;
      patterns[61759] = 29'b1_111000100111_111_1_111000100111;
      patterns[61760] = 29'b1_111000101000_000_1_111000101000;
      patterns[61761] = 29'b1_111000101000_001_1_101000111000;
      patterns[61762] = 29'b1_111000101000_010_1_110001010001;
      patterns[61763] = 29'b1_111000101000_011_1_100010100011;
      patterns[61764] = 29'b1_111000101000_100_0_111100010100;
      patterns[61765] = 29'b1_111000101000_101_0_011110001010;
      patterns[61766] = 29'b1_111000101000_110_1_111000101000;
      patterns[61767] = 29'b1_111000101000_111_1_111000101000;
      patterns[61768] = 29'b1_111000101001_000_1_111000101001;
      patterns[61769] = 29'b1_111000101001_001_1_101001111000;
      patterns[61770] = 29'b1_111000101001_010_1_110001010011;
      patterns[61771] = 29'b1_111000101001_011_1_100010100111;
      patterns[61772] = 29'b1_111000101001_100_1_111100010100;
      patterns[61773] = 29'b1_111000101001_101_0_111110001010;
      patterns[61774] = 29'b1_111000101001_110_1_111000101001;
      patterns[61775] = 29'b1_111000101001_111_1_111000101001;
      patterns[61776] = 29'b1_111000101010_000_1_111000101010;
      patterns[61777] = 29'b1_111000101010_001_1_101010111000;
      patterns[61778] = 29'b1_111000101010_010_1_110001010101;
      patterns[61779] = 29'b1_111000101010_011_1_100010101011;
      patterns[61780] = 29'b1_111000101010_100_0_111100010101;
      patterns[61781] = 29'b1_111000101010_101_1_011110001010;
      patterns[61782] = 29'b1_111000101010_110_1_111000101010;
      patterns[61783] = 29'b1_111000101010_111_1_111000101010;
      patterns[61784] = 29'b1_111000101011_000_1_111000101011;
      patterns[61785] = 29'b1_111000101011_001_1_101011111000;
      patterns[61786] = 29'b1_111000101011_010_1_110001010111;
      patterns[61787] = 29'b1_111000101011_011_1_100010101111;
      patterns[61788] = 29'b1_111000101011_100_1_111100010101;
      patterns[61789] = 29'b1_111000101011_101_1_111110001010;
      patterns[61790] = 29'b1_111000101011_110_1_111000101011;
      patterns[61791] = 29'b1_111000101011_111_1_111000101011;
      patterns[61792] = 29'b1_111000101100_000_1_111000101100;
      patterns[61793] = 29'b1_111000101100_001_1_101100111000;
      patterns[61794] = 29'b1_111000101100_010_1_110001011001;
      patterns[61795] = 29'b1_111000101100_011_1_100010110011;
      patterns[61796] = 29'b1_111000101100_100_0_111100010110;
      patterns[61797] = 29'b1_111000101100_101_0_011110001011;
      patterns[61798] = 29'b1_111000101100_110_1_111000101100;
      patterns[61799] = 29'b1_111000101100_111_1_111000101100;
      patterns[61800] = 29'b1_111000101101_000_1_111000101101;
      patterns[61801] = 29'b1_111000101101_001_1_101101111000;
      patterns[61802] = 29'b1_111000101101_010_1_110001011011;
      patterns[61803] = 29'b1_111000101101_011_1_100010110111;
      patterns[61804] = 29'b1_111000101101_100_1_111100010110;
      patterns[61805] = 29'b1_111000101101_101_0_111110001011;
      patterns[61806] = 29'b1_111000101101_110_1_111000101101;
      patterns[61807] = 29'b1_111000101101_111_1_111000101101;
      patterns[61808] = 29'b1_111000101110_000_1_111000101110;
      patterns[61809] = 29'b1_111000101110_001_1_101110111000;
      patterns[61810] = 29'b1_111000101110_010_1_110001011101;
      patterns[61811] = 29'b1_111000101110_011_1_100010111011;
      patterns[61812] = 29'b1_111000101110_100_0_111100010111;
      patterns[61813] = 29'b1_111000101110_101_1_011110001011;
      patterns[61814] = 29'b1_111000101110_110_1_111000101110;
      patterns[61815] = 29'b1_111000101110_111_1_111000101110;
      patterns[61816] = 29'b1_111000101111_000_1_111000101111;
      patterns[61817] = 29'b1_111000101111_001_1_101111111000;
      patterns[61818] = 29'b1_111000101111_010_1_110001011111;
      patterns[61819] = 29'b1_111000101111_011_1_100010111111;
      patterns[61820] = 29'b1_111000101111_100_1_111100010111;
      patterns[61821] = 29'b1_111000101111_101_1_111110001011;
      patterns[61822] = 29'b1_111000101111_110_1_111000101111;
      patterns[61823] = 29'b1_111000101111_111_1_111000101111;
      patterns[61824] = 29'b1_111000110000_000_1_111000110000;
      patterns[61825] = 29'b1_111000110000_001_1_110000111000;
      patterns[61826] = 29'b1_111000110000_010_1_110001100001;
      patterns[61827] = 29'b1_111000110000_011_1_100011000011;
      patterns[61828] = 29'b1_111000110000_100_0_111100011000;
      patterns[61829] = 29'b1_111000110000_101_0_011110001100;
      patterns[61830] = 29'b1_111000110000_110_1_111000110000;
      patterns[61831] = 29'b1_111000110000_111_1_111000110000;
      patterns[61832] = 29'b1_111000110001_000_1_111000110001;
      patterns[61833] = 29'b1_111000110001_001_1_110001111000;
      patterns[61834] = 29'b1_111000110001_010_1_110001100011;
      patterns[61835] = 29'b1_111000110001_011_1_100011000111;
      patterns[61836] = 29'b1_111000110001_100_1_111100011000;
      patterns[61837] = 29'b1_111000110001_101_0_111110001100;
      patterns[61838] = 29'b1_111000110001_110_1_111000110001;
      patterns[61839] = 29'b1_111000110001_111_1_111000110001;
      patterns[61840] = 29'b1_111000110010_000_1_111000110010;
      patterns[61841] = 29'b1_111000110010_001_1_110010111000;
      patterns[61842] = 29'b1_111000110010_010_1_110001100101;
      patterns[61843] = 29'b1_111000110010_011_1_100011001011;
      patterns[61844] = 29'b1_111000110010_100_0_111100011001;
      patterns[61845] = 29'b1_111000110010_101_1_011110001100;
      patterns[61846] = 29'b1_111000110010_110_1_111000110010;
      patterns[61847] = 29'b1_111000110010_111_1_111000110010;
      patterns[61848] = 29'b1_111000110011_000_1_111000110011;
      patterns[61849] = 29'b1_111000110011_001_1_110011111000;
      patterns[61850] = 29'b1_111000110011_010_1_110001100111;
      patterns[61851] = 29'b1_111000110011_011_1_100011001111;
      patterns[61852] = 29'b1_111000110011_100_1_111100011001;
      patterns[61853] = 29'b1_111000110011_101_1_111110001100;
      patterns[61854] = 29'b1_111000110011_110_1_111000110011;
      patterns[61855] = 29'b1_111000110011_111_1_111000110011;
      patterns[61856] = 29'b1_111000110100_000_1_111000110100;
      patterns[61857] = 29'b1_111000110100_001_1_110100111000;
      patterns[61858] = 29'b1_111000110100_010_1_110001101001;
      patterns[61859] = 29'b1_111000110100_011_1_100011010011;
      patterns[61860] = 29'b1_111000110100_100_0_111100011010;
      patterns[61861] = 29'b1_111000110100_101_0_011110001101;
      patterns[61862] = 29'b1_111000110100_110_1_111000110100;
      patterns[61863] = 29'b1_111000110100_111_1_111000110100;
      patterns[61864] = 29'b1_111000110101_000_1_111000110101;
      patterns[61865] = 29'b1_111000110101_001_1_110101111000;
      patterns[61866] = 29'b1_111000110101_010_1_110001101011;
      patterns[61867] = 29'b1_111000110101_011_1_100011010111;
      patterns[61868] = 29'b1_111000110101_100_1_111100011010;
      patterns[61869] = 29'b1_111000110101_101_0_111110001101;
      patterns[61870] = 29'b1_111000110101_110_1_111000110101;
      patterns[61871] = 29'b1_111000110101_111_1_111000110101;
      patterns[61872] = 29'b1_111000110110_000_1_111000110110;
      patterns[61873] = 29'b1_111000110110_001_1_110110111000;
      patterns[61874] = 29'b1_111000110110_010_1_110001101101;
      patterns[61875] = 29'b1_111000110110_011_1_100011011011;
      patterns[61876] = 29'b1_111000110110_100_0_111100011011;
      patterns[61877] = 29'b1_111000110110_101_1_011110001101;
      patterns[61878] = 29'b1_111000110110_110_1_111000110110;
      patterns[61879] = 29'b1_111000110110_111_1_111000110110;
      patterns[61880] = 29'b1_111000110111_000_1_111000110111;
      patterns[61881] = 29'b1_111000110111_001_1_110111111000;
      patterns[61882] = 29'b1_111000110111_010_1_110001101111;
      patterns[61883] = 29'b1_111000110111_011_1_100011011111;
      patterns[61884] = 29'b1_111000110111_100_1_111100011011;
      patterns[61885] = 29'b1_111000110111_101_1_111110001101;
      patterns[61886] = 29'b1_111000110111_110_1_111000110111;
      patterns[61887] = 29'b1_111000110111_111_1_111000110111;
      patterns[61888] = 29'b1_111000111000_000_1_111000111000;
      patterns[61889] = 29'b1_111000111000_001_1_111000111000;
      patterns[61890] = 29'b1_111000111000_010_1_110001110001;
      patterns[61891] = 29'b1_111000111000_011_1_100011100011;
      patterns[61892] = 29'b1_111000111000_100_0_111100011100;
      patterns[61893] = 29'b1_111000111000_101_0_011110001110;
      patterns[61894] = 29'b1_111000111000_110_1_111000111000;
      patterns[61895] = 29'b1_111000111000_111_1_111000111000;
      patterns[61896] = 29'b1_111000111001_000_1_111000111001;
      patterns[61897] = 29'b1_111000111001_001_1_111001111000;
      patterns[61898] = 29'b1_111000111001_010_1_110001110011;
      patterns[61899] = 29'b1_111000111001_011_1_100011100111;
      patterns[61900] = 29'b1_111000111001_100_1_111100011100;
      patterns[61901] = 29'b1_111000111001_101_0_111110001110;
      patterns[61902] = 29'b1_111000111001_110_1_111000111001;
      patterns[61903] = 29'b1_111000111001_111_1_111000111001;
      patterns[61904] = 29'b1_111000111010_000_1_111000111010;
      patterns[61905] = 29'b1_111000111010_001_1_111010111000;
      patterns[61906] = 29'b1_111000111010_010_1_110001110101;
      patterns[61907] = 29'b1_111000111010_011_1_100011101011;
      patterns[61908] = 29'b1_111000111010_100_0_111100011101;
      patterns[61909] = 29'b1_111000111010_101_1_011110001110;
      patterns[61910] = 29'b1_111000111010_110_1_111000111010;
      patterns[61911] = 29'b1_111000111010_111_1_111000111010;
      patterns[61912] = 29'b1_111000111011_000_1_111000111011;
      patterns[61913] = 29'b1_111000111011_001_1_111011111000;
      patterns[61914] = 29'b1_111000111011_010_1_110001110111;
      patterns[61915] = 29'b1_111000111011_011_1_100011101111;
      patterns[61916] = 29'b1_111000111011_100_1_111100011101;
      patterns[61917] = 29'b1_111000111011_101_1_111110001110;
      patterns[61918] = 29'b1_111000111011_110_1_111000111011;
      patterns[61919] = 29'b1_111000111011_111_1_111000111011;
      patterns[61920] = 29'b1_111000111100_000_1_111000111100;
      patterns[61921] = 29'b1_111000111100_001_1_111100111000;
      patterns[61922] = 29'b1_111000111100_010_1_110001111001;
      patterns[61923] = 29'b1_111000111100_011_1_100011110011;
      patterns[61924] = 29'b1_111000111100_100_0_111100011110;
      patterns[61925] = 29'b1_111000111100_101_0_011110001111;
      patterns[61926] = 29'b1_111000111100_110_1_111000111100;
      patterns[61927] = 29'b1_111000111100_111_1_111000111100;
      patterns[61928] = 29'b1_111000111101_000_1_111000111101;
      patterns[61929] = 29'b1_111000111101_001_1_111101111000;
      patterns[61930] = 29'b1_111000111101_010_1_110001111011;
      patterns[61931] = 29'b1_111000111101_011_1_100011110111;
      patterns[61932] = 29'b1_111000111101_100_1_111100011110;
      patterns[61933] = 29'b1_111000111101_101_0_111110001111;
      patterns[61934] = 29'b1_111000111101_110_1_111000111101;
      patterns[61935] = 29'b1_111000111101_111_1_111000111101;
      patterns[61936] = 29'b1_111000111110_000_1_111000111110;
      patterns[61937] = 29'b1_111000111110_001_1_111110111000;
      patterns[61938] = 29'b1_111000111110_010_1_110001111101;
      patterns[61939] = 29'b1_111000111110_011_1_100011111011;
      patterns[61940] = 29'b1_111000111110_100_0_111100011111;
      patterns[61941] = 29'b1_111000111110_101_1_011110001111;
      patterns[61942] = 29'b1_111000111110_110_1_111000111110;
      patterns[61943] = 29'b1_111000111110_111_1_111000111110;
      patterns[61944] = 29'b1_111000111111_000_1_111000111111;
      patterns[61945] = 29'b1_111000111111_001_1_111111111000;
      patterns[61946] = 29'b1_111000111111_010_1_110001111111;
      patterns[61947] = 29'b1_111000111111_011_1_100011111111;
      patterns[61948] = 29'b1_111000111111_100_1_111100011111;
      patterns[61949] = 29'b1_111000111111_101_1_111110001111;
      patterns[61950] = 29'b1_111000111111_110_1_111000111111;
      patterns[61951] = 29'b1_111000111111_111_1_111000111111;
      patterns[61952] = 29'b1_111001000000_000_1_111001000000;
      patterns[61953] = 29'b1_111001000000_001_1_000000111001;
      patterns[61954] = 29'b1_111001000000_010_1_110010000001;
      patterns[61955] = 29'b1_111001000000_011_1_100100000011;
      patterns[61956] = 29'b1_111001000000_100_0_111100100000;
      patterns[61957] = 29'b1_111001000000_101_0_011110010000;
      patterns[61958] = 29'b1_111001000000_110_1_111001000000;
      patterns[61959] = 29'b1_111001000000_111_1_111001000000;
      patterns[61960] = 29'b1_111001000001_000_1_111001000001;
      patterns[61961] = 29'b1_111001000001_001_1_000001111001;
      patterns[61962] = 29'b1_111001000001_010_1_110010000011;
      patterns[61963] = 29'b1_111001000001_011_1_100100000111;
      patterns[61964] = 29'b1_111001000001_100_1_111100100000;
      patterns[61965] = 29'b1_111001000001_101_0_111110010000;
      patterns[61966] = 29'b1_111001000001_110_1_111001000001;
      patterns[61967] = 29'b1_111001000001_111_1_111001000001;
      patterns[61968] = 29'b1_111001000010_000_1_111001000010;
      patterns[61969] = 29'b1_111001000010_001_1_000010111001;
      patterns[61970] = 29'b1_111001000010_010_1_110010000101;
      patterns[61971] = 29'b1_111001000010_011_1_100100001011;
      patterns[61972] = 29'b1_111001000010_100_0_111100100001;
      patterns[61973] = 29'b1_111001000010_101_1_011110010000;
      patterns[61974] = 29'b1_111001000010_110_1_111001000010;
      patterns[61975] = 29'b1_111001000010_111_1_111001000010;
      patterns[61976] = 29'b1_111001000011_000_1_111001000011;
      patterns[61977] = 29'b1_111001000011_001_1_000011111001;
      patterns[61978] = 29'b1_111001000011_010_1_110010000111;
      patterns[61979] = 29'b1_111001000011_011_1_100100001111;
      patterns[61980] = 29'b1_111001000011_100_1_111100100001;
      patterns[61981] = 29'b1_111001000011_101_1_111110010000;
      patterns[61982] = 29'b1_111001000011_110_1_111001000011;
      patterns[61983] = 29'b1_111001000011_111_1_111001000011;
      patterns[61984] = 29'b1_111001000100_000_1_111001000100;
      patterns[61985] = 29'b1_111001000100_001_1_000100111001;
      patterns[61986] = 29'b1_111001000100_010_1_110010001001;
      patterns[61987] = 29'b1_111001000100_011_1_100100010011;
      patterns[61988] = 29'b1_111001000100_100_0_111100100010;
      patterns[61989] = 29'b1_111001000100_101_0_011110010001;
      patterns[61990] = 29'b1_111001000100_110_1_111001000100;
      patterns[61991] = 29'b1_111001000100_111_1_111001000100;
      patterns[61992] = 29'b1_111001000101_000_1_111001000101;
      patterns[61993] = 29'b1_111001000101_001_1_000101111001;
      patterns[61994] = 29'b1_111001000101_010_1_110010001011;
      patterns[61995] = 29'b1_111001000101_011_1_100100010111;
      patterns[61996] = 29'b1_111001000101_100_1_111100100010;
      patterns[61997] = 29'b1_111001000101_101_0_111110010001;
      patterns[61998] = 29'b1_111001000101_110_1_111001000101;
      patterns[61999] = 29'b1_111001000101_111_1_111001000101;
      patterns[62000] = 29'b1_111001000110_000_1_111001000110;
      patterns[62001] = 29'b1_111001000110_001_1_000110111001;
      patterns[62002] = 29'b1_111001000110_010_1_110010001101;
      patterns[62003] = 29'b1_111001000110_011_1_100100011011;
      patterns[62004] = 29'b1_111001000110_100_0_111100100011;
      patterns[62005] = 29'b1_111001000110_101_1_011110010001;
      patterns[62006] = 29'b1_111001000110_110_1_111001000110;
      patterns[62007] = 29'b1_111001000110_111_1_111001000110;
      patterns[62008] = 29'b1_111001000111_000_1_111001000111;
      patterns[62009] = 29'b1_111001000111_001_1_000111111001;
      patterns[62010] = 29'b1_111001000111_010_1_110010001111;
      patterns[62011] = 29'b1_111001000111_011_1_100100011111;
      patterns[62012] = 29'b1_111001000111_100_1_111100100011;
      patterns[62013] = 29'b1_111001000111_101_1_111110010001;
      patterns[62014] = 29'b1_111001000111_110_1_111001000111;
      patterns[62015] = 29'b1_111001000111_111_1_111001000111;
      patterns[62016] = 29'b1_111001001000_000_1_111001001000;
      patterns[62017] = 29'b1_111001001000_001_1_001000111001;
      patterns[62018] = 29'b1_111001001000_010_1_110010010001;
      patterns[62019] = 29'b1_111001001000_011_1_100100100011;
      patterns[62020] = 29'b1_111001001000_100_0_111100100100;
      patterns[62021] = 29'b1_111001001000_101_0_011110010010;
      patterns[62022] = 29'b1_111001001000_110_1_111001001000;
      patterns[62023] = 29'b1_111001001000_111_1_111001001000;
      patterns[62024] = 29'b1_111001001001_000_1_111001001001;
      patterns[62025] = 29'b1_111001001001_001_1_001001111001;
      patterns[62026] = 29'b1_111001001001_010_1_110010010011;
      patterns[62027] = 29'b1_111001001001_011_1_100100100111;
      patterns[62028] = 29'b1_111001001001_100_1_111100100100;
      patterns[62029] = 29'b1_111001001001_101_0_111110010010;
      patterns[62030] = 29'b1_111001001001_110_1_111001001001;
      patterns[62031] = 29'b1_111001001001_111_1_111001001001;
      patterns[62032] = 29'b1_111001001010_000_1_111001001010;
      patterns[62033] = 29'b1_111001001010_001_1_001010111001;
      patterns[62034] = 29'b1_111001001010_010_1_110010010101;
      patterns[62035] = 29'b1_111001001010_011_1_100100101011;
      patterns[62036] = 29'b1_111001001010_100_0_111100100101;
      patterns[62037] = 29'b1_111001001010_101_1_011110010010;
      patterns[62038] = 29'b1_111001001010_110_1_111001001010;
      patterns[62039] = 29'b1_111001001010_111_1_111001001010;
      patterns[62040] = 29'b1_111001001011_000_1_111001001011;
      patterns[62041] = 29'b1_111001001011_001_1_001011111001;
      patterns[62042] = 29'b1_111001001011_010_1_110010010111;
      patterns[62043] = 29'b1_111001001011_011_1_100100101111;
      patterns[62044] = 29'b1_111001001011_100_1_111100100101;
      patterns[62045] = 29'b1_111001001011_101_1_111110010010;
      patterns[62046] = 29'b1_111001001011_110_1_111001001011;
      patterns[62047] = 29'b1_111001001011_111_1_111001001011;
      patterns[62048] = 29'b1_111001001100_000_1_111001001100;
      patterns[62049] = 29'b1_111001001100_001_1_001100111001;
      patterns[62050] = 29'b1_111001001100_010_1_110010011001;
      patterns[62051] = 29'b1_111001001100_011_1_100100110011;
      patterns[62052] = 29'b1_111001001100_100_0_111100100110;
      patterns[62053] = 29'b1_111001001100_101_0_011110010011;
      patterns[62054] = 29'b1_111001001100_110_1_111001001100;
      patterns[62055] = 29'b1_111001001100_111_1_111001001100;
      patterns[62056] = 29'b1_111001001101_000_1_111001001101;
      patterns[62057] = 29'b1_111001001101_001_1_001101111001;
      patterns[62058] = 29'b1_111001001101_010_1_110010011011;
      patterns[62059] = 29'b1_111001001101_011_1_100100110111;
      patterns[62060] = 29'b1_111001001101_100_1_111100100110;
      patterns[62061] = 29'b1_111001001101_101_0_111110010011;
      patterns[62062] = 29'b1_111001001101_110_1_111001001101;
      patterns[62063] = 29'b1_111001001101_111_1_111001001101;
      patterns[62064] = 29'b1_111001001110_000_1_111001001110;
      patterns[62065] = 29'b1_111001001110_001_1_001110111001;
      patterns[62066] = 29'b1_111001001110_010_1_110010011101;
      patterns[62067] = 29'b1_111001001110_011_1_100100111011;
      patterns[62068] = 29'b1_111001001110_100_0_111100100111;
      patterns[62069] = 29'b1_111001001110_101_1_011110010011;
      patterns[62070] = 29'b1_111001001110_110_1_111001001110;
      patterns[62071] = 29'b1_111001001110_111_1_111001001110;
      patterns[62072] = 29'b1_111001001111_000_1_111001001111;
      patterns[62073] = 29'b1_111001001111_001_1_001111111001;
      patterns[62074] = 29'b1_111001001111_010_1_110010011111;
      patterns[62075] = 29'b1_111001001111_011_1_100100111111;
      patterns[62076] = 29'b1_111001001111_100_1_111100100111;
      patterns[62077] = 29'b1_111001001111_101_1_111110010011;
      patterns[62078] = 29'b1_111001001111_110_1_111001001111;
      patterns[62079] = 29'b1_111001001111_111_1_111001001111;
      patterns[62080] = 29'b1_111001010000_000_1_111001010000;
      patterns[62081] = 29'b1_111001010000_001_1_010000111001;
      patterns[62082] = 29'b1_111001010000_010_1_110010100001;
      patterns[62083] = 29'b1_111001010000_011_1_100101000011;
      patterns[62084] = 29'b1_111001010000_100_0_111100101000;
      patterns[62085] = 29'b1_111001010000_101_0_011110010100;
      patterns[62086] = 29'b1_111001010000_110_1_111001010000;
      patterns[62087] = 29'b1_111001010000_111_1_111001010000;
      patterns[62088] = 29'b1_111001010001_000_1_111001010001;
      patterns[62089] = 29'b1_111001010001_001_1_010001111001;
      patterns[62090] = 29'b1_111001010001_010_1_110010100011;
      patterns[62091] = 29'b1_111001010001_011_1_100101000111;
      patterns[62092] = 29'b1_111001010001_100_1_111100101000;
      patterns[62093] = 29'b1_111001010001_101_0_111110010100;
      patterns[62094] = 29'b1_111001010001_110_1_111001010001;
      patterns[62095] = 29'b1_111001010001_111_1_111001010001;
      patterns[62096] = 29'b1_111001010010_000_1_111001010010;
      patterns[62097] = 29'b1_111001010010_001_1_010010111001;
      patterns[62098] = 29'b1_111001010010_010_1_110010100101;
      patterns[62099] = 29'b1_111001010010_011_1_100101001011;
      patterns[62100] = 29'b1_111001010010_100_0_111100101001;
      patterns[62101] = 29'b1_111001010010_101_1_011110010100;
      patterns[62102] = 29'b1_111001010010_110_1_111001010010;
      patterns[62103] = 29'b1_111001010010_111_1_111001010010;
      patterns[62104] = 29'b1_111001010011_000_1_111001010011;
      patterns[62105] = 29'b1_111001010011_001_1_010011111001;
      patterns[62106] = 29'b1_111001010011_010_1_110010100111;
      patterns[62107] = 29'b1_111001010011_011_1_100101001111;
      patterns[62108] = 29'b1_111001010011_100_1_111100101001;
      patterns[62109] = 29'b1_111001010011_101_1_111110010100;
      patterns[62110] = 29'b1_111001010011_110_1_111001010011;
      patterns[62111] = 29'b1_111001010011_111_1_111001010011;
      patterns[62112] = 29'b1_111001010100_000_1_111001010100;
      patterns[62113] = 29'b1_111001010100_001_1_010100111001;
      patterns[62114] = 29'b1_111001010100_010_1_110010101001;
      patterns[62115] = 29'b1_111001010100_011_1_100101010011;
      patterns[62116] = 29'b1_111001010100_100_0_111100101010;
      patterns[62117] = 29'b1_111001010100_101_0_011110010101;
      patterns[62118] = 29'b1_111001010100_110_1_111001010100;
      patterns[62119] = 29'b1_111001010100_111_1_111001010100;
      patterns[62120] = 29'b1_111001010101_000_1_111001010101;
      patterns[62121] = 29'b1_111001010101_001_1_010101111001;
      patterns[62122] = 29'b1_111001010101_010_1_110010101011;
      patterns[62123] = 29'b1_111001010101_011_1_100101010111;
      patterns[62124] = 29'b1_111001010101_100_1_111100101010;
      patterns[62125] = 29'b1_111001010101_101_0_111110010101;
      patterns[62126] = 29'b1_111001010101_110_1_111001010101;
      patterns[62127] = 29'b1_111001010101_111_1_111001010101;
      patterns[62128] = 29'b1_111001010110_000_1_111001010110;
      patterns[62129] = 29'b1_111001010110_001_1_010110111001;
      patterns[62130] = 29'b1_111001010110_010_1_110010101101;
      patterns[62131] = 29'b1_111001010110_011_1_100101011011;
      patterns[62132] = 29'b1_111001010110_100_0_111100101011;
      patterns[62133] = 29'b1_111001010110_101_1_011110010101;
      patterns[62134] = 29'b1_111001010110_110_1_111001010110;
      patterns[62135] = 29'b1_111001010110_111_1_111001010110;
      patterns[62136] = 29'b1_111001010111_000_1_111001010111;
      patterns[62137] = 29'b1_111001010111_001_1_010111111001;
      patterns[62138] = 29'b1_111001010111_010_1_110010101111;
      patterns[62139] = 29'b1_111001010111_011_1_100101011111;
      patterns[62140] = 29'b1_111001010111_100_1_111100101011;
      patterns[62141] = 29'b1_111001010111_101_1_111110010101;
      patterns[62142] = 29'b1_111001010111_110_1_111001010111;
      patterns[62143] = 29'b1_111001010111_111_1_111001010111;
      patterns[62144] = 29'b1_111001011000_000_1_111001011000;
      patterns[62145] = 29'b1_111001011000_001_1_011000111001;
      patterns[62146] = 29'b1_111001011000_010_1_110010110001;
      patterns[62147] = 29'b1_111001011000_011_1_100101100011;
      patterns[62148] = 29'b1_111001011000_100_0_111100101100;
      patterns[62149] = 29'b1_111001011000_101_0_011110010110;
      patterns[62150] = 29'b1_111001011000_110_1_111001011000;
      patterns[62151] = 29'b1_111001011000_111_1_111001011000;
      patterns[62152] = 29'b1_111001011001_000_1_111001011001;
      patterns[62153] = 29'b1_111001011001_001_1_011001111001;
      patterns[62154] = 29'b1_111001011001_010_1_110010110011;
      patterns[62155] = 29'b1_111001011001_011_1_100101100111;
      patterns[62156] = 29'b1_111001011001_100_1_111100101100;
      patterns[62157] = 29'b1_111001011001_101_0_111110010110;
      patterns[62158] = 29'b1_111001011001_110_1_111001011001;
      patterns[62159] = 29'b1_111001011001_111_1_111001011001;
      patterns[62160] = 29'b1_111001011010_000_1_111001011010;
      patterns[62161] = 29'b1_111001011010_001_1_011010111001;
      patterns[62162] = 29'b1_111001011010_010_1_110010110101;
      patterns[62163] = 29'b1_111001011010_011_1_100101101011;
      patterns[62164] = 29'b1_111001011010_100_0_111100101101;
      patterns[62165] = 29'b1_111001011010_101_1_011110010110;
      patterns[62166] = 29'b1_111001011010_110_1_111001011010;
      patterns[62167] = 29'b1_111001011010_111_1_111001011010;
      patterns[62168] = 29'b1_111001011011_000_1_111001011011;
      patterns[62169] = 29'b1_111001011011_001_1_011011111001;
      patterns[62170] = 29'b1_111001011011_010_1_110010110111;
      patterns[62171] = 29'b1_111001011011_011_1_100101101111;
      patterns[62172] = 29'b1_111001011011_100_1_111100101101;
      patterns[62173] = 29'b1_111001011011_101_1_111110010110;
      patterns[62174] = 29'b1_111001011011_110_1_111001011011;
      patterns[62175] = 29'b1_111001011011_111_1_111001011011;
      patterns[62176] = 29'b1_111001011100_000_1_111001011100;
      patterns[62177] = 29'b1_111001011100_001_1_011100111001;
      patterns[62178] = 29'b1_111001011100_010_1_110010111001;
      patterns[62179] = 29'b1_111001011100_011_1_100101110011;
      patterns[62180] = 29'b1_111001011100_100_0_111100101110;
      patterns[62181] = 29'b1_111001011100_101_0_011110010111;
      patterns[62182] = 29'b1_111001011100_110_1_111001011100;
      patterns[62183] = 29'b1_111001011100_111_1_111001011100;
      patterns[62184] = 29'b1_111001011101_000_1_111001011101;
      patterns[62185] = 29'b1_111001011101_001_1_011101111001;
      patterns[62186] = 29'b1_111001011101_010_1_110010111011;
      patterns[62187] = 29'b1_111001011101_011_1_100101110111;
      patterns[62188] = 29'b1_111001011101_100_1_111100101110;
      patterns[62189] = 29'b1_111001011101_101_0_111110010111;
      patterns[62190] = 29'b1_111001011101_110_1_111001011101;
      patterns[62191] = 29'b1_111001011101_111_1_111001011101;
      patterns[62192] = 29'b1_111001011110_000_1_111001011110;
      patterns[62193] = 29'b1_111001011110_001_1_011110111001;
      patterns[62194] = 29'b1_111001011110_010_1_110010111101;
      patterns[62195] = 29'b1_111001011110_011_1_100101111011;
      patterns[62196] = 29'b1_111001011110_100_0_111100101111;
      patterns[62197] = 29'b1_111001011110_101_1_011110010111;
      patterns[62198] = 29'b1_111001011110_110_1_111001011110;
      patterns[62199] = 29'b1_111001011110_111_1_111001011110;
      patterns[62200] = 29'b1_111001011111_000_1_111001011111;
      patterns[62201] = 29'b1_111001011111_001_1_011111111001;
      patterns[62202] = 29'b1_111001011111_010_1_110010111111;
      patterns[62203] = 29'b1_111001011111_011_1_100101111111;
      patterns[62204] = 29'b1_111001011111_100_1_111100101111;
      patterns[62205] = 29'b1_111001011111_101_1_111110010111;
      patterns[62206] = 29'b1_111001011111_110_1_111001011111;
      patterns[62207] = 29'b1_111001011111_111_1_111001011111;
      patterns[62208] = 29'b1_111001100000_000_1_111001100000;
      patterns[62209] = 29'b1_111001100000_001_1_100000111001;
      patterns[62210] = 29'b1_111001100000_010_1_110011000001;
      patterns[62211] = 29'b1_111001100000_011_1_100110000011;
      patterns[62212] = 29'b1_111001100000_100_0_111100110000;
      patterns[62213] = 29'b1_111001100000_101_0_011110011000;
      patterns[62214] = 29'b1_111001100000_110_1_111001100000;
      patterns[62215] = 29'b1_111001100000_111_1_111001100000;
      patterns[62216] = 29'b1_111001100001_000_1_111001100001;
      patterns[62217] = 29'b1_111001100001_001_1_100001111001;
      patterns[62218] = 29'b1_111001100001_010_1_110011000011;
      patterns[62219] = 29'b1_111001100001_011_1_100110000111;
      patterns[62220] = 29'b1_111001100001_100_1_111100110000;
      patterns[62221] = 29'b1_111001100001_101_0_111110011000;
      patterns[62222] = 29'b1_111001100001_110_1_111001100001;
      patterns[62223] = 29'b1_111001100001_111_1_111001100001;
      patterns[62224] = 29'b1_111001100010_000_1_111001100010;
      patterns[62225] = 29'b1_111001100010_001_1_100010111001;
      patterns[62226] = 29'b1_111001100010_010_1_110011000101;
      patterns[62227] = 29'b1_111001100010_011_1_100110001011;
      patterns[62228] = 29'b1_111001100010_100_0_111100110001;
      patterns[62229] = 29'b1_111001100010_101_1_011110011000;
      patterns[62230] = 29'b1_111001100010_110_1_111001100010;
      patterns[62231] = 29'b1_111001100010_111_1_111001100010;
      patterns[62232] = 29'b1_111001100011_000_1_111001100011;
      patterns[62233] = 29'b1_111001100011_001_1_100011111001;
      patterns[62234] = 29'b1_111001100011_010_1_110011000111;
      patterns[62235] = 29'b1_111001100011_011_1_100110001111;
      patterns[62236] = 29'b1_111001100011_100_1_111100110001;
      patterns[62237] = 29'b1_111001100011_101_1_111110011000;
      patterns[62238] = 29'b1_111001100011_110_1_111001100011;
      patterns[62239] = 29'b1_111001100011_111_1_111001100011;
      patterns[62240] = 29'b1_111001100100_000_1_111001100100;
      patterns[62241] = 29'b1_111001100100_001_1_100100111001;
      patterns[62242] = 29'b1_111001100100_010_1_110011001001;
      patterns[62243] = 29'b1_111001100100_011_1_100110010011;
      patterns[62244] = 29'b1_111001100100_100_0_111100110010;
      patterns[62245] = 29'b1_111001100100_101_0_011110011001;
      patterns[62246] = 29'b1_111001100100_110_1_111001100100;
      patterns[62247] = 29'b1_111001100100_111_1_111001100100;
      patterns[62248] = 29'b1_111001100101_000_1_111001100101;
      patterns[62249] = 29'b1_111001100101_001_1_100101111001;
      patterns[62250] = 29'b1_111001100101_010_1_110011001011;
      patterns[62251] = 29'b1_111001100101_011_1_100110010111;
      patterns[62252] = 29'b1_111001100101_100_1_111100110010;
      patterns[62253] = 29'b1_111001100101_101_0_111110011001;
      patterns[62254] = 29'b1_111001100101_110_1_111001100101;
      patterns[62255] = 29'b1_111001100101_111_1_111001100101;
      patterns[62256] = 29'b1_111001100110_000_1_111001100110;
      patterns[62257] = 29'b1_111001100110_001_1_100110111001;
      patterns[62258] = 29'b1_111001100110_010_1_110011001101;
      patterns[62259] = 29'b1_111001100110_011_1_100110011011;
      patterns[62260] = 29'b1_111001100110_100_0_111100110011;
      patterns[62261] = 29'b1_111001100110_101_1_011110011001;
      patterns[62262] = 29'b1_111001100110_110_1_111001100110;
      patterns[62263] = 29'b1_111001100110_111_1_111001100110;
      patterns[62264] = 29'b1_111001100111_000_1_111001100111;
      patterns[62265] = 29'b1_111001100111_001_1_100111111001;
      patterns[62266] = 29'b1_111001100111_010_1_110011001111;
      patterns[62267] = 29'b1_111001100111_011_1_100110011111;
      patterns[62268] = 29'b1_111001100111_100_1_111100110011;
      patterns[62269] = 29'b1_111001100111_101_1_111110011001;
      patterns[62270] = 29'b1_111001100111_110_1_111001100111;
      patterns[62271] = 29'b1_111001100111_111_1_111001100111;
      patterns[62272] = 29'b1_111001101000_000_1_111001101000;
      patterns[62273] = 29'b1_111001101000_001_1_101000111001;
      patterns[62274] = 29'b1_111001101000_010_1_110011010001;
      patterns[62275] = 29'b1_111001101000_011_1_100110100011;
      patterns[62276] = 29'b1_111001101000_100_0_111100110100;
      patterns[62277] = 29'b1_111001101000_101_0_011110011010;
      patterns[62278] = 29'b1_111001101000_110_1_111001101000;
      patterns[62279] = 29'b1_111001101000_111_1_111001101000;
      patterns[62280] = 29'b1_111001101001_000_1_111001101001;
      patterns[62281] = 29'b1_111001101001_001_1_101001111001;
      patterns[62282] = 29'b1_111001101001_010_1_110011010011;
      patterns[62283] = 29'b1_111001101001_011_1_100110100111;
      patterns[62284] = 29'b1_111001101001_100_1_111100110100;
      patterns[62285] = 29'b1_111001101001_101_0_111110011010;
      patterns[62286] = 29'b1_111001101001_110_1_111001101001;
      patterns[62287] = 29'b1_111001101001_111_1_111001101001;
      patterns[62288] = 29'b1_111001101010_000_1_111001101010;
      patterns[62289] = 29'b1_111001101010_001_1_101010111001;
      patterns[62290] = 29'b1_111001101010_010_1_110011010101;
      patterns[62291] = 29'b1_111001101010_011_1_100110101011;
      patterns[62292] = 29'b1_111001101010_100_0_111100110101;
      patterns[62293] = 29'b1_111001101010_101_1_011110011010;
      patterns[62294] = 29'b1_111001101010_110_1_111001101010;
      patterns[62295] = 29'b1_111001101010_111_1_111001101010;
      patterns[62296] = 29'b1_111001101011_000_1_111001101011;
      patterns[62297] = 29'b1_111001101011_001_1_101011111001;
      patterns[62298] = 29'b1_111001101011_010_1_110011010111;
      patterns[62299] = 29'b1_111001101011_011_1_100110101111;
      patterns[62300] = 29'b1_111001101011_100_1_111100110101;
      patterns[62301] = 29'b1_111001101011_101_1_111110011010;
      patterns[62302] = 29'b1_111001101011_110_1_111001101011;
      patterns[62303] = 29'b1_111001101011_111_1_111001101011;
      patterns[62304] = 29'b1_111001101100_000_1_111001101100;
      patterns[62305] = 29'b1_111001101100_001_1_101100111001;
      patterns[62306] = 29'b1_111001101100_010_1_110011011001;
      patterns[62307] = 29'b1_111001101100_011_1_100110110011;
      patterns[62308] = 29'b1_111001101100_100_0_111100110110;
      patterns[62309] = 29'b1_111001101100_101_0_011110011011;
      patterns[62310] = 29'b1_111001101100_110_1_111001101100;
      patterns[62311] = 29'b1_111001101100_111_1_111001101100;
      patterns[62312] = 29'b1_111001101101_000_1_111001101101;
      patterns[62313] = 29'b1_111001101101_001_1_101101111001;
      patterns[62314] = 29'b1_111001101101_010_1_110011011011;
      patterns[62315] = 29'b1_111001101101_011_1_100110110111;
      patterns[62316] = 29'b1_111001101101_100_1_111100110110;
      patterns[62317] = 29'b1_111001101101_101_0_111110011011;
      patterns[62318] = 29'b1_111001101101_110_1_111001101101;
      patterns[62319] = 29'b1_111001101101_111_1_111001101101;
      patterns[62320] = 29'b1_111001101110_000_1_111001101110;
      patterns[62321] = 29'b1_111001101110_001_1_101110111001;
      patterns[62322] = 29'b1_111001101110_010_1_110011011101;
      patterns[62323] = 29'b1_111001101110_011_1_100110111011;
      patterns[62324] = 29'b1_111001101110_100_0_111100110111;
      patterns[62325] = 29'b1_111001101110_101_1_011110011011;
      patterns[62326] = 29'b1_111001101110_110_1_111001101110;
      patterns[62327] = 29'b1_111001101110_111_1_111001101110;
      patterns[62328] = 29'b1_111001101111_000_1_111001101111;
      patterns[62329] = 29'b1_111001101111_001_1_101111111001;
      patterns[62330] = 29'b1_111001101111_010_1_110011011111;
      patterns[62331] = 29'b1_111001101111_011_1_100110111111;
      patterns[62332] = 29'b1_111001101111_100_1_111100110111;
      patterns[62333] = 29'b1_111001101111_101_1_111110011011;
      patterns[62334] = 29'b1_111001101111_110_1_111001101111;
      patterns[62335] = 29'b1_111001101111_111_1_111001101111;
      patterns[62336] = 29'b1_111001110000_000_1_111001110000;
      patterns[62337] = 29'b1_111001110000_001_1_110000111001;
      patterns[62338] = 29'b1_111001110000_010_1_110011100001;
      patterns[62339] = 29'b1_111001110000_011_1_100111000011;
      patterns[62340] = 29'b1_111001110000_100_0_111100111000;
      patterns[62341] = 29'b1_111001110000_101_0_011110011100;
      patterns[62342] = 29'b1_111001110000_110_1_111001110000;
      patterns[62343] = 29'b1_111001110000_111_1_111001110000;
      patterns[62344] = 29'b1_111001110001_000_1_111001110001;
      patterns[62345] = 29'b1_111001110001_001_1_110001111001;
      patterns[62346] = 29'b1_111001110001_010_1_110011100011;
      patterns[62347] = 29'b1_111001110001_011_1_100111000111;
      patterns[62348] = 29'b1_111001110001_100_1_111100111000;
      patterns[62349] = 29'b1_111001110001_101_0_111110011100;
      patterns[62350] = 29'b1_111001110001_110_1_111001110001;
      patterns[62351] = 29'b1_111001110001_111_1_111001110001;
      patterns[62352] = 29'b1_111001110010_000_1_111001110010;
      patterns[62353] = 29'b1_111001110010_001_1_110010111001;
      patterns[62354] = 29'b1_111001110010_010_1_110011100101;
      patterns[62355] = 29'b1_111001110010_011_1_100111001011;
      patterns[62356] = 29'b1_111001110010_100_0_111100111001;
      patterns[62357] = 29'b1_111001110010_101_1_011110011100;
      patterns[62358] = 29'b1_111001110010_110_1_111001110010;
      patterns[62359] = 29'b1_111001110010_111_1_111001110010;
      patterns[62360] = 29'b1_111001110011_000_1_111001110011;
      patterns[62361] = 29'b1_111001110011_001_1_110011111001;
      patterns[62362] = 29'b1_111001110011_010_1_110011100111;
      patterns[62363] = 29'b1_111001110011_011_1_100111001111;
      patterns[62364] = 29'b1_111001110011_100_1_111100111001;
      patterns[62365] = 29'b1_111001110011_101_1_111110011100;
      patterns[62366] = 29'b1_111001110011_110_1_111001110011;
      patterns[62367] = 29'b1_111001110011_111_1_111001110011;
      patterns[62368] = 29'b1_111001110100_000_1_111001110100;
      patterns[62369] = 29'b1_111001110100_001_1_110100111001;
      patterns[62370] = 29'b1_111001110100_010_1_110011101001;
      patterns[62371] = 29'b1_111001110100_011_1_100111010011;
      patterns[62372] = 29'b1_111001110100_100_0_111100111010;
      patterns[62373] = 29'b1_111001110100_101_0_011110011101;
      patterns[62374] = 29'b1_111001110100_110_1_111001110100;
      patterns[62375] = 29'b1_111001110100_111_1_111001110100;
      patterns[62376] = 29'b1_111001110101_000_1_111001110101;
      patterns[62377] = 29'b1_111001110101_001_1_110101111001;
      patterns[62378] = 29'b1_111001110101_010_1_110011101011;
      patterns[62379] = 29'b1_111001110101_011_1_100111010111;
      patterns[62380] = 29'b1_111001110101_100_1_111100111010;
      patterns[62381] = 29'b1_111001110101_101_0_111110011101;
      patterns[62382] = 29'b1_111001110101_110_1_111001110101;
      patterns[62383] = 29'b1_111001110101_111_1_111001110101;
      patterns[62384] = 29'b1_111001110110_000_1_111001110110;
      patterns[62385] = 29'b1_111001110110_001_1_110110111001;
      patterns[62386] = 29'b1_111001110110_010_1_110011101101;
      patterns[62387] = 29'b1_111001110110_011_1_100111011011;
      patterns[62388] = 29'b1_111001110110_100_0_111100111011;
      patterns[62389] = 29'b1_111001110110_101_1_011110011101;
      patterns[62390] = 29'b1_111001110110_110_1_111001110110;
      patterns[62391] = 29'b1_111001110110_111_1_111001110110;
      patterns[62392] = 29'b1_111001110111_000_1_111001110111;
      patterns[62393] = 29'b1_111001110111_001_1_110111111001;
      patterns[62394] = 29'b1_111001110111_010_1_110011101111;
      patterns[62395] = 29'b1_111001110111_011_1_100111011111;
      patterns[62396] = 29'b1_111001110111_100_1_111100111011;
      patterns[62397] = 29'b1_111001110111_101_1_111110011101;
      patterns[62398] = 29'b1_111001110111_110_1_111001110111;
      patterns[62399] = 29'b1_111001110111_111_1_111001110111;
      patterns[62400] = 29'b1_111001111000_000_1_111001111000;
      patterns[62401] = 29'b1_111001111000_001_1_111000111001;
      patterns[62402] = 29'b1_111001111000_010_1_110011110001;
      patterns[62403] = 29'b1_111001111000_011_1_100111100011;
      patterns[62404] = 29'b1_111001111000_100_0_111100111100;
      patterns[62405] = 29'b1_111001111000_101_0_011110011110;
      patterns[62406] = 29'b1_111001111000_110_1_111001111000;
      patterns[62407] = 29'b1_111001111000_111_1_111001111000;
      patterns[62408] = 29'b1_111001111001_000_1_111001111001;
      patterns[62409] = 29'b1_111001111001_001_1_111001111001;
      patterns[62410] = 29'b1_111001111001_010_1_110011110011;
      patterns[62411] = 29'b1_111001111001_011_1_100111100111;
      patterns[62412] = 29'b1_111001111001_100_1_111100111100;
      patterns[62413] = 29'b1_111001111001_101_0_111110011110;
      patterns[62414] = 29'b1_111001111001_110_1_111001111001;
      patterns[62415] = 29'b1_111001111001_111_1_111001111001;
      patterns[62416] = 29'b1_111001111010_000_1_111001111010;
      patterns[62417] = 29'b1_111001111010_001_1_111010111001;
      patterns[62418] = 29'b1_111001111010_010_1_110011110101;
      patterns[62419] = 29'b1_111001111010_011_1_100111101011;
      patterns[62420] = 29'b1_111001111010_100_0_111100111101;
      patterns[62421] = 29'b1_111001111010_101_1_011110011110;
      patterns[62422] = 29'b1_111001111010_110_1_111001111010;
      patterns[62423] = 29'b1_111001111010_111_1_111001111010;
      patterns[62424] = 29'b1_111001111011_000_1_111001111011;
      patterns[62425] = 29'b1_111001111011_001_1_111011111001;
      patterns[62426] = 29'b1_111001111011_010_1_110011110111;
      patterns[62427] = 29'b1_111001111011_011_1_100111101111;
      patterns[62428] = 29'b1_111001111011_100_1_111100111101;
      patterns[62429] = 29'b1_111001111011_101_1_111110011110;
      patterns[62430] = 29'b1_111001111011_110_1_111001111011;
      patterns[62431] = 29'b1_111001111011_111_1_111001111011;
      patterns[62432] = 29'b1_111001111100_000_1_111001111100;
      patterns[62433] = 29'b1_111001111100_001_1_111100111001;
      patterns[62434] = 29'b1_111001111100_010_1_110011111001;
      patterns[62435] = 29'b1_111001111100_011_1_100111110011;
      patterns[62436] = 29'b1_111001111100_100_0_111100111110;
      patterns[62437] = 29'b1_111001111100_101_0_011110011111;
      patterns[62438] = 29'b1_111001111100_110_1_111001111100;
      patterns[62439] = 29'b1_111001111100_111_1_111001111100;
      patterns[62440] = 29'b1_111001111101_000_1_111001111101;
      patterns[62441] = 29'b1_111001111101_001_1_111101111001;
      patterns[62442] = 29'b1_111001111101_010_1_110011111011;
      patterns[62443] = 29'b1_111001111101_011_1_100111110111;
      patterns[62444] = 29'b1_111001111101_100_1_111100111110;
      patterns[62445] = 29'b1_111001111101_101_0_111110011111;
      patterns[62446] = 29'b1_111001111101_110_1_111001111101;
      patterns[62447] = 29'b1_111001111101_111_1_111001111101;
      patterns[62448] = 29'b1_111001111110_000_1_111001111110;
      patterns[62449] = 29'b1_111001111110_001_1_111110111001;
      patterns[62450] = 29'b1_111001111110_010_1_110011111101;
      patterns[62451] = 29'b1_111001111110_011_1_100111111011;
      patterns[62452] = 29'b1_111001111110_100_0_111100111111;
      patterns[62453] = 29'b1_111001111110_101_1_011110011111;
      patterns[62454] = 29'b1_111001111110_110_1_111001111110;
      patterns[62455] = 29'b1_111001111110_111_1_111001111110;
      patterns[62456] = 29'b1_111001111111_000_1_111001111111;
      patterns[62457] = 29'b1_111001111111_001_1_111111111001;
      patterns[62458] = 29'b1_111001111111_010_1_110011111111;
      patterns[62459] = 29'b1_111001111111_011_1_100111111111;
      patterns[62460] = 29'b1_111001111111_100_1_111100111111;
      patterns[62461] = 29'b1_111001111111_101_1_111110011111;
      patterns[62462] = 29'b1_111001111111_110_1_111001111111;
      patterns[62463] = 29'b1_111001111111_111_1_111001111111;
      patterns[62464] = 29'b1_111010000000_000_1_111010000000;
      patterns[62465] = 29'b1_111010000000_001_1_000000111010;
      patterns[62466] = 29'b1_111010000000_010_1_110100000001;
      patterns[62467] = 29'b1_111010000000_011_1_101000000011;
      patterns[62468] = 29'b1_111010000000_100_0_111101000000;
      patterns[62469] = 29'b1_111010000000_101_0_011110100000;
      patterns[62470] = 29'b1_111010000000_110_1_111010000000;
      patterns[62471] = 29'b1_111010000000_111_1_111010000000;
      patterns[62472] = 29'b1_111010000001_000_1_111010000001;
      patterns[62473] = 29'b1_111010000001_001_1_000001111010;
      patterns[62474] = 29'b1_111010000001_010_1_110100000011;
      patterns[62475] = 29'b1_111010000001_011_1_101000000111;
      patterns[62476] = 29'b1_111010000001_100_1_111101000000;
      patterns[62477] = 29'b1_111010000001_101_0_111110100000;
      patterns[62478] = 29'b1_111010000001_110_1_111010000001;
      patterns[62479] = 29'b1_111010000001_111_1_111010000001;
      patterns[62480] = 29'b1_111010000010_000_1_111010000010;
      patterns[62481] = 29'b1_111010000010_001_1_000010111010;
      patterns[62482] = 29'b1_111010000010_010_1_110100000101;
      patterns[62483] = 29'b1_111010000010_011_1_101000001011;
      patterns[62484] = 29'b1_111010000010_100_0_111101000001;
      patterns[62485] = 29'b1_111010000010_101_1_011110100000;
      patterns[62486] = 29'b1_111010000010_110_1_111010000010;
      patterns[62487] = 29'b1_111010000010_111_1_111010000010;
      patterns[62488] = 29'b1_111010000011_000_1_111010000011;
      patterns[62489] = 29'b1_111010000011_001_1_000011111010;
      patterns[62490] = 29'b1_111010000011_010_1_110100000111;
      patterns[62491] = 29'b1_111010000011_011_1_101000001111;
      patterns[62492] = 29'b1_111010000011_100_1_111101000001;
      patterns[62493] = 29'b1_111010000011_101_1_111110100000;
      patterns[62494] = 29'b1_111010000011_110_1_111010000011;
      patterns[62495] = 29'b1_111010000011_111_1_111010000011;
      patterns[62496] = 29'b1_111010000100_000_1_111010000100;
      patterns[62497] = 29'b1_111010000100_001_1_000100111010;
      patterns[62498] = 29'b1_111010000100_010_1_110100001001;
      patterns[62499] = 29'b1_111010000100_011_1_101000010011;
      patterns[62500] = 29'b1_111010000100_100_0_111101000010;
      patterns[62501] = 29'b1_111010000100_101_0_011110100001;
      patterns[62502] = 29'b1_111010000100_110_1_111010000100;
      patterns[62503] = 29'b1_111010000100_111_1_111010000100;
      patterns[62504] = 29'b1_111010000101_000_1_111010000101;
      patterns[62505] = 29'b1_111010000101_001_1_000101111010;
      patterns[62506] = 29'b1_111010000101_010_1_110100001011;
      patterns[62507] = 29'b1_111010000101_011_1_101000010111;
      patterns[62508] = 29'b1_111010000101_100_1_111101000010;
      patterns[62509] = 29'b1_111010000101_101_0_111110100001;
      patterns[62510] = 29'b1_111010000101_110_1_111010000101;
      patterns[62511] = 29'b1_111010000101_111_1_111010000101;
      patterns[62512] = 29'b1_111010000110_000_1_111010000110;
      patterns[62513] = 29'b1_111010000110_001_1_000110111010;
      patterns[62514] = 29'b1_111010000110_010_1_110100001101;
      patterns[62515] = 29'b1_111010000110_011_1_101000011011;
      patterns[62516] = 29'b1_111010000110_100_0_111101000011;
      patterns[62517] = 29'b1_111010000110_101_1_011110100001;
      patterns[62518] = 29'b1_111010000110_110_1_111010000110;
      patterns[62519] = 29'b1_111010000110_111_1_111010000110;
      patterns[62520] = 29'b1_111010000111_000_1_111010000111;
      patterns[62521] = 29'b1_111010000111_001_1_000111111010;
      patterns[62522] = 29'b1_111010000111_010_1_110100001111;
      patterns[62523] = 29'b1_111010000111_011_1_101000011111;
      patterns[62524] = 29'b1_111010000111_100_1_111101000011;
      patterns[62525] = 29'b1_111010000111_101_1_111110100001;
      patterns[62526] = 29'b1_111010000111_110_1_111010000111;
      patterns[62527] = 29'b1_111010000111_111_1_111010000111;
      patterns[62528] = 29'b1_111010001000_000_1_111010001000;
      patterns[62529] = 29'b1_111010001000_001_1_001000111010;
      patterns[62530] = 29'b1_111010001000_010_1_110100010001;
      patterns[62531] = 29'b1_111010001000_011_1_101000100011;
      patterns[62532] = 29'b1_111010001000_100_0_111101000100;
      patterns[62533] = 29'b1_111010001000_101_0_011110100010;
      patterns[62534] = 29'b1_111010001000_110_1_111010001000;
      patterns[62535] = 29'b1_111010001000_111_1_111010001000;
      patterns[62536] = 29'b1_111010001001_000_1_111010001001;
      patterns[62537] = 29'b1_111010001001_001_1_001001111010;
      patterns[62538] = 29'b1_111010001001_010_1_110100010011;
      patterns[62539] = 29'b1_111010001001_011_1_101000100111;
      patterns[62540] = 29'b1_111010001001_100_1_111101000100;
      patterns[62541] = 29'b1_111010001001_101_0_111110100010;
      patterns[62542] = 29'b1_111010001001_110_1_111010001001;
      patterns[62543] = 29'b1_111010001001_111_1_111010001001;
      patterns[62544] = 29'b1_111010001010_000_1_111010001010;
      patterns[62545] = 29'b1_111010001010_001_1_001010111010;
      patterns[62546] = 29'b1_111010001010_010_1_110100010101;
      patterns[62547] = 29'b1_111010001010_011_1_101000101011;
      patterns[62548] = 29'b1_111010001010_100_0_111101000101;
      patterns[62549] = 29'b1_111010001010_101_1_011110100010;
      patterns[62550] = 29'b1_111010001010_110_1_111010001010;
      patterns[62551] = 29'b1_111010001010_111_1_111010001010;
      patterns[62552] = 29'b1_111010001011_000_1_111010001011;
      patterns[62553] = 29'b1_111010001011_001_1_001011111010;
      patterns[62554] = 29'b1_111010001011_010_1_110100010111;
      patterns[62555] = 29'b1_111010001011_011_1_101000101111;
      patterns[62556] = 29'b1_111010001011_100_1_111101000101;
      patterns[62557] = 29'b1_111010001011_101_1_111110100010;
      patterns[62558] = 29'b1_111010001011_110_1_111010001011;
      patterns[62559] = 29'b1_111010001011_111_1_111010001011;
      patterns[62560] = 29'b1_111010001100_000_1_111010001100;
      patterns[62561] = 29'b1_111010001100_001_1_001100111010;
      patterns[62562] = 29'b1_111010001100_010_1_110100011001;
      patterns[62563] = 29'b1_111010001100_011_1_101000110011;
      patterns[62564] = 29'b1_111010001100_100_0_111101000110;
      patterns[62565] = 29'b1_111010001100_101_0_011110100011;
      patterns[62566] = 29'b1_111010001100_110_1_111010001100;
      patterns[62567] = 29'b1_111010001100_111_1_111010001100;
      patterns[62568] = 29'b1_111010001101_000_1_111010001101;
      patterns[62569] = 29'b1_111010001101_001_1_001101111010;
      patterns[62570] = 29'b1_111010001101_010_1_110100011011;
      patterns[62571] = 29'b1_111010001101_011_1_101000110111;
      patterns[62572] = 29'b1_111010001101_100_1_111101000110;
      patterns[62573] = 29'b1_111010001101_101_0_111110100011;
      patterns[62574] = 29'b1_111010001101_110_1_111010001101;
      patterns[62575] = 29'b1_111010001101_111_1_111010001101;
      patterns[62576] = 29'b1_111010001110_000_1_111010001110;
      patterns[62577] = 29'b1_111010001110_001_1_001110111010;
      patterns[62578] = 29'b1_111010001110_010_1_110100011101;
      patterns[62579] = 29'b1_111010001110_011_1_101000111011;
      patterns[62580] = 29'b1_111010001110_100_0_111101000111;
      patterns[62581] = 29'b1_111010001110_101_1_011110100011;
      patterns[62582] = 29'b1_111010001110_110_1_111010001110;
      patterns[62583] = 29'b1_111010001110_111_1_111010001110;
      patterns[62584] = 29'b1_111010001111_000_1_111010001111;
      patterns[62585] = 29'b1_111010001111_001_1_001111111010;
      patterns[62586] = 29'b1_111010001111_010_1_110100011111;
      patterns[62587] = 29'b1_111010001111_011_1_101000111111;
      patterns[62588] = 29'b1_111010001111_100_1_111101000111;
      patterns[62589] = 29'b1_111010001111_101_1_111110100011;
      patterns[62590] = 29'b1_111010001111_110_1_111010001111;
      patterns[62591] = 29'b1_111010001111_111_1_111010001111;
      patterns[62592] = 29'b1_111010010000_000_1_111010010000;
      patterns[62593] = 29'b1_111010010000_001_1_010000111010;
      patterns[62594] = 29'b1_111010010000_010_1_110100100001;
      patterns[62595] = 29'b1_111010010000_011_1_101001000011;
      patterns[62596] = 29'b1_111010010000_100_0_111101001000;
      patterns[62597] = 29'b1_111010010000_101_0_011110100100;
      patterns[62598] = 29'b1_111010010000_110_1_111010010000;
      patterns[62599] = 29'b1_111010010000_111_1_111010010000;
      patterns[62600] = 29'b1_111010010001_000_1_111010010001;
      patterns[62601] = 29'b1_111010010001_001_1_010001111010;
      patterns[62602] = 29'b1_111010010001_010_1_110100100011;
      patterns[62603] = 29'b1_111010010001_011_1_101001000111;
      patterns[62604] = 29'b1_111010010001_100_1_111101001000;
      patterns[62605] = 29'b1_111010010001_101_0_111110100100;
      patterns[62606] = 29'b1_111010010001_110_1_111010010001;
      patterns[62607] = 29'b1_111010010001_111_1_111010010001;
      patterns[62608] = 29'b1_111010010010_000_1_111010010010;
      patterns[62609] = 29'b1_111010010010_001_1_010010111010;
      patterns[62610] = 29'b1_111010010010_010_1_110100100101;
      patterns[62611] = 29'b1_111010010010_011_1_101001001011;
      patterns[62612] = 29'b1_111010010010_100_0_111101001001;
      patterns[62613] = 29'b1_111010010010_101_1_011110100100;
      patterns[62614] = 29'b1_111010010010_110_1_111010010010;
      patterns[62615] = 29'b1_111010010010_111_1_111010010010;
      patterns[62616] = 29'b1_111010010011_000_1_111010010011;
      patterns[62617] = 29'b1_111010010011_001_1_010011111010;
      patterns[62618] = 29'b1_111010010011_010_1_110100100111;
      patterns[62619] = 29'b1_111010010011_011_1_101001001111;
      patterns[62620] = 29'b1_111010010011_100_1_111101001001;
      patterns[62621] = 29'b1_111010010011_101_1_111110100100;
      patterns[62622] = 29'b1_111010010011_110_1_111010010011;
      patterns[62623] = 29'b1_111010010011_111_1_111010010011;
      patterns[62624] = 29'b1_111010010100_000_1_111010010100;
      patterns[62625] = 29'b1_111010010100_001_1_010100111010;
      patterns[62626] = 29'b1_111010010100_010_1_110100101001;
      patterns[62627] = 29'b1_111010010100_011_1_101001010011;
      patterns[62628] = 29'b1_111010010100_100_0_111101001010;
      patterns[62629] = 29'b1_111010010100_101_0_011110100101;
      patterns[62630] = 29'b1_111010010100_110_1_111010010100;
      patterns[62631] = 29'b1_111010010100_111_1_111010010100;
      patterns[62632] = 29'b1_111010010101_000_1_111010010101;
      patterns[62633] = 29'b1_111010010101_001_1_010101111010;
      patterns[62634] = 29'b1_111010010101_010_1_110100101011;
      patterns[62635] = 29'b1_111010010101_011_1_101001010111;
      patterns[62636] = 29'b1_111010010101_100_1_111101001010;
      patterns[62637] = 29'b1_111010010101_101_0_111110100101;
      patterns[62638] = 29'b1_111010010101_110_1_111010010101;
      patterns[62639] = 29'b1_111010010101_111_1_111010010101;
      patterns[62640] = 29'b1_111010010110_000_1_111010010110;
      patterns[62641] = 29'b1_111010010110_001_1_010110111010;
      patterns[62642] = 29'b1_111010010110_010_1_110100101101;
      patterns[62643] = 29'b1_111010010110_011_1_101001011011;
      patterns[62644] = 29'b1_111010010110_100_0_111101001011;
      patterns[62645] = 29'b1_111010010110_101_1_011110100101;
      patterns[62646] = 29'b1_111010010110_110_1_111010010110;
      patterns[62647] = 29'b1_111010010110_111_1_111010010110;
      patterns[62648] = 29'b1_111010010111_000_1_111010010111;
      patterns[62649] = 29'b1_111010010111_001_1_010111111010;
      patterns[62650] = 29'b1_111010010111_010_1_110100101111;
      patterns[62651] = 29'b1_111010010111_011_1_101001011111;
      patterns[62652] = 29'b1_111010010111_100_1_111101001011;
      patterns[62653] = 29'b1_111010010111_101_1_111110100101;
      patterns[62654] = 29'b1_111010010111_110_1_111010010111;
      patterns[62655] = 29'b1_111010010111_111_1_111010010111;
      patterns[62656] = 29'b1_111010011000_000_1_111010011000;
      patterns[62657] = 29'b1_111010011000_001_1_011000111010;
      patterns[62658] = 29'b1_111010011000_010_1_110100110001;
      patterns[62659] = 29'b1_111010011000_011_1_101001100011;
      patterns[62660] = 29'b1_111010011000_100_0_111101001100;
      patterns[62661] = 29'b1_111010011000_101_0_011110100110;
      patterns[62662] = 29'b1_111010011000_110_1_111010011000;
      patterns[62663] = 29'b1_111010011000_111_1_111010011000;
      patterns[62664] = 29'b1_111010011001_000_1_111010011001;
      patterns[62665] = 29'b1_111010011001_001_1_011001111010;
      patterns[62666] = 29'b1_111010011001_010_1_110100110011;
      patterns[62667] = 29'b1_111010011001_011_1_101001100111;
      patterns[62668] = 29'b1_111010011001_100_1_111101001100;
      patterns[62669] = 29'b1_111010011001_101_0_111110100110;
      patterns[62670] = 29'b1_111010011001_110_1_111010011001;
      patterns[62671] = 29'b1_111010011001_111_1_111010011001;
      patterns[62672] = 29'b1_111010011010_000_1_111010011010;
      patterns[62673] = 29'b1_111010011010_001_1_011010111010;
      patterns[62674] = 29'b1_111010011010_010_1_110100110101;
      patterns[62675] = 29'b1_111010011010_011_1_101001101011;
      patterns[62676] = 29'b1_111010011010_100_0_111101001101;
      patterns[62677] = 29'b1_111010011010_101_1_011110100110;
      patterns[62678] = 29'b1_111010011010_110_1_111010011010;
      patterns[62679] = 29'b1_111010011010_111_1_111010011010;
      patterns[62680] = 29'b1_111010011011_000_1_111010011011;
      patterns[62681] = 29'b1_111010011011_001_1_011011111010;
      patterns[62682] = 29'b1_111010011011_010_1_110100110111;
      patterns[62683] = 29'b1_111010011011_011_1_101001101111;
      patterns[62684] = 29'b1_111010011011_100_1_111101001101;
      patterns[62685] = 29'b1_111010011011_101_1_111110100110;
      patterns[62686] = 29'b1_111010011011_110_1_111010011011;
      patterns[62687] = 29'b1_111010011011_111_1_111010011011;
      patterns[62688] = 29'b1_111010011100_000_1_111010011100;
      patterns[62689] = 29'b1_111010011100_001_1_011100111010;
      patterns[62690] = 29'b1_111010011100_010_1_110100111001;
      patterns[62691] = 29'b1_111010011100_011_1_101001110011;
      patterns[62692] = 29'b1_111010011100_100_0_111101001110;
      patterns[62693] = 29'b1_111010011100_101_0_011110100111;
      patterns[62694] = 29'b1_111010011100_110_1_111010011100;
      patterns[62695] = 29'b1_111010011100_111_1_111010011100;
      patterns[62696] = 29'b1_111010011101_000_1_111010011101;
      patterns[62697] = 29'b1_111010011101_001_1_011101111010;
      patterns[62698] = 29'b1_111010011101_010_1_110100111011;
      patterns[62699] = 29'b1_111010011101_011_1_101001110111;
      patterns[62700] = 29'b1_111010011101_100_1_111101001110;
      patterns[62701] = 29'b1_111010011101_101_0_111110100111;
      patterns[62702] = 29'b1_111010011101_110_1_111010011101;
      patterns[62703] = 29'b1_111010011101_111_1_111010011101;
      patterns[62704] = 29'b1_111010011110_000_1_111010011110;
      patterns[62705] = 29'b1_111010011110_001_1_011110111010;
      patterns[62706] = 29'b1_111010011110_010_1_110100111101;
      patterns[62707] = 29'b1_111010011110_011_1_101001111011;
      patterns[62708] = 29'b1_111010011110_100_0_111101001111;
      patterns[62709] = 29'b1_111010011110_101_1_011110100111;
      patterns[62710] = 29'b1_111010011110_110_1_111010011110;
      patterns[62711] = 29'b1_111010011110_111_1_111010011110;
      patterns[62712] = 29'b1_111010011111_000_1_111010011111;
      patterns[62713] = 29'b1_111010011111_001_1_011111111010;
      patterns[62714] = 29'b1_111010011111_010_1_110100111111;
      patterns[62715] = 29'b1_111010011111_011_1_101001111111;
      patterns[62716] = 29'b1_111010011111_100_1_111101001111;
      patterns[62717] = 29'b1_111010011111_101_1_111110100111;
      patterns[62718] = 29'b1_111010011111_110_1_111010011111;
      patterns[62719] = 29'b1_111010011111_111_1_111010011111;
      patterns[62720] = 29'b1_111010100000_000_1_111010100000;
      patterns[62721] = 29'b1_111010100000_001_1_100000111010;
      patterns[62722] = 29'b1_111010100000_010_1_110101000001;
      patterns[62723] = 29'b1_111010100000_011_1_101010000011;
      patterns[62724] = 29'b1_111010100000_100_0_111101010000;
      patterns[62725] = 29'b1_111010100000_101_0_011110101000;
      patterns[62726] = 29'b1_111010100000_110_1_111010100000;
      patterns[62727] = 29'b1_111010100000_111_1_111010100000;
      patterns[62728] = 29'b1_111010100001_000_1_111010100001;
      patterns[62729] = 29'b1_111010100001_001_1_100001111010;
      patterns[62730] = 29'b1_111010100001_010_1_110101000011;
      patterns[62731] = 29'b1_111010100001_011_1_101010000111;
      patterns[62732] = 29'b1_111010100001_100_1_111101010000;
      patterns[62733] = 29'b1_111010100001_101_0_111110101000;
      patterns[62734] = 29'b1_111010100001_110_1_111010100001;
      patterns[62735] = 29'b1_111010100001_111_1_111010100001;
      patterns[62736] = 29'b1_111010100010_000_1_111010100010;
      patterns[62737] = 29'b1_111010100010_001_1_100010111010;
      patterns[62738] = 29'b1_111010100010_010_1_110101000101;
      patterns[62739] = 29'b1_111010100010_011_1_101010001011;
      patterns[62740] = 29'b1_111010100010_100_0_111101010001;
      patterns[62741] = 29'b1_111010100010_101_1_011110101000;
      patterns[62742] = 29'b1_111010100010_110_1_111010100010;
      patterns[62743] = 29'b1_111010100010_111_1_111010100010;
      patterns[62744] = 29'b1_111010100011_000_1_111010100011;
      patterns[62745] = 29'b1_111010100011_001_1_100011111010;
      patterns[62746] = 29'b1_111010100011_010_1_110101000111;
      patterns[62747] = 29'b1_111010100011_011_1_101010001111;
      patterns[62748] = 29'b1_111010100011_100_1_111101010001;
      patterns[62749] = 29'b1_111010100011_101_1_111110101000;
      patterns[62750] = 29'b1_111010100011_110_1_111010100011;
      patterns[62751] = 29'b1_111010100011_111_1_111010100011;
      patterns[62752] = 29'b1_111010100100_000_1_111010100100;
      patterns[62753] = 29'b1_111010100100_001_1_100100111010;
      patterns[62754] = 29'b1_111010100100_010_1_110101001001;
      patterns[62755] = 29'b1_111010100100_011_1_101010010011;
      patterns[62756] = 29'b1_111010100100_100_0_111101010010;
      patterns[62757] = 29'b1_111010100100_101_0_011110101001;
      patterns[62758] = 29'b1_111010100100_110_1_111010100100;
      patterns[62759] = 29'b1_111010100100_111_1_111010100100;
      patterns[62760] = 29'b1_111010100101_000_1_111010100101;
      patterns[62761] = 29'b1_111010100101_001_1_100101111010;
      patterns[62762] = 29'b1_111010100101_010_1_110101001011;
      patterns[62763] = 29'b1_111010100101_011_1_101010010111;
      patterns[62764] = 29'b1_111010100101_100_1_111101010010;
      patterns[62765] = 29'b1_111010100101_101_0_111110101001;
      patterns[62766] = 29'b1_111010100101_110_1_111010100101;
      patterns[62767] = 29'b1_111010100101_111_1_111010100101;
      patterns[62768] = 29'b1_111010100110_000_1_111010100110;
      patterns[62769] = 29'b1_111010100110_001_1_100110111010;
      patterns[62770] = 29'b1_111010100110_010_1_110101001101;
      patterns[62771] = 29'b1_111010100110_011_1_101010011011;
      patterns[62772] = 29'b1_111010100110_100_0_111101010011;
      patterns[62773] = 29'b1_111010100110_101_1_011110101001;
      patterns[62774] = 29'b1_111010100110_110_1_111010100110;
      patterns[62775] = 29'b1_111010100110_111_1_111010100110;
      patterns[62776] = 29'b1_111010100111_000_1_111010100111;
      patterns[62777] = 29'b1_111010100111_001_1_100111111010;
      patterns[62778] = 29'b1_111010100111_010_1_110101001111;
      patterns[62779] = 29'b1_111010100111_011_1_101010011111;
      patterns[62780] = 29'b1_111010100111_100_1_111101010011;
      patterns[62781] = 29'b1_111010100111_101_1_111110101001;
      patterns[62782] = 29'b1_111010100111_110_1_111010100111;
      patterns[62783] = 29'b1_111010100111_111_1_111010100111;
      patterns[62784] = 29'b1_111010101000_000_1_111010101000;
      patterns[62785] = 29'b1_111010101000_001_1_101000111010;
      patterns[62786] = 29'b1_111010101000_010_1_110101010001;
      patterns[62787] = 29'b1_111010101000_011_1_101010100011;
      patterns[62788] = 29'b1_111010101000_100_0_111101010100;
      patterns[62789] = 29'b1_111010101000_101_0_011110101010;
      patterns[62790] = 29'b1_111010101000_110_1_111010101000;
      patterns[62791] = 29'b1_111010101000_111_1_111010101000;
      patterns[62792] = 29'b1_111010101001_000_1_111010101001;
      patterns[62793] = 29'b1_111010101001_001_1_101001111010;
      patterns[62794] = 29'b1_111010101001_010_1_110101010011;
      patterns[62795] = 29'b1_111010101001_011_1_101010100111;
      patterns[62796] = 29'b1_111010101001_100_1_111101010100;
      patterns[62797] = 29'b1_111010101001_101_0_111110101010;
      patterns[62798] = 29'b1_111010101001_110_1_111010101001;
      patterns[62799] = 29'b1_111010101001_111_1_111010101001;
      patterns[62800] = 29'b1_111010101010_000_1_111010101010;
      patterns[62801] = 29'b1_111010101010_001_1_101010111010;
      patterns[62802] = 29'b1_111010101010_010_1_110101010101;
      patterns[62803] = 29'b1_111010101010_011_1_101010101011;
      patterns[62804] = 29'b1_111010101010_100_0_111101010101;
      patterns[62805] = 29'b1_111010101010_101_1_011110101010;
      patterns[62806] = 29'b1_111010101010_110_1_111010101010;
      patterns[62807] = 29'b1_111010101010_111_1_111010101010;
      patterns[62808] = 29'b1_111010101011_000_1_111010101011;
      patterns[62809] = 29'b1_111010101011_001_1_101011111010;
      patterns[62810] = 29'b1_111010101011_010_1_110101010111;
      patterns[62811] = 29'b1_111010101011_011_1_101010101111;
      patterns[62812] = 29'b1_111010101011_100_1_111101010101;
      patterns[62813] = 29'b1_111010101011_101_1_111110101010;
      patterns[62814] = 29'b1_111010101011_110_1_111010101011;
      patterns[62815] = 29'b1_111010101011_111_1_111010101011;
      patterns[62816] = 29'b1_111010101100_000_1_111010101100;
      patterns[62817] = 29'b1_111010101100_001_1_101100111010;
      patterns[62818] = 29'b1_111010101100_010_1_110101011001;
      patterns[62819] = 29'b1_111010101100_011_1_101010110011;
      patterns[62820] = 29'b1_111010101100_100_0_111101010110;
      patterns[62821] = 29'b1_111010101100_101_0_011110101011;
      patterns[62822] = 29'b1_111010101100_110_1_111010101100;
      patterns[62823] = 29'b1_111010101100_111_1_111010101100;
      patterns[62824] = 29'b1_111010101101_000_1_111010101101;
      patterns[62825] = 29'b1_111010101101_001_1_101101111010;
      patterns[62826] = 29'b1_111010101101_010_1_110101011011;
      patterns[62827] = 29'b1_111010101101_011_1_101010110111;
      patterns[62828] = 29'b1_111010101101_100_1_111101010110;
      patterns[62829] = 29'b1_111010101101_101_0_111110101011;
      patterns[62830] = 29'b1_111010101101_110_1_111010101101;
      patterns[62831] = 29'b1_111010101101_111_1_111010101101;
      patterns[62832] = 29'b1_111010101110_000_1_111010101110;
      patterns[62833] = 29'b1_111010101110_001_1_101110111010;
      patterns[62834] = 29'b1_111010101110_010_1_110101011101;
      patterns[62835] = 29'b1_111010101110_011_1_101010111011;
      patterns[62836] = 29'b1_111010101110_100_0_111101010111;
      patterns[62837] = 29'b1_111010101110_101_1_011110101011;
      patterns[62838] = 29'b1_111010101110_110_1_111010101110;
      patterns[62839] = 29'b1_111010101110_111_1_111010101110;
      patterns[62840] = 29'b1_111010101111_000_1_111010101111;
      patterns[62841] = 29'b1_111010101111_001_1_101111111010;
      patterns[62842] = 29'b1_111010101111_010_1_110101011111;
      patterns[62843] = 29'b1_111010101111_011_1_101010111111;
      patterns[62844] = 29'b1_111010101111_100_1_111101010111;
      patterns[62845] = 29'b1_111010101111_101_1_111110101011;
      patterns[62846] = 29'b1_111010101111_110_1_111010101111;
      patterns[62847] = 29'b1_111010101111_111_1_111010101111;
      patterns[62848] = 29'b1_111010110000_000_1_111010110000;
      patterns[62849] = 29'b1_111010110000_001_1_110000111010;
      patterns[62850] = 29'b1_111010110000_010_1_110101100001;
      patterns[62851] = 29'b1_111010110000_011_1_101011000011;
      patterns[62852] = 29'b1_111010110000_100_0_111101011000;
      patterns[62853] = 29'b1_111010110000_101_0_011110101100;
      patterns[62854] = 29'b1_111010110000_110_1_111010110000;
      patterns[62855] = 29'b1_111010110000_111_1_111010110000;
      patterns[62856] = 29'b1_111010110001_000_1_111010110001;
      patterns[62857] = 29'b1_111010110001_001_1_110001111010;
      patterns[62858] = 29'b1_111010110001_010_1_110101100011;
      patterns[62859] = 29'b1_111010110001_011_1_101011000111;
      patterns[62860] = 29'b1_111010110001_100_1_111101011000;
      patterns[62861] = 29'b1_111010110001_101_0_111110101100;
      patterns[62862] = 29'b1_111010110001_110_1_111010110001;
      patterns[62863] = 29'b1_111010110001_111_1_111010110001;
      patterns[62864] = 29'b1_111010110010_000_1_111010110010;
      patterns[62865] = 29'b1_111010110010_001_1_110010111010;
      patterns[62866] = 29'b1_111010110010_010_1_110101100101;
      patterns[62867] = 29'b1_111010110010_011_1_101011001011;
      patterns[62868] = 29'b1_111010110010_100_0_111101011001;
      patterns[62869] = 29'b1_111010110010_101_1_011110101100;
      patterns[62870] = 29'b1_111010110010_110_1_111010110010;
      patterns[62871] = 29'b1_111010110010_111_1_111010110010;
      patterns[62872] = 29'b1_111010110011_000_1_111010110011;
      patterns[62873] = 29'b1_111010110011_001_1_110011111010;
      patterns[62874] = 29'b1_111010110011_010_1_110101100111;
      patterns[62875] = 29'b1_111010110011_011_1_101011001111;
      patterns[62876] = 29'b1_111010110011_100_1_111101011001;
      patterns[62877] = 29'b1_111010110011_101_1_111110101100;
      patterns[62878] = 29'b1_111010110011_110_1_111010110011;
      patterns[62879] = 29'b1_111010110011_111_1_111010110011;
      patterns[62880] = 29'b1_111010110100_000_1_111010110100;
      patterns[62881] = 29'b1_111010110100_001_1_110100111010;
      patterns[62882] = 29'b1_111010110100_010_1_110101101001;
      patterns[62883] = 29'b1_111010110100_011_1_101011010011;
      patterns[62884] = 29'b1_111010110100_100_0_111101011010;
      patterns[62885] = 29'b1_111010110100_101_0_011110101101;
      patterns[62886] = 29'b1_111010110100_110_1_111010110100;
      patterns[62887] = 29'b1_111010110100_111_1_111010110100;
      patterns[62888] = 29'b1_111010110101_000_1_111010110101;
      patterns[62889] = 29'b1_111010110101_001_1_110101111010;
      patterns[62890] = 29'b1_111010110101_010_1_110101101011;
      patterns[62891] = 29'b1_111010110101_011_1_101011010111;
      patterns[62892] = 29'b1_111010110101_100_1_111101011010;
      patterns[62893] = 29'b1_111010110101_101_0_111110101101;
      patterns[62894] = 29'b1_111010110101_110_1_111010110101;
      patterns[62895] = 29'b1_111010110101_111_1_111010110101;
      patterns[62896] = 29'b1_111010110110_000_1_111010110110;
      patterns[62897] = 29'b1_111010110110_001_1_110110111010;
      patterns[62898] = 29'b1_111010110110_010_1_110101101101;
      patterns[62899] = 29'b1_111010110110_011_1_101011011011;
      patterns[62900] = 29'b1_111010110110_100_0_111101011011;
      patterns[62901] = 29'b1_111010110110_101_1_011110101101;
      patterns[62902] = 29'b1_111010110110_110_1_111010110110;
      patterns[62903] = 29'b1_111010110110_111_1_111010110110;
      patterns[62904] = 29'b1_111010110111_000_1_111010110111;
      patterns[62905] = 29'b1_111010110111_001_1_110111111010;
      patterns[62906] = 29'b1_111010110111_010_1_110101101111;
      patterns[62907] = 29'b1_111010110111_011_1_101011011111;
      patterns[62908] = 29'b1_111010110111_100_1_111101011011;
      patterns[62909] = 29'b1_111010110111_101_1_111110101101;
      patterns[62910] = 29'b1_111010110111_110_1_111010110111;
      patterns[62911] = 29'b1_111010110111_111_1_111010110111;
      patterns[62912] = 29'b1_111010111000_000_1_111010111000;
      patterns[62913] = 29'b1_111010111000_001_1_111000111010;
      patterns[62914] = 29'b1_111010111000_010_1_110101110001;
      patterns[62915] = 29'b1_111010111000_011_1_101011100011;
      patterns[62916] = 29'b1_111010111000_100_0_111101011100;
      patterns[62917] = 29'b1_111010111000_101_0_011110101110;
      patterns[62918] = 29'b1_111010111000_110_1_111010111000;
      patterns[62919] = 29'b1_111010111000_111_1_111010111000;
      patterns[62920] = 29'b1_111010111001_000_1_111010111001;
      patterns[62921] = 29'b1_111010111001_001_1_111001111010;
      patterns[62922] = 29'b1_111010111001_010_1_110101110011;
      patterns[62923] = 29'b1_111010111001_011_1_101011100111;
      patterns[62924] = 29'b1_111010111001_100_1_111101011100;
      patterns[62925] = 29'b1_111010111001_101_0_111110101110;
      patterns[62926] = 29'b1_111010111001_110_1_111010111001;
      patterns[62927] = 29'b1_111010111001_111_1_111010111001;
      patterns[62928] = 29'b1_111010111010_000_1_111010111010;
      patterns[62929] = 29'b1_111010111010_001_1_111010111010;
      patterns[62930] = 29'b1_111010111010_010_1_110101110101;
      patterns[62931] = 29'b1_111010111010_011_1_101011101011;
      patterns[62932] = 29'b1_111010111010_100_0_111101011101;
      patterns[62933] = 29'b1_111010111010_101_1_011110101110;
      patterns[62934] = 29'b1_111010111010_110_1_111010111010;
      patterns[62935] = 29'b1_111010111010_111_1_111010111010;
      patterns[62936] = 29'b1_111010111011_000_1_111010111011;
      patterns[62937] = 29'b1_111010111011_001_1_111011111010;
      patterns[62938] = 29'b1_111010111011_010_1_110101110111;
      patterns[62939] = 29'b1_111010111011_011_1_101011101111;
      patterns[62940] = 29'b1_111010111011_100_1_111101011101;
      patterns[62941] = 29'b1_111010111011_101_1_111110101110;
      patterns[62942] = 29'b1_111010111011_110_1_111010111011;
      patterns[62943] = 29'b1_111010111011_111_1_111010111011;
      patterns[62944] = 29'b1_111010111100_000_1_111010111100;
      patterns[62945] = 29'b1_111010111100_001_1_111100111010;
      patterns[62946] = 29'b1_111010111100_010_1_110101111001;
      patterns[62947] = 29'b1_111010111100_011_1_101011110011;
      patterns[62948] = 29'b1_111010111100_100_0_111101011110;
      patterns[62949] = 29'b1_111010111100_101_0_011110101111;
      patterns[62950] = 29'b1_111010111100_110_1_111010111100;
      patterns[62951] = 29'b1_111010111100_111_1_111010111100;
      patterns[62952] = 29'b1_111010111101_000_1_111010111101;
      patterns[62953] = 29'b1_111010111101_001_1_111101111010;
      patterns[62954] = 29'b1_111010111101_010_1_110101111011;
      patterns[62955] = 29'b1_111010111101_011_1_101011110111;
      patterns[62956] = 29'b1_111010111101_100_1_111101011110;
      patterns[62957] = 29'b1_111010111101_101_0_111110101111;
      patterns[62958] = 29'b1_111010111101_110_1_111010111101;
      patterns[62959] = 29'b1_111010111101_111_1_111010111101;
      patterns[62960] = 29'b1_111010111110_000_1_111010111110;
      patterns[62961] = 29'b1_111010111110_001_1_111110111010;
      patterns[62962] = 29'b1_111010111110_010_1_110101111101;
      patterns[62963] = 29'b1_111010111110_011_1_101011111011;
      patterns[62964] = 29'b1_111010111110_100_0_111101011111;
      patterns[62965] = 29'b1_111010111110_101_1_011110101111;
      patterns[62966] = 29'b1_111010111110_110_1_111010111110;
      patterns[62967] = 29'b1_111010111110_111_1_111010111110;
      patterns[62968] = 29'b1_111010111111_000_1_111010111111;
      patterns[62969] = 29'b1_111010111111_001_1_111111111010;
      patterns[62970] = 29'b1_111010111111_010_1_110101111111;
      patterns[62971] = 29'b1_111010111111_011_1_101011111111;
      patterns[62972] = 29'b1_111010111111_100_1_111101011111;
      patterns[62973] = 29'b1_111010111111_101_1_111110101111;
      patterns[62974] = 29'b1_111010111111_110_1_111010111111;
      patterns[62975] = 29'b1_111010111111_111_1_111010111111;
      patterns[62976] = 29'b1_111011000000_000_1_111011000000;
      patterns[62977] = 29'b1_111011000000_001_1_000000111011;
      patterns[62978] = 29'b1_111011000000_010_1_110110000001;
      patterns[62979] = 29'b1_111011000000_011_1_101100000011;
      patterns[62980] = 29'b1_111011000000_100_0_111101100000;
      patterns[62981] = 29'b1_111011000000_101_0_011110110000;
      patterns[62982] = 29'b1_111011000000_110_1_111011000000;
      patterns[62983] = 29'b1_111011000000_111_1_111011000000;
      patterns[62984] = 29'b1_111011000001_000_1_111011000001;
      patterns[62985] = 29'b1_111011000001_001_1_000001111011;
      patterns[62986] = 29'b1_111011000001_010_1_110110000011;
      patterns[62987] = 29'b1_111011000001_011_1_101100000111;
      patterns[62988] = 29'b1_111011000001_100_1_111101100000;
      patterns[62989] = 29'b1_111011000001_101_0_111110110000;
      patterns[62990] = 29'b1_111011000001_110_1_111011000001;
      patterns[62991] = 29'b1_111011000001_111_1_111011000001;
      patterns[62992] = 29'b1_111011000010_000_1_111011000010;
      patterns[62993] = 29'b1_111011000010_001_1_000010111011;
      patterns[62994] = 29'b1_111011000010_010_1_110110000101;
      patterns[62995] = 29'b1_111011000010_011_1_101100001011;
      patterns[62996] = 29'b1_111011000010_100_0_111101100001;
      patterns[62997] = 29'b1_111011000010_101_1_011110110000;
      patterns[62998] = 29'b1_111011000010_110_1_111011000010;
      patterns[62999] = 29'b1_111011000010_111_1_111011000010;
      patterns[63000] = 29'b1_111011000011_000_1_111011000011;
      patterns[63001] = 29'b1_111011000011_001_1_000011111011;
      patterns[63002] = 29'b1_111011000011_010_1_110110000111;
      patterns[63003] = 29'b1_111011000011_011_1_101100001111;
      patterns[63004] = 29'b1_111011000011_100_1_111101100001;
      patterns[63005] = 29'b1_111011000011_101_1_111110110000;
      patterns[63006] = 29'b1_111011000011_110_1_111011000011;
      patterns[63007] = 29'b1_111011000011_111_1_111011000011;
      patterns[63008] = 29'b1_111011000100_000_1_111011000100;
      patterns[63009] = 29'b1_111011000100_001_1_000100111011;
      patterns[63010] = 29'b1_111011000100_010_1_110110001001;
      patterns[63011] = 29'b1_111011000100_011_1_101100010011;
      patterns[63012] = 29'b1_111011000100_100_0_111101100010;
      patterns[63013] = 29'b1_111011000100_101_0_011110110001;
      patterns[63014] = 29'b1_111011000100_110_1_111011000100;
      patterns[63015] = 29'b1_111011000100_111_1_111011000100;
      patterns[63016] = 29'b1_111011000101_000_1_111011000101;
      patterns[63017] = 29'b1_111011000101_001_1_000101111011;
      patterns[63018] = 29'b1_111011000101_010_1_110110001011;
      patterns[63019] = 29'b1_111011000101_011_1_101100010111;
      patterns[63020] = 29'b1_111011000101_100_1_111101100010;
      patterns[63021] = 29'b1_111011000101_101_0_111110110001;
      patterns[63022] = 29'b1_111011000101_110_1_111011000101;
      patterns[63023] = 29'b1_111011000101_111_1_111011000101;
      patterns[63024] = 29'b1_111011000110_000_1_111011000110;
      patterns[63025] = 29'b1_111011000110_001_1_000110111011;
      patterns[63026] = 29'b1_111011000110_010_1_110110001101;
      patterns[63027] = 29'b1_111011000110_011_1_101100011011;
      patterns[63028] = 29'b1_111011000110_100_0_111101100011;
      patterns[63029] = 29'b1_111011000110_101_1_011110110001;
      patterns[63030] = 29'b1_111011000110_110_1_111011000110;
      patterns[63031] = 29'b1_111011000110_111_1_111011000110;
      patterns[63032] = 29'b1_111011000111_000_1_111011000111;
      patterns[63033] = 29'b1_111011000111_001_1_000111111011;
      patterns[63034] = 29'b1_111011000111_010_1_110110001111;
      patterns[63035] = 29'b1_111011000111_011_1_101100011111;
      patterns[63036] = 29'b1_111011000111_100_1_111101100011;
      patterns[63037] = 29'b1_111011000111_101_1_111110110001;
      patterns[63038] = 29'b1_111011000111_110_1_111011000111;
      patterns[63039] = 29'b1_111011000111_111_1_111011000111;
      patterns[63040] = 29'b1_111011001000_000_1_111011001000;
      patterns[63041] = 29'b1_111011001000_001_1_001000111011;
      patterns[63042] = 29'b1_111011001000_010_1_110110010001;
      patterns[63043] = 29'b1_111011001000_011_1_101100100011;
      patterns[63044] = 29'b1_111011001000_100_0_111101100100;
      patterns[63045] = 29'b1_111011001000_101_0_011110110010;
      patterns[63046] = 29'b1_111011001000_110_1_111011001000;
      patterns[63047] = 29'b1_111011001000_111_1_111011001000;
      patterns[63048] = 29'b1_111011001001_000_1_111011001001;
      patterns[63049] = 29'b1_111011001001_001_1_001001111011;
      patterns[63050] = 29'b1_111011001001_010_1_110110010011;
      patterns[63051] = 29'b1_111011001001_011_1_101100100111;
      patterns[63052] = 29'b1_111011001001_100_1_111101100100;
      patterns[63053] = 29'b1_111011001001_101_0_111110110010;
      patterns[63054] = 29'b1_111011001001_110_1_111011001001;
      patterns[63055] = 29'b1_111011001001_111_1_111011001001;
      patterns[63056] = 29'b1_111011001010_000_1_111011001010;
      patterns[63057] = 29'b1_111011001010_001_1_001010111011;
      patterns[63058] = 29'b1_111011001010_010_1_110110010101;
      patterns[63059] = 29'b1_111011001010_011_1_101100101011;
      patterns[63060] = 29'b1_111011001010_100_0_111101100101;
      patterns[63061] = 29'b1_111011001010_101_1_011110110010;
      patterns[63062] = 29'b1_111011001010_110_1_111011001010;
      patterns[63063] = 29'b1_111011001010_111_1_111011001010;
      patterns[63064] = 29'b1_111011001011_000_1_111011001011;
      patterns[63065] = 29'b1_111011001011_001_1_001011111011;
      patterns[63066] = 29'b1_111011001011_010_1_110110010111;
      patterns[63067] = 29'b1_111011001011_011_1_101100101111;
      patterns[63068] = 29'b1_111011001011_100_1_111101100101;
      patterns[63069] = 29'b1_111011001011_101_1_111110110010;
      patterns[63070] = 29'b1_111011001011_110_1_111011001011;
      patterns[63071] = 29'b1_111011001011_111_1_111011001011;
      patterns[63072] = 29'b1_111011001100_000_1_111011001100;
      patterns[63073] = 29'b1_111011001100_001_1_001100111011;
      patterns[63074] = 29'b1_111011001100_010_1_110110011001;
      patterns[63075] = 29'b1_111011001100_011_1_101100110011;
      patterns[63076] = 29'b1_111011001100_100_0_111101100110;
      patterns[63077] = 29'b1_111011001100_101_0_011110110011;
      patterns[63078] = 29'b1_111011001100_110_1_111011001100;
      patterns[63079] = 29'b1_111011001100_111_1_111011001100;
      patterns[63080] = 29'b1_111011001101_000_1_111011001101;
      patterns[63081] = 29'b1_111011001101_001_1_001101111011;
      patterns[63082] = 29'b1_111011001101_010_1_110110011011;
      patterns[63083] = 29'b1_111011001101_011_1_101100110111;
      patterns[63084] = 29'b1_111011001101_100_1_111101100110;
      patterns[63085] = 29'b1_111011001101_101_0_111110110011;
      patterns[63086] = 29'b1_111011001101_110_1_111011001101;
      patterns[63087] = 29'b1_111011001101_111_1_111011001101;
      patterns[63088] = 29'b1_111011001110_000_1_111011001110;
      patterns[63089] = 29'b1_111011001110_001_1_001110111011;
      patterns[63090] = 29'b1_111011001110_010_1_110110011101;
      patterns[63091] = 29'b1_111011001110_011_1_101100111011;
      patterns[63092] = 29'b1_111011001110_100_0_111101100111;
      patterns[63093] = 29'b1_111011001110_101_1_011110110011;
      patterns[63094] = 29'b1_111011001110_110_1_111011001110;
      patterns[63095] = 29'b1_111011001110_111_1_111011001110;
      patterns[63096] = 29'b1_111011001111_000_1_111011001111;
      patterns[63097] = 29'b1_111011001111_001_1_001111111011;
      patterns[63098] = 29'b1_111011001111_010_1_110110011111;
      patterns[63099] = 29'b1_111011001111_011_1_101100111111;
      patterns[63100] = 29'b1_111011001111_100_1_111101100111;
      patterns[63101] = 29'b1_111011001111_101_1_111110110011;
      patterns[63102] = 29'b1_111011001111_110_1_111011001111;
      patterns[63103] = 29'b1_111011001111_111_1_111011001111;
      patterns[63104] = 29'b1_111011010000_000_1_111011010000;
      patterns[63105] = 29'b1_111011010000_001_1_010000111011;
      patterns[63106] = 29'b1_111011010000_010_1_110110100001;
      patterns[63107] = 29'b1_111011010000_011_1_101101000011;
      patterns[63108] = 29'b1_111011010000_100_0_111101101000;
      patterns[63109] = 29'b1_111011010000_101_0_011110110100;
      patterns[63110] = 29'b1_111011010000_110_1_111011010000;
      patterns[63111] = 29'b1_111011010000_111_1_111011010000;
      patterns[63112] = 29'b1_111011010001_000_1_111011010001;
      patterns[63113] = 29'b1_111011010001_001_1_010001111011;
      patterns[63114] = 29'b1_111011010001_010_1_110110100011;
      patterns[63115] = 29'b1_111011010001_011_1_101101000111;
      patterns[63116] = 29'b1_111011010001_100_1_111101101000;
      patterns[63117] = 29'b1_111011010001_101_0_111110110100;
      patterns[63118] = 29'b1_111011010001_110_1_111011010001;
      patterns[63119] = 29'b1_111011010001_111_1_111011010001;
      patterns[63120] = 29'b1_111011010010_000_1_111011010010;
      patterns[63121] = 29'b1_111011010010_001_1_010010111011;
      patterns[63122] = 29'b1_111011010010_010_1_110110100101;
      patterns[63123] = 29'b1_111011010010_011_1_101101001011;
      patterns[63124] = 29'b1_111011010010_100_0_111101101001;
      patterns[63125] = 29'b1_111011010010_101_1_011110110100;
      patterns[63126] = 29'b1_111011010010_110_1_111011010010;
      patterns[63127] = 29'b1_111011010010_111_1_111011010010;
      patterns[63128] = 29'b1_111011010011_000_1_111011010011;
      patterns[63129] = 29'b1_111011010011_001_1_010011111011;
      patterns[63130] = 29'b1_111011010011_010_1_110110100111;
      patterns[63131] = 29'b1_111011010011_011_1_101101001111;
      patterns[63132] = 29'b1_111011010011_100_1_111101101001;
      patterns[63133] = 29'b1_111011010011_101_1_111110110100;
      patterns[63134] = 29'b1_111011010011_110_1_111011010011;
      patterns[63135] = 29'b1_111011010011_111_1_111011010011;
      patterns[63136] = 29'b1_111011010100_000_1_111011010100;
      patterns[63137] = 29'b1_111011010100_001_1_010100111011;
      patterns[63138] = 29'b1_111011010100_010_1_110110101001;
      patterns[63139] = 29'b1_111011010100_011_1_101101010011;
      patterns[63140] = 29'b1_111011010100_100_0_111101101010;
      patterns[63141] = 29'b1_111011010100_101_0_011110110101;
      patterns[63142] = 29'b1_111011010100_110_1_111011010100;
      patterns[63143] = 29'b1_111011010100_111_1_111011010100;
      patterns[63144] = 29'b1_111011010101_000_1_111011010101;
      patterns[63145] = 29'b1_111011010101_001_1_010101111011;
      patterns[63146] = 29'b1_111011010101_010_1_110110101011;
      patterns[63147] = 29'b1_111011010101_011_1_101101010111;
      patterns[63148] = 29'b1_111011010101_100_1_111101101010;
      patterns[63149] = 29'b1_111011010101_101_0_111110110101;
      patterns[63150] = 29'b1_111011010101_110_1_111011010101;
      patterns[63151] = 29'b1_111011010101_111_1_111011010101;
      patterns[63152] = 29'b1_111011010110_000_1_111011010110;
      patterns[63153] = 29'b1_111011010110_001_1_010110111011;
      patterns[63154] = 29'b1_111011010110_010_1_110110101101;
      patterns[63155] = 29'b1_111011010110_011_1_101101011011;
      patterns[63156] = 29'b1_111011010110_100_0_111101101011;
      patterns[63157] = 29'b1_111011010110_101_1_011110110101;
      patterns[63158] = 29'b1_111011010110_110_1_111011010110;
      patterns[63159] = 29'b1_111011010110_111_1_111011010110;
      patterns[63160] = 29'b1_111011010111_000_1_111011010111;
      patterns[63161] = 29'b1_111011010111_001_1_010111111011;
      patterns[63162] = 29'b1_111011010111_010_1_110110101111;
      patterns[63163] = 29'b1_111011010111_011_1_101101011111;
      patterns[63164] = 29'b1_111011010111_100_1_111101101011;
      patterns[63165] = 29'b1_111011010111_101_1_111110110101;
      patterns[63166] = 29'b1_111011010111_110_1_111011010111;
      patterns[63167] = 29'b1_111011010111_111_1_111011010111;
      patterns[63168] = 29'b1_111011011000_000_1_111011011000;
      patterns[63169] = 29'b1_111011011000_001_1_011000111011;
      patterns[63170] = 29'b1_111011011000_010_1_110110110001;
      patterns[63171] = 29'b1_111011011000_011_1_101101100011;
      patterns[63172] = 29'b1_111011011000_100_0_111101101100;
      patterns[63173] = 29'b1_111011011000_101_0_011110110110;
      patterns[63174] = 29'b1_111011011000_110_1_111011011000;
      patterns[63175] = 29'b1_111011011000_111_1_111011011000;
      patterns[63176] = 29'b1_111011011001_000_1_111011011001;
      patterns[63177] = 29'b1_111011011001_001_1_011001111011;
      patterns[63178] = 29'b1_111011011001_010_1_110110110011;
      patterns[63179] = 29'b1_111011011001_011_1_101101100111;
      patterns[63180] = 29'b1_111011011001_100_1_111101101100;
      patterns[63181] = 29'b1_111011011001_101_0_111110110110;
      patterns[63182] = 29'b1_111011011001_110_1_111011011001;
      patterns[63183] = 29'b1_111011011001_111_1_111011011001;
      patterns[63184] = 29'b1_111011011010_000_1_111011011010;
      patterns[63185] = 29'b1_111011011010_001_1_011010111011;
      patterns[63186] = 29'b1_111011011010_010_1_110110110101;
      patterns[63187] = 29'b1_111011011010_011_1_101101101011;
      patterns[63188] = 29'b1_111011011010_100_0_111101101101;
      patterns[63189] = 29'b1_111011011010_101_1_011110110110;
      patterns[63190] = 29'b1_111011011010_110_1_111011011010;
      patterns[63191] = 29'b1_111011011010_111_1_111011011010;
      patterns[63192] = 29'b1_111011011011_000_1_111011011011;
      patterns[63193] = 29'b1_111011011011_001_1_011011111011;
      patterns[63194] = 29'b1_111011011011_010_1_110110110111;
      patterns[63195] = 29'b1_111011011011_011_1_101101101111;
      patterns[63196] = 29'b1_111011011011_100_1_111101101101;
      patterns[63197] = 29'b1_111011011011_101_1_111110110110;
      patterns[63198] = 29'b1_111011011011_110_1_111011011011;
      patterns[63199] = 29'b1_111011011011_111_1_111011011011;
      patterns[63200] = 29'b1_111011011100_000_1_111011011100;
      patterns[63201] = 29'b1_111011011100_001_1_011100111011;
      patterns[63202] = 29'b1_111011011100_010_1_110110111001;
      patterns[63203] = 29'b1_111011011100_011_1_101101110011;
      patterns[63204] = 29'b1_111011011100_100_0_111101101110;
      patterns[63205] = 29'b1_111011011100_101_0_011110110111;
      patterns[63206] = 29'b1_111011011100_110_1_111011011100;
      patterns[63207] = 29'b1_111011011100_111_1_111011011100;
      patterns[63208] = 29'b1_111011011101_000_1_111011011101;
      patterns[63209] = 29'b1_111011011101_001_1_011101111011;
      patterns[63210] = 29'b1_111011011101_010_1_110110111011;
      patterns[63211] = 29'b1_111011011101_011_1_101101110111;
      patterns[63212] = 29'b1_111011011101_100_1_111101101110;
      patterns[63213] = 29'b1_111011011101_101_0_111110110111;
      patterns[63214] = 29'b1_111011011101_110_1_111011011101;
      patterns[63215] = 29'b1_111011011101_111_1_111011011101;
      patterns[63216] = 29'b1_111011011110_000_1_111011011110;
      patterns[63217] = 29'b1_111011011110_001_1_011110111011;
      patterns[63218] = 29'b1_111011011110_010_1_110110111101;
      patterns[63219] = 29'b1_111011011110_011_1_101101111011;
      patterns[63220] = 29'b1_111011011110_100_0_111101101111;
      patterns[63221] = 29'b1_111011011110_101_1_011110110111;
      patterns[63222] = 29'b1_111011011110_110_1_111011011110;
      patterns[63223] = 29'b1_111011011110_111_1_111011011110;
      patterns[63224] = 29'b1_111011011111_000_1_111011011111;
      patterns[63225] = 29'b1_111011011111_001_1_011111111011;
      patterns[63226] = 29'b1_111011011111_010_1_110110111111;
      patterns[63227] = 29'b1_111011011111_011_1_101101111111;
      patterns[63228] = 29'b1_111011011111_100_1_111101101111;
      patterns[63229] = 29'b1_111011011111_101_1_111110110111;
      patterns[63230] = 29'b1_111011011111_110_1_111011011111;
      patterns[63231] = 29'b1_111011011111_111_1_111011011111;
      patterns[63232] = 29'b1_111011100000_000_1_111011100000;
      patterns[63233] = 29'b1_111011100000_001_1_100000111011;
      patterns[63234] = 29'b1_111011100000_010_1_110111000001;
      patterns[63235] = 29'b1_111011100000_011_1_101110000011;
      patterns[63236] = 29'b1_111011100000_100_0_111101110000;
      patterns[63237] = 29'b1_111011100000_101_0_011110111000;
      patterns[63238] = 29'b1_111011100000_110_1_111011100000;
      patterns[63239] = 29'b1_111011100000_111_1_111011100000;
      patterns[63240] = 29'b1_111011100001_000_1_111011100001;
      patterns[63241] = 29'b1_111011100001_001_1_100001111011;
      patterns[63242] = 29'b1_111011100001_010_1_110111000011;
      patterns[63243] = 29'b1_111011100001_011_1_101110000111;
      patterns[63244] = 29'b1_111011100001_100_1_111101110000;
      patterns[63245] = 29'b1_111011100001_101_0_111110111000;
      patterns[63246] = 29'b1_111011100001_110_1_111011100001;
      patterns[63247] = 29'b1_111011100001_111_1_111011100001;
      patterns[63248] = 29'b1_111011100010_000_1_111011100010;
      patterns[63249] = 29'b1_111011100010_001_1_100010111011;
      patterns[63250] = 29'b1_111011100010_010_1_110111000101;
      patterns[63251] = 29'b1_111011100010_011_1_101110001011;
      patterns[63252] = 29'b1_111011100010_100_0_111101110001;
      patterns[63253] = 29'b1_111011100010_101_1_011110111000;
      patterns[63254] = 29'b1_111011100010_110_1_111011100010;
      patterns[63255] = 29'b1_111011100010_111_1_111011100010;
      patterns[63256] = 29'b1_111011100011_000_1_111011100011;
      patterns[63257] = 29'b1_111011100011_001_1_100011111011;
      patterns[63258] = 29'b1_111011100011_010_1_110111000111;
      patterns[63259] = 29'b1_111011100011_011_1_101110001111;
      patterns[63260] = 29'b1_111011100011_100_1_111101110001;
      patterns[63261] = 29'b1_111011100011_101_1_111110111000;
      patterns[63262] = 29'b1_111011100011_110_1_111011100011;
      patterns[63263] = 29'b1_111011100011_111_1_111011100011;
      patterns[63264] = 29'b1_111011100100_000_1_111011100100;
      patterns[63265] = 29'b1_111011100100_001_1_100100111011;
      patterns[63266] = 29'b1_111011100100_010_1_110111001001;
      patterns[63267] = 29'b1_111011100100_011_1_101110010011;
      patterns[63268] = 29'b1_111011100100_100_0_111101110010;
      patterns[63269] = 29'b1_111011100100_101_0_011110111001;
      patterns[63270] = 29'b1_111011100100_110_1_111011100100;
      patterns[63271] = 29'b1_111011100100_111_1_111011100100;
      patterns[63272] = 29'b1_111011100101_000_1_111011100101;
      patterns[63273] = 29'b1_111011100101_001_1_100101111011;
      patterns[63274] = 29'b1_111011100101_010_1_110111001011;
      patterns[63275] = 29'b1_111011100101_011_1_101110010111;
      patterns[63276] = 29'b1_111011100101_100_1_111101110010;
      patterns[63277] = 29'b1_111011100101_101_0_111110111001;
      patterns[63278] = 29'b1_111011100101_110_1_111011100101;
      patterns[63279] = 29'b1_111011100101_111_1_111011100101;
      patterns[63280] = 29'b1_111011100110_000_1_111011100110;
      patterns[63281] = 29'b1_111011100110_001_1_100110111011;
      patterns[63282] = 29'b1_111011100110_010_1_110111001101;
      patterns[63283] = 29'b1_111011100110_011_1_101110011011;
      patterns[63284] = 29'b1_111011100110_100_0_111101110011;
      patterns[63285] = 29'b1_111011100110_101_1_011110111001;
      patterns[63286] = 29'b1_111011100110_110_1_111011100110;
      patterns[63287] = 29'b1_111011100110_111_1_111011100110;
      patterns[63288] = 29'b1_111011100111_000_1_111011100111;
      patterns[63289] = 29'b1_111011100111_001_1_100111111011;
      patterns[63290] = 29'b1_111011100111_010_1_110111001111;
      patterns[63291] = 29'b1_111011100111_011_1_101110011111;
      patterns[63292] = 29'b1_111011100111_100_1_111101110011;
      patterns[63293] = 29'b1_111011100111_101_1_111110111001;
      patterns[63294] = 29'b1_111011100111_110_1_111011100111;
      patterns[63295] = 29'b1_111011100111_111_1_111011100111;
      patterns[63296] = 29'b1_111011101000_000_1_111011101000;
      patterns[63297] = 29'b1_111011101000_001_1_101000111011;
      patterns[63298] = 29'b1_111011101000_010_1_110111010001;
      patterns[63299] = 29'b1_111011101000_011_1_101110100011;
      patterns[63300] = 29'b1_111011101000_100_0_111101110100;
      patterns[63301] = 29'b1_111011101000_101_0_011110111010;
      patterns[63302] = 29'b1_111011101000_110_1_111011101000;
      patterns[63303] = 29'b1_111011101000_111_1_111011101000;
      patterns[63304] = 29'b1_111011101001_000_1_111011101001;
      patterns[63305] = 29'b1_111011101001_001_1_101001111011;
      patterns[63306] = 29'b1_111011101001_010_1_110111010011;
      patterns[63307] = 29'b1_111011101001_011_1_101110100111;
      patterns[63308] = 29'b1_111011101001_100_1_111101110100;
      patterns[63309] = 29'b1_111011101001_101_0_111110111010;
      patterns[63310] = 29'b1_111011101001_110_1_111011101001;
      patterns[63311] = 29'b1_111011101001_111_1_111011101001;
      patterns[63312] = 29'b1_111011101010_000_1_111011101010;
      patterns[63313] = 29'b1_111011101010_001_1_101010111011;
      patterns[63314] = 29'b1_111011101010_010_1_110111010101;
      patterns[63315] = 29'b1_111011101010_011_1_101110101011;
      patterns[63316] = 29'b1_111011101010_100_0_111101110101;
      patterns[63317] = 29'b1_111011101010_101_1_011110111010;
      patterns[63318] = 29'b1_111011101010_110_1_111011101010;
      patterns[63319] = 29'b1_111011101010_111_1_111011101010;
      patterns[63320] = 29'b1_111011101011_000_1_111011101011;
      patterns[63321] = 29'b1_111011101011_001_1_101011111011;
      patterns[63322] = 29'b1_111011101011_010_1_110111010111;
      patterns[63323] = 29'b1_111011101011_011_1_101110101111;
      patterns[63324] = 29'b1_111011101011_100_1_111101110101;
      patterns[63325] = 29'b1_111011101011_101_1_111110111010;
      patterns[63326] = 29'b1_111011101011_110_1_111011101011;
      patterns[63327] = 29'b1_111011101011_111_1_111011101011;
      patterns[63328] = 29'b1_111011101100_000_1_111011101100;
      patterns[63329] = 29'b1_111011101100_001_1_101100111011;
      patterns[63330] = 29'b1_111011101100_010_1_110111011001;
      patterns[63331] = 29'b1_111011101100_011_1_101110110011;
      patterns[63332] = 29'b1_111011101100_100_0_111101110110;
      patterns[63333] = 29'b1_111011101100_101_0_011110111011;
      patterns[63334] = 29'b1_111011101100_110_1_111011101100;
      patterns[63335] = 29'b1_111011101100_111_1_111011101100;
      patterns[63336] = 29'b1_111011101101_000_1_111011101101;
      patterns[63337] = 29'b1_111011101101_001_1_101101111011;
      patterns[63338] = 29'b1_111011101101_010_1_110111011011;
      patterns[63339] = 29'b1_111011101101_011_1_101110110111;
      patterns[63340] = 29'b1_111011101101_100_1_111101110110;
      patterns[63341] = 29'b1_111011101101_101_0_111110111011;
      patterns[63342] = 29'b1_111011101101_110_1_111011101101;
      patterns[63343] = 29'b1_111011101101_111_1_111011101101;
      patterns[63344] = 29'b1_111011101110_000_1_111011101110;
      patterns[63345] = 29'b1_111011101110_001_1_101110111011;
      patterns[63346] = 29'b1_111011101110_010_1_110111011101;
      patterns[63347] = 29'b1_111011101110_011_1_101110111011;
      patterns[63348] = 29'b1_111011101110_100_0_111101110111;
      patterns[63349] = 29'b1_111011101110_101_1_011110111011;
      patterns[63350] = 29'b1_111011101110_110_1_111011101110;
      patterns[63351] = 29'b1_111011101110_111_1_111011101110;
      patterns[63352] = 29'b1_111011101111_000_1_111011101111;
      patterns[63353] = 29'b1_111011101111_001_1_101111111011;
      patterns[63354] = 29'b1_111011101111_010_1_110111011111;
      patterns[63355] = 29'b1_111011101111_011_1_101110111111;
      patterns[63356] = 29'b1_111011101111_100_1_111101110111;
      patterns[63357] = 29'b1_111011101111_101_1_111110111011;
      patterns[63358] = 29'b1_111011101111_110_1_111011101111;
      patterns[63359] = 29'b1_111011101111_111_1_111011101111;
      patterns[63360] = 29'b1_111011110000_000_1_111011110000;
      patterns[63361] = 29'b1_111011110000_001_1_110000111011;
      patterns[63362] = 29'b1_111011110000_010_1_110111100001;
      patterns[63363] = 29'b1_111011110000_011_1_101111000011;
      patterns[63364] = 29'b1_111011110000_100_0_111101111000;
      patterns[63365] = 29'b1_111011110000_101_0_011110111100;
      patterns[63366] = 29'b1_111011110000_110_1_111011110000;
      patterns[63367] = 29'b1_111011110000_111_1_111011110000;
      patterns[63368] = 29'b1_111011110001_000_1_111011110001;
      patterns[63369] = 29'b1_111011110001_001_1_110001111011;
      patterns[63370] = 29'b1_111011110001_010_1_110111100011;
      patterns[63371] = 29'b1_111011110001_011_1_101111000111;
      patterns[63372] = 29'b1_111011110001_100_1_111101111000;
      patterns[63373] = 29'b1_111011110001_101_0_111110111100;
      patterns[63374] = 29'b1_111011110001_110_1_111011110001;
      patterns[63375] = 29'b1_111011110001_111_1_111011110001;
      patterns[63376] = 29'b1_111011110010_000_1_111011110010;
      patterns[63377] = 29'b1_111011110010_001_1_110010111011;
      patterns[63378] = 29'b1_111011110010_010_1_110111100101;
      patterns[63379] = 29'b1_111011110010_011_1_101111001011;
      patterns[63380] = 29'b1_111011110010_100_0_111101111001;
      patterns[63381] = 29'b1_111011110010_101_1_011110111100;
      patterns[63382] = 29'b1_111011110010_110_1_111011110010;
      patterns[63383] = 29'b1_111011110010_111_1_111011110010;
      patterns[63384] = 29'b1_111011110011_000_1_111011110011;
      patterns[63385] = 29'b1_111011110011_001_1_110011111011;
      patterns[63386] = 29'b1_111011110011_010_1_110111100111;
      patterns[63387] = 29'b1_111011110011_011_1_101111001111;
      patterns[63388] = 29'b1_111011110011_100_1_111101111001;
      patterns[63389] = 29'b1_111011110011_101_1_111110111100;
      patterns[63390] = 29'b1_111011110011_110_1_111011110011;
      patterns[63391] = 29'b1_111011110011_111_1_111011110011;
      patterns[63392] = 29'b1_111011110100_000_1_111011110100;
      patterns[63393] = 29'b1_111011110100_001_1_110100111011;
      patterns[63394] = 29'b1_111011110100_010_1_110111101001;
      patterns[63395] = 29'b1_111011110100_011_1_101111010011;
      patterns[63396] = 29'b1_111011110100_100_0_111101111010;
      patterns[63397] = 29'b1_111011110100_101_0_011110111101;
      patterns[63398] = 29'b1_111011110100_110_1_111011110100;
      patterns[63399] = 29'b1_111011110100_111_1_111011110100;
      patterns[63400] = 29'b1_111011110101_000_1_111011110101;
      patterns[63401] = 29'b1_111011110101_001_1_110101111011;
      patterns[63402] = 29'b1_111011110101_010_1_110111101011;
      patterns[63403] = 29'b1_111011110101_011_1_101111010111;
      patterns[63404] = 29'b1_111011110101_100_1_111101111010;
      patterns[63405] = 29'b1_111011110101_101_0_111110111101;
      patterns[63406] = 29'b1_111011110101_110_1_111011110101;
      patterns[63407] = 29'b1_111011110101_111_1_111011110101;
      patterns[63408] = 29'b1_111011110110_000_1_111011110110;
      patterns[63409] = 29'b1_111011110110_001_1_110110111011;
      patterns[63410] = 29'b1_111011110110_010_1_110111101101;
      patterns[63411] = 29'b1_111011110110_011_1_101111011011;
      patterns[63412] = 29'b1_111011110110_100_0_111101111011;
      patterns[63413] = 29'b1_111011110110_101_1_011110111101;
      patterns[63414] = 29'b1_111011110110_110_1_111011110110;
      patterns[63415] = 29'b1_111011110110_111_1_111011110110;
      patterns[63416] = 29'b1_111011110111_000_1_111011110111;
      patterns[63417] = 29'b1_111011110111_001_1_110111111011;
      patterns[63418] = 29'b1_111011110111_010_1_110111101111;
      patterns[63419] = 29'b1_111011110111_011_1_101111011111;
      patterns[63420] = 29'b1_111011110111_100_1_111101111011;
      patterns[63421] = 29'b1_111011110111_101_1_111110111101;
      patterns[63422] = 29'b1_111011110111_110_1_111011110111;
      patterns[63423] = 29'b1_111011110111_111_1_111011110111;
      patterns[63424] = 29'b1_111011111000_000_1_111011111000;
      patterns[63425] = 29'b1_111011111000_001_1_111000111011;
      patterns[63426] = 29'b1_111011111000_010_1_110111110001;
      patterns[63427] = 29'b1_111011111000_011_1_101111100011;
      patterns[63428] = 29'b1_111011111000_100_0_111101111100;
      patterns[63429] = 29'b1_111011111000_101_0_011110111110;
      patterns[63430] = 29'b1_111011111000_110_1_111011111000;
      patterns[63431] = 29'b1_111011111000_111_1_111011111000;
      patterns[63432] = 29'b1_111011111001_000_1_111011111001;
      patterns[63433] = 29'b1_111011111001_001_1_111001111011;
      patterns[63434] = 29'b1_111011111001_010_1_110111110011;
      patterns[63435] = 29'b1_111011111001_011_1_101111100111;
      patterns[63436] = 29'b1_111011111001_100_1_111101111100;
      patterns[63437] = 29'b1_111011111001_101_0_111110111110;
      patterns[63438] = 29'b1_111011111001_110_1_111011111001;
      patterns[63439] = 29'b1_111011111001_111_1_111011111001;
      patterns[63440] = 29'b1_111011111010_000_1_111011111010;
      patterns[63441] = 29'b1_111011111010_001_1_111010111011;
      patterns[63442] = 29'b1_111011111010_010_1_110111110101;
      patterns[63443] = 29'b1_111011111010_011_1_101111101011;
      patterns[63444] = 29'b1_111011111010_100_0_111101111101;
      patterns[63445] = 29'b1_111011111010_101_1_011110111110;
      patterns[63446] = 29'b1_111011111010_110_1_111011111010;
      patterns[63447] = 29'b1_111011111010_111_1_111011111010;
      patterns[63448] = 29'b1_111011111011_000_1_111011111011;
      patterns[63449] = 29'b1_111011111011_001_1_111011111011;
      patterns[63450] = 29'b1_111011111011_010_1_110111110111;
      patterns[63451] = 29'b1_111011111011_011_1_101111101111;
      patterns[63452] = 29'b1_111011111011_100_1_111101111101;
      patterns[63453] = 29'b1_111011111011_101_1_111110111110;
      patterns[63454] = 29'b1_111011111011_110_1_111011111011;
      patterns[63455] = 29'b1_111011111011_111_1_111011111011;
      patterns[63456] = 29'b1_111011111100_000_1_111011111100;
      patterns[63457] = 29'b1_111011111100_001_1_111100111011;
      patterns[63458] = 29'b1_111011111100_010_1_110111111001;
      patterns[63459] = 29'b1_111011111100_011_1_101111110011;
      patterns[63460] = 29'b1_111011111100_100_0_111101111110;
      patterns[63461] = 29'b1_111011111100_101_0_011110111111;
      patterns[63462] = 29'b1_111011111100_110_1_111011111100;
      patterns[63463] = 29'b1_111011111100_111_1_111011111100;
      patterns[63464] = 29'b1_111011111101_000_1_111011111101;
      patterns[63465] = 29'b1_111011111101_001_1_111101111011;
      patterns[63466] = 29'b1_111011111101_010_1_110111111011;
      patterns[63467] = 29'b1_111011111101_011_1_101111110111;
      patterns[63468] = 29'b1_111011111101_100_1_111101111110;
      patterns[63469] = 29'b1_111011111101_101_0_111110111111;
      patterns[63470] = 29'b1_111011111101_110_1_111011111101;
      patterns[63471] = 29'b1_111011111101_111_1_111011111101;
      patterns[63472] = 29'b1_111011111110_000_1_111011111110;
      patterns[63473] = 29'b1_111011111110_001_1_111110111011;
      patterns[63474] = 29'b1_111011111110_010_1_110111111101;
      patterns[63475] = 29'b1_111011111110_011_1_101111111011;
      patterns[63476] = 29'b1_111011111110_100_0_111101111111;
      patterns[63477] = 29'b1_111011111110_101_1_011110111111;
      patterns[63478] = 29'b1_111011111110_110_1_111011111110;
      patterns[63479] = 29'b1_111011111110_111_1_111011111110;
      patterns[63480] = 29'b1_111011111111_000_1_111011111111;
      patterns[63481] = 29'b1_111011111111_001_1_111111111011;
      patterns[63482] = 29'b1_111011111111_010_1_110111111111;
      patterns[63483] = 29'b1_111011111111_011_1_101111111111;
      patterns[63484] = 29'b1_111011111111_100_1_111101111111;
      patterns[63485] = 29'b1_111011111111_101_1_111110111111;
      patterns[63486] = 29'b1_111011111111_110_1_111011111111;
      patterns[63487] = 29'b1_111011111111_111_1_111011111111;
      patterns[63488] = 29'b1_111100000000_000_1_111100000000;
      patterns[63489] = 29'b1_111100000000_001_1_000000111100;
      patterns[63490] = 29'b1_111100000000_010_1_111000000001;
      patterns[63491] = 29'b1_111100000000_011_1_110000000011;
      patterns[63492] = 29'b1_111100000000_100_0_111110000000;
      patterns[63493] = 29'b1_111100000000_101_0_011111000000;
      patterns[63494] = 29'b1_111100000000_110_1_111100000000;
      patterns[63495] = 29'b1_111100000000_111_1_111100000000;
      patterns[63496] = 29'b1_111100000001_000_1_111100000001;
      patterns[63497] = 29'b1_111100000001_001_1_000001111100;
      patterns[63498] = 29'b1_111100000001_010_1_111000000011;
      patterns[63499] = 29'b1_111100000001_011_1_110000000111;
      patterns[63500] = 29'b1_111100000001_100_1_111110000000;
      patterns[63501] = 29'b1_111100000001_101_0_111111000000;
      patterns[63502] = 29'b1_111100000001_110_1_111100000001;
      patterns[63503] = 29'b1_111100000001_111_1_111100000001;
      patterns[63504] = 29'b1_111100000010_000_1_111100000010;
      patterns[63505] = 29'b1_111100000010_001_1_000010111100;
      patterns[63506] = 29'b1_111100000010_010_1_111000000101;
      patterns[63507] = 29'b1_111100000010_011_1_110000001011;
      patterns[63508] = 29'b1_111100000010_100_0_111110000001;
      patterns[63509] = 29'b1_111100000010_101_1_011111000000;
      patterns[63510] = 29'b1_111100000010_110_1_111100000010;
      patterns[63511] = 29'b1_111100000010_111_1_111100000010;
      patterns[63512] = 29'b1_111100000011_000_1_111100000011;
      patterns[63513] = 29'b1_111100000011_001_1_000011111100;
      patterns[63514] = 29'b1_111100000011_010_1_111000000111;
      patterns[63515] = 29'b1_111100000011_011_1_110000001111;
      patterns[63516] = 29'b1_111100000011_100_1_111110000001;
      patterns[63517] = 29'b1_111100000011_101_1_111111000000;
      patterns[63518] = 29'b1_111100000011_110_1_111100000011;
      patterns[63519] = 29'b1_111100000011_111_1_111100000011;
      patterns[63520] = 29'b1_111100000100_000_1_111100000100;
      patterns[63521] = 29'b1_111100000100_001_1_000100111100;
      patterns[63522] = 29'b1_111100000100_010_1_111000001001;
      patterns[63523] = 29'b1_111100000100_011_1_110000010011;
      patterns[63524] = 29'b1_111100000100_100_0_111110000010;
      patterns[63525] = 29'b1_111100000100_101_0_011111000001;
      patterns[63526] = 29'b1_111100000100_110_1_111100000100;
      patterns[63527] = 29'b1_111100000100_111_1_111100000100;
      patterns[63528] = 29'b1_111100000101_000_1_111100000101;
      patterns[63529] = 29'b1_111100000101_001_1_000101111100;
      patterns[63530] = 29'b1_111100000101_010_1_111000001011;
      patterns[63531] = 29'b1_111100000101_011_1_110000010111;
      patterns[63532] = 29'b1_111100000101_100_1_111110000010;
      patterns[63533] = 29'b1_111100000101_101_0_111111000001;
      patterns[63534] = 29'b1_111100000101_110_1_111100000101;
      patterns[63535] = 29'b1_111100000101_111_1_111100000101;
      patterns[63536] = 29'b1_111100000110_000_1_111100000110;
      patterns[63537] = 29'b1_111100000110_001_1_000110111100;
      patterns[63538] = 29'b1_111100000110_010_1_111000001101;
      patterns[63539] = 29'b1_111100000110_011_1_110000011011;
      patterns[63540] = 29'b1_111100000110_100_0_111110000011;
      patterns[63541] = 29'b1_111100000110_101_1_011111000001;
      patterns[63542] = 29'b1_111100000110_110_1_111100000110;
      patterns[63543] = 29'b1_111100000110_111_1_111100000110;
      patterns[63544] = 29'b1_111100000111_000_1_111100000111;
      patterns[63545] = 29'b1_111100000111_001_1_000111111100;
      patterns[63546] = 29'b1_111100000111_010_1_111000001111;
      patterns[63547] = 29'b1_111100000111_011_1_110000011111;
      patterns[63548] = 29'b1_111100000111_100_1_111110000011;
      patterns[63549] = 29'b1_111100000111_101_1_111111000001;
      patterns[63550] = 29'b1_111100000111_110_1_111100000111;
      patterns[63551] = 29'b1_111100000111_111_1_111100000111;
      patterns[63552] = 29'b1_111100001000_000_1_111100001000;
      patterns[63553] = 29'b1_111100001000_001_1_001000111100;
      patterns[63554] = 29'b1_111100001000_010_1_111000010001;
      patterns[63555] = 29'b1_111100001000_011_1_110000100011;
      patterns[63556] = 29'b1_111100001000_100_0_111110000100;
      patterns[63557] = 29'b1_111100001000_101_0_011111000010;
      patterns[63558] = 29'b1_111100001000_110_1_111100001000;
      patterns[63559] = 29'b1_111100001000_111_1_111100001000;
      patterns[63560] = 29'b1_111100001001_000_1_111100001001;
      patterns[63561] = 29'b1_111100001001_001_1_001001111100;
      patterns[63562] = 29'b1_111100001001_010_1_111000010011;
      patterns[63563] = 29'b1_111100001001_011_1_110000100111;
      patterns[63564] = 29'b1_111100001001_100_1_111110000100;
      patterns[63565] = 29'b1_111100001001_101_0_111111000010;
      patterns[63566] = 29'b1_111100001001_110_1_111100001001;
      patterns[63567] = 29'b1_111100001001_111_1_111100001001;
      patterns[63568] = 29'b1_111100001010_000_1_111100001010;
      patterns[63569] = 29'b1_111100001010_001_1_001010111100;
      patterns[63570] = 29'b1_111100001010_010_1_111000010101;
      patterns[63571] = 29'b1_111100001010_011_1_110000101011;
      patterns[63572] = 29'b1_111100001010_100_0_111110000101;
      patterns[63573] = 29'b1_111100001010_101_1_011111000010;
      patterns[63574] = 29'b1_111100001010_110_1_111100001010;
      patterns[63575] = 29'b1_111100001010_111_1_111100001010;
      patterns[63576] = 29'b1_111100001011_000_1_111100001011;
      patterns[63577] = 29'b1_111100001011_001_1_001011111100;
      patterns[63578] = 29'b1_111100001011_010_1_111000010111;
      patterns[63579] = 29'b1_111100001011_011_1_110000101111;
      patterns[63580] = 29'b1_111100001011_100_1_111110000101;
      patterns[63581] = 29'b1_111100001011_101_1_111111000010;
      patterns[63582] = 29'b1_111100001011_110_1_111100001011;
      patterns[63583] = 29'b1_111100001011_111_1_111100001011;
      patterns[63584] = 29'b1_111100001100_000_1_111100001100;
      patterns[63585] = 29'b1_111100001100_001_1_001100111100;
      patterns[63586] = 29'b1_111100001100_010_1_111000011001;
      patterns[63587] = 29'b1_111100001100_011_1_110000110011;
      patterns[63588] = 29'b1_111100001100_100_0_111110000110;
      patterns[63589] = 29'b1_111100001100_101_0_011111000011;
      patterns[63590] = 29'b1_111100001100_110_1_111100001100;
      patterns[63591] = 29'b1_111100001100_111_1_111100001100;
      patterns[63592] = 29'b1_111100001101_000_1_111100001101;
      patterns[63593] = 29'b1_111100001101_001_1_001101111100;
      patterns[63594] = 29'b1_111100001101_010_1_111000011011;
      patterns[63595] = 29'b1_111100001101_011_1_110000110111;
      patterns[63596] = 29'b1_111100001101_100_1_111110000110;
      patterns[63597] = 29'b1_111100001101_101_0_111111000011;
      patterns[63598] = 29'b1_111100001101_110_1_111100001101;
      patterns[63599] = 29'b1_111100001101_111_1_111100001101;
      patterns[63600] = 29'b1_111100001110_000_1_111100001110;
      patterns[63601] = 29'b1_111100001110_001_1_001110111100;
      patterns[63602] = 29'b1_111100001110_010_1_111000011101;
      patterns[63603] = 29'b1_111100001110_011_1_110000111011;
      patterns[63604] = 29'b1_111100001110_100_0_111110000111;
      patterns[63605] = 29'b1_111100001110_101_1_011111000011;
      patterns[63606] = 29'b1_111100001110_110_1_111100001110;
      patterns[63607] = 29'b1_111100001110_111_1_111100001110;
      patterns[63608] = 29'b1_111100001111_000_1_111100001111;
      patterns[63609] = 29'b1_111100001111_001_1_001111111100;
      patterns[63610] = 29'b1_111100001111_010_1_111000011111;
      patterns[63611] = 29'b1_111100001111_011_1_110000111111;
      patterns[63612] = 29'b1_111100001111_100_1_111110000111;
      patterns[63613] = 29'b1_111100001111_101_1_111111000011;
      patterns[63614] = 29'b1_111100001111_110_1_111100001111;
      patterns[63615] = 29'b1_111100001111_111_1_111100001111;
      patterns[63616] = 29'b1_111100010000_000_1_111100010000;
      patterns[63617] = 29'b1_111100010000_001_1_010000111100;
      patterns[63618] = 29'b1_111100010000_010_1_111000100001;
      patterns[63619] = 29'b1_111100010000_011_1_110001000011;
      patterns[63620] = 29'b1_111100010000_100_0_111110001000;
      patterns[63621] = 29'b1_111100010000_101_0_011111000100;
      patterns[63622] = 29'b1_111100010000_110_1_111100010000;
      patterns[63623] = 29'b1_111100010000_111_1_111100010000;
      patterns[63624] = 29'b1_111100010001_000_1_111100010001;
      patterns[63625] = 29'b1_111100010001_001_1_010001111100;
      patterns[63626] = 29'b1_111100010001_010_1_111000100011;
      patterns[63627] = 29'b1_111100010001_011_1_110001000111;
      patterns[63628] = 29'b1_111100010001_100_1_111110001000;
      patterns[63629] = 29'b1_111100010001_101_0_111111000100;
      patterns[63630] = 29'b1_111100010001_110_1_111100010001;
      patterns[63631] = 29'b1_111100010001_111_1_111100010001;
      patterns[63632] = 29'b1_111100010010_000_1_111100010010;
      patterns[63633] = 29'b1_111100010010_001_1_010010111100;
      patterns[63634] = 29'b1_111100010010_010_1_111000100101;
      patterns[63635] = 29'b1_111100010010_011_1_110001001011;
      patterns[63636] = 29'b1_111100010010_100_0_111110001001;
      patterns[63637] = 29'b1_111100010010_101_1_011111000100;
      patterns[63638] = 29'b1_111100010010_110_1_111100010010;
      patterns[63639] = 29'b1_111100010010_111_1_111100010010;
      patterns[63640] = 29'b1_111100010011_000_1_111100010011;
      patterns[63641] = 29'b1_111100010011_001_1_010011111100;
      patterns[63642] = 29'b1_111100010011_010_1_111000100111;
      patterns[63643] = 29'b1_111100010011_011_1_110001001111;
      patterns[63644] = 29'b1_111100010011_100_1_111110001001;
      patterns[63645] = 29'b1_111100010011_101_1_111111000100;
      patterns[63646] = 29'b1_111100010011_110_1_111100010011;
      patterns[63647] = 29'b1_111100010011_111_1_111100010011;
      patterns[63648] = 29'b1_111100010100_000_1_111100010100;
      patterns[63649] = 29'b1_111100010100_001_1_010100111100;
      patterns[63650] = 29'b1_111100010100_010_1_111000101001;
      patterns[63651] = 29'b1_111100010100_011_1_110001010011;
      patterns[63652] = 29'b1_111100010100_100_0_111110001010;
      patterns[63653] = 29'b1_111100010100_101_0_011111000101;
      patterns[63654] = 29'b1_111100010100_110_1_111100010100;
      patterns[63655] = 29'b1_111100010100_111_1_111100010100;
      patterns[63656] = 29'b1_111100010101_000_1_111100010101;
      patterns[63657] = 29'b1_111100010101_001_1_010101111100;
      patterns[63658] = 29'b1_111100010101_010_1_111000101011;
      patterns[63659] = 29'b1_111100010101_011_1_110001010111;
      patterns[63660] = 29'b1_111100010101_100_1_111110001010;
      patterns[63661] = 29'b1_111100010101_101_0_111111000101;
      patterns[63662] = 29'b1_111100010101_110_1_111100010101;
      patterns[63663] = 29'b1_111100010101_111_1_111100010101;
      patterns[63664] = 29'b1_111100010110_000_1_111100010110;
      patterns[63665] = 29'b1_111100010110_001_1_010110111100;
      patterns[63666] = 29'b1_111100010110_010_1_111000101101;
      patterns[63667] = 29'b1_111100010110_011_1_110001011011;
      patterns[63668] = 29'b1_111100010110_100_0_111110001011;
      patterns[63669] = 29'b1_111100010110_101_1_011111000101;
      patterns[63670] = 29'b1_111100010110_110_1_111100010110;
      patterns[63671] = 29'b1_111100010110_111_1_111100010110;
      patterns[63672] = 29'b1_111100010111_000_1_111100010111;
      patterns[63673] = 29'b1_111100010111_001_1_010111111100;
      patterns[63674] = 29'b1_111100010111_010_1_111000101111;
      patterns[63675] = 29'b1_111100010111_011_1_110001011111;
      patterns[63676] = 29'b1_111100010111_100_1_111110001011;
      patterns[63677] = 29'b1_111100010111_101_1_111111000101;
      patterns[63678] = 29'b1_111100010111_110_1_111100010111;
      patterns[63679] = 29'b1_111100010111_111_1_111100010111;
      patterns[63680] = 29'b1_111100011000_000_1_111100011000;
      patterns[63681] = 29'b1_111100011000_001_1_011000111100;
      patterns[63682] = 29'b1_111100011000_010_1_111000110001;
      patterns[63683] = 29'b1_111100011000_011_1_110001100011;
      patterns[63684] = 29'b1_111100011000_100_0_111110001100;
      patterns[63685] = 29'b1_111100011000_101_0_011111000110;
      patterns[63686] = 29'b1_111100011000_110_1_111100011000;
      patterns[63687] = 29'b1_111100011000_111_1_111100011000;
      patterns[63688] = 29'b1_111100011001_000_1_111100011001;
      patterns[63689] = 29'b1_111100011001_001_1_011001111100;
      patterns[63690] = 29'b1_111100011001_010_1_111000110011;
      patterns[63691] = 29'b1_111100011001_011_1_110001100111;
      patterns[63692] = 29'b1_111100011001_100_1_111110001100;
      patterns[63693] = 29'b1_111100011001_101_0_111111000110;
      patterns[63694] = 29'b1_111100011001_110_1_111100011001;
      patterns[63695] = 29'b1_111100011001_111_1_111100011001;
      patterns[63696] = 29'b1_111100011010_000_1_111100011010;
      patterns[63697] = 29'b1_111100011010_001_1_011010111100;
      patterns[63698] = 29'b1_111100011010_010_1_111000110101;
      patterns[63699] = 29'b1_111100011010_011_1_110001101011;
      patterns[63700] = 29'b1_111100011010_100_0_111110001101;
      patterns[63701] = 29'b1_111100011010_101_1_011111000110;
      patterns[63702] = 29'b1_111100011010_110_1_111100011010;
      patterns[63703] = 29'b1_111100011010_111_1_111100011010;
      patterns[63704] = 29'b1_111100011011_000_1_111100011011;
      patterns[63705] = 29'b1_111100011011_001_1_011011111100;
      patterns[63706] = 29'b1_111100011011_010_1_111000110111;
      patterns[63707] = 29'b1_111100011011_011_1_110001101111;
      patterns[63708] = 29'b1_111100011011_100_1_111110001101;
      patterns[63709] = 29'b1_111100011011_101_1_111111000110;
      patterns[63710] = 29'b1_111100011011_110_1_111100011011;
      patterns[63711] = 29'b1_111100011011_111_1_111100011011;
      patterns[63712] = 29'b1_111100011100_000_1_111100011100;
      patterns[63713] = 29'b1_111100011100_001_1_011100111100;
      patterns[63714] = 29'b1_111100011100_010_1_111000111001;
      patterns[63715] = 29'b1_111100011100_011_1_110001110011;
      patterns[63716] = 29'b1_111100011100_100_0_111110001110;
      patterns[63717] = 29'b1_111100011100_101_0_011111000111;
      patterns[63718] = 29'b1_111100011100_110_1_111100011100;
      patterns[63719] = 29'b1_111100011100_111_1_111100011100;
      patterns[63720] = 29'b1_111100011101_000_1_111100011101;
      patterns[63721] = 29'b1_111100011101_001_1_011101111100;
      patterns[63722] = 29'b1_111100011101_010_1_111000111011;
      patterns[63723] = 29'b1_111100011101_011_1_110001110111;
      patterns[63724] = 29'b1_111100011101_100_1_111110001110;
      patterns[63725] = 29'b1_111100011101_101_0_111111000111;
      patterns[63726] = 29'b1_111100011101_110_1_111100011101;
      patterns[63727] = 29'b1_111100011101_111_1_111100011101;
      patterns[63728] = 29'b1_111100011110_000_1_111100011110;
      patterns[63729] = 29'b1_111100011110_001_1_011110111100;
      patterns[63730] = 29'b1_111100011110_010_1_111000111101;
      patterns[63731] = 29'b1_111100011110_011_1_110001111011;
      patterns[63732] = 29'b1_111100011110_100_0_111110001111;
      patterns[63733] = 29'b1_111100011110_101_1_011111000111;
      patterns[63734] = 29'b1_111100011110_110_1_111100011110;
      patterns[63735] = 29'b1_111100011110_111_1_111100011110;
      patterns[63736] = 29'b1_111100011111_000_1_111100011111;
      patterns[63737] = 29'b1_111100011111_001_1_011111111100;
      patterns[63738] = 29'b1_111100011111_010_1_111000111111;
      patterns[63739] = 29'b1_111100011111_011_1_110001111111;
      patterns[63740] = 29'b1_111100011111_100_1_111110001111;
      patterns[63741] = 29'b1_111100011111_101_1_111111000111;
      patterns[63742] = 29'b1_111100011111_110_1_111100011111;
      patterns[63743] = 29'b1_111100011111_111_1_111100011111;
      patterns[63744] = 29'b1_111100100000_000_1_111100100000;
      patterns[63745] = 29'b1_111100100000_001_1_100000111100;
      patterns[63746] = 29'b1_111100100000_010_1_111001000001;
      patterns[63747] = 29'b1_111100100000_011_1_110010000011;
      patterns[63748] = 29'b1_111100100000_100_0_111110010000;
      patterns[63749] = 29'b1_111100100000_101_0_011111001000;
      patterns[63750] = 29'b1_111100100000_110_1_111100100000;
      patterns[63751] = 29'b1_111100100000_111_1_111100100000;
      patterns[63752] = 29'b1_111100100001_000_1_111100100001;
      patterns[63753] = 29'b1_111100100001_001_1_100001111100;
      patterns[63754] = 29'b1_111100100001_010_1_111001000011;
      patterns[63755] = 29'b1_111100100001_011_1_110010000111;
      patterns[63756] = 29'b1_111100100001_100_1_111110010000;
      patterns[63757] = 29'b1_111100100001_101_0_111111001000;
      patterns[63758] = 29'b1_111100100001_110_1_111100100001;
      patterns[63759] = 29'b1_111100100001_111_1_111100100001;
      patterns[63760] = 29'b1_111100100010_000_1_111100100010;
      patterns[63761] = 29'b1_111100100010_001_1_100010111100;
      patterns[63762] = 29'b1_111100100010_010_1_111001000101;
      patterns[63763] = 29'b1_111100100010_011_1_110010001011;
      patterns[63764] = 29'b1_111100100010_100_0_111110010001;
      patterns[63765] = 29'b1_111100100010_101_1_011111001000;
      patterns[63766] = 29'b1_111100100010_110_1_111100100010;
      patterns[63767] = 29'b1_111100100010_111_1_111100100010;
      patterns[63768] = 29'b1_111100100011_000_1_111100100011;
      patterns[63769] = 29'b1_111100100011_001_1_100011111100;
      patterns[63770] = 29'b1_111100100011_010_1_111001000111;
      patterns[63771] = 29'b1_111100100011_011_1_110010001111;
      patterns[63772] = 29'b1_111100100011_100_1_111110010001;
      patterns[63773] = 29'b1_111100100011_101_1_111111001000;
      patterns[63774] = 29'b1_111100100011_110_1_111100100011;
      patterns[63775] = 29'b1_111100100011_111_1_111100100011;
      patterns[63776] = 29'b1_111100100100_000_1_111100100100;
      patterns[63777] = 29'b1_111100100100_001_1_100100111100;
      patterns[63778] = 29'b1_111100100100_010_1_111001001001;
      patterns[63779] = 29'b1_111100100100_011_1_110010010011;
      patterns[63780] = 29'b1_111100100100_100_0_111110010010;
      patterns[63781] = 29'b1_111100100100_101_0_011111001001;
      patterns[63782] = 29'b1_111100100100_110_1_111100100100;
      patterns[63783] = 29'b1_111100100100_111_1_111100100100;
      patterns[63784] = 29'b1_111100100101_000_1_111100100101;
      patterns[63785] = 29'b1_111100100101_001_1_100101111100;
      patterns[63786] = 29'b1_111100100101_010_1_111001001011;
      patterns[63787] = 29'b1_111100100101_011_1_110010010111;
      patterns[63788] = 29'b1_111100100101_100_1_111110010010;
      patterns[63789] = 29'b1_111100100101_101_0_111111001001;
      patterns[63790] = 29'b1_111100100101_110_1_111100100101;
      patterns[63791] = 29'b1_111100100101_111_1_111100100101;
      patterns[63792] = 29'b1_111100100110_000_1_111100100110;
      patterns[63793] = 29'b1_111100100110_001_1_100110111100;
      patterns[63794] = 29'b1_111100100110_010_1_111001001101;
      patterns[63795] = 29'b1_111100100110_011_1_110010011011;
      patterns[63796] = 29'b1_111100100110_100_0_111110010011;
      patterns[63797] = 29'b1_111100100110_101_1_011111001001;
      patterns[63798] = 29'b1_111100100110_110_1_111100100110;
      patterns[63799] = 29'b1_111100100110_111_1_111100100110;
      patterns[63800] = 29'b1_111100100111_000_1_111100100111;
      patterns[63801] = 29'b1_111100100111_001_1_100111111100;
      patterns[63802] = 29'b1_111100100111_010_1_111001001111;
      patterns[63803] = 29'b1_111100100111_011_1_110010011111;
      patterns[63804] = 29'b1_111100100111_100_1_111110010011;
      patterns[63805] = 29'b1_111100100111_101_1_111111001001;
      patterns[63806] = 29'b1_111100100111_110_1_111100100111;
      patterns[63807] = 29'b1_111100100111_111_1_111100100111;
      patterns[63808] = 29'b1_111100101000_000_1_111100101000;
      patterns[63809] = 29'b1_111100101000_001_1_101000111100;
      patterns[63810] = 29'b1_111100101000_010_1_111001010001;
      patterns[63811] = 29'b1_111100101000_011_1_110010100011;
      patterns[63812] = 29'b1_111100101000_100_0_111110010100;
      patterns[63813] = 29'b1_111100101000_101_0_011111001010;
      patterns[63814] = 29'b1_111100101000_110_1_111100101000;
      patterns[63815] = 29'b1_111100101000_111_1_111100101000;
      patterns[63816] = 29'b1_111100101001_000_1_111100101001;
      patterns[63817] = 29'b1_111100101001_001_1_101001111100;
      patterns[63818] = 29'b1_111100101001_010_1_111001010011;
      patterns[63819] = 29'b1_111100101001_011_1_110010100111;
      patterns[63820] = 29'b1_111100101001_100_1_111110010100;
      patterns[63821] = 29'b1_111100101001_101_0_111111001010;
      patterns[63822] = 29'b1_111100101001_110_1_111100101001;
      patterns[63823] = 29'b1_111100101001_111_1_111100101001;
      patterns[63824] = 29'b1_111100101010_000_1_111100101010;
      patterns[63825] = 29'b1_111100101010_001_1_101010111100;
      patterns[63826] = 29'b1_111100101010_010_1_111001010101;
      patterns[63827] = 29'b1_111100101010_011_1_110010101011;
      patterns[63828] = 29'b1_111100101010_100_0_111110010101;
      patterns[63829] = 29'b1_111100101010_101_1_011111001010;
      patterns[63830] = 29'b1_111100101010_110_1_111100101010;
      patterns[63831] = 29'b1_111100101010_111_1_111100101010;
      patterns[63832] = 29'b1_111100101011_000_1_111100101011;
      patterns[63833] = 29'b1_111100101011_001_1_101011111100;
      patterns[63834] = 29'b1_111100101011_010_1_111001010111;
      patterns[63835] = 29'b1_111100101011_011_1_110010101111;
      patterns[63836] = 29'b1_111100101011_100_1_111110010101;
      patterns[63837] = 29'b1_111100101011_101_1_111111001010;
      patterns[63838] = 29'b1_111100101011_110_1_111100101011;
      patterns[63839] = 29'b1_111100101011_111_1_111100101011;
      patterns[63840] = 29'b1_111100101100_000_1_111100101100;
      patterns[63841] = 29'b1_111100101100_001_1_101100111100;
      patterns[63842] = 29'b1_111100101100_010_1_111001011001;
      patterns[63843] = 29'b1_111100101100_011_1_110010110011;
      patterns[63844] = 29'b1_111100101100_100_0_111110010110;
      patterns[63845] = 29'b1_111100101100_101_0_011111001011;
      patterns[63846] = 29'b1_111100101100_110_1_111100101100;
      patterns[63847] = 29'b1_111100101100_111_1_111100101100;
      patterns[63848] = 29'b1_111100101101_000_1_111100101101;
      patterns[63849] = 29'b1_111100101101_001_1_101101111100;
      patterns[63850] = 29'b1_111100101101_010_1_111001011011;
      patterns[63851] = 29'b1_111100101101_011_1_110010110111;
      patterns[63852] = 29'b1_111100101101_100_1_111110010110;
      patterns[63853] = 29'b1_111100101101_101_0_111111001011;
      patterns[63854] = 29'b1_111100101101_110_1_111100101101;
      patterns[63855] = 29'b1_111100101101_111_1_111100101101;
      patterns[63856] = 29'b1_111100101110_000_1_111100101110;
      patterns[63857] = 29'b1_111100101110_001_1_101110111100;
      patterns[63858] = 29'b1_111100101110_010_1_111001011101;
      patterns[63859] = 29'b1_111100101110_011_1_110010111011;
      patterns[63860] = 29'b1_111100101110_100_0_111110010111;
      patterns[63861] = 29'b1_111100101110_101_1_011111001011;
      patterns[63862] = 29'b1_111100101110_110_1_111100101110;
      patterns[63863] = 29'b1_111100101110_111_1_111100101110;
      patterns[63864] = 29'b1_111100101111_000_1_111100101111;
      patterns[63865] = 29'b1_111100101111_001_1_101111111100;
      patterns[63866] = 29'b1_111100101111_010_1_111001011111;
      patterns[63867] = 29'b1_111100101111_011_1_110010111111;
      patterns[63868] = 29'b1_111100101111_100_1_111110010111;
      patterns[63869] = 29'b1_111100101111_101_1_111111001011;
      patterns[63870] = 29'b1_111100101111_110_1_111100101111;
      patterns[63871] = 29'b1_111100101111_111_1_111100101111;
      patterns[63872] = 29'b1_111100110000_000_1_111100110000;
      patterns[63873] = 29'b1_111100110000_001_1_110000111100;
      patterns[63874] = 29'b1_111100110000_010_1_111001100001;
      patterns[63875] = 29'b1_111100110000_011_1_110011000011;
      patterns[63876] = 29'b1_111100110000_100_0_111110011000;
      patterns[63877] = 29'b1_111100110000_101_0_011111001100;
      patterns[63878] = 29'b1_111100110000_110_1_111100110000;
      patterns[63879] = 29'b1_111100110000_111_1_111100110000;
      patterns[63880] = 29'b1_111100110001_000_1_111100110001;
      patterns[63881] = 29'b1_111100110001_001_1_110001111100;
      patterns[63882] = 29'b1_111100110001_010_1_111001100011;
      patterns[63883] = 29'b1_111100110001_011_1_110011000111;
      patterns[63884] = 29'b1_111100110001_100_1_111110011000;
      patterns[63885] = 29'b1_111100110001_101_0_111111001100;
      patterns[63886] = 29'b1_111100110001_110_1_111100110001;
      patterns[63887] = 29'b1_111100110001_111_1_111100110001;
      patterns[63888] = 29'b1_111100110010_000_1_111100110010;
      patterns[63889] = 29'b1_111100110010_001_1_110010111100;
      patterns[63890] = 29'b1_111100110010_010_1_111001100101;
      patterns[63891] = 29'b1_111100110010_011_1_110011001011;
      patterns[63892] = 29'b1_111100110010_100_0_111110011001;
      patterns[63893] = 29'b1_111100110010_101_1_011111001100;
      patterns[63894] = 29'b1_111100110010_110_1_111100110010;
      patterns[63895] = 29'b1_111100110010_111_1_111100110010;
      patterns[63896] = 29'b1_111100110011_000_1_111100110011;
      patterns[63897] = 29'b1_111100110011_001_1_110011111100;
      patterns[63898] = 29'b1_111100110011_010_1_111001100111;
      patterns[63899] = 29'b1_111100110011_011_1_110011001111;
      patterns[63900] = 29'b1_111100110011_100_1_111110011001;
      patterns[63901] = 29'b1_111100110011_101_1_111111001100;
      patterns[63902] = 29'b1_111100110011_110_1_111100110011;
      patterns[63903] = 29'b1_111100110011_111_1_111100110011;
      patterns[63904] = 29'b1_111100110100_000_1_111100110100;
      patterns[63905] = 29'b1_111100110100_001_1_110100111100;
      patterns[63906] = 29'b1_111100110100_010_1_111001101001;
      patterns[63907] = 29'b1_111100110100_011_1_110011010011;
      patterns[63908] = 29'b1_111100110100_100_0_111110011010;
      patterns[63909] = 29'b1_111100110100_101_0_011111001101;
      patterns[63910] = 29'b1_111100110100_110_1_111100110100;
      patterns[63911] = 29'b1_111100110100_111_1_111100110100;
      patterns[63912] = 29'b1_111100110101_000_1_111100110101;
      patterns[63913] = 29'b1_111100110101_001_1_110101111100;
      patterns[63914] = 29'b1_111100110101_010_1_111001101011;
      patterns[63915] = 29'b1_111100110101_011_1_110011010111;
      patterns[63916] = 29'b1_111100110101_100_1_111110011010;
      patterns[63917] = 29'b1_111100110101_101_0_111111001101;
      patterns[63918] = 29'b1_111100110101_110_1_111100110101;
      patterns[63919] = 29'b1_111100110101_111_1_111100110101;
      patterns[63920] = 29'b1_111100110110_000_1_111100110110;
      patterns[63921] = 29'b1_111100110110_001_1_110110111100;
      patterns[63922] = 29'b1_111100110110_010_1_111001101101;
      patterns[63923] = 29'b1_111100110110_011_1_110011011011;
      patterns[63924] = 29'b1_111100110110_100_0_111110011011;
      patterns[63925] = 29'b1_111100110110_101_1_011111001101;
      patterns[63926] = 29'b1_111100110110_110_1_111100110110;
      patterns[63927] = 29'b1_111100110110_111_1_111100110110;
      patterns[63928] = 29'b1_111100110111_000_1_111100110111;
      patterns[63929] = 29'b1_111100110111_001_1_110111111100;
      patterns[63930] = 29'b1_111100110111_010_1_111001101111;
      patterns[63931] = 29'b1_111100110111_011_1_110011011111;
      patterns[63932] = 29'b1_111100110111_100_1_111110011011;
      patterns[63933] = 29'b1_111100110111_101_1_111111001101;
      patterns[63934] = 29'b1_111100110111_110_1_111100110111;
      patterns[63935] = 29'b1_111100110111_111_1_111100110111;
      patterns[63936] = 29'b1_111100111000_000_1_111100111000;
      patterns[63937] = 29'b1_111100111000_001_1_111000111100;
      patterns[63938] = 29'b1_111100111000_010_1_111001110001;
      patterns[63939] = 29'b1_111100111000_011_1_110011100011;
      patterns[63940] = 29'b1_111100111000_100_0_111110011100;
      patterns[63941] = 29'b1_111100111000_101_0_011111001110;
      patterns[63942] = 29'b1_111100111000_110_1_111100111000;
      patterns[63943] = 29'b1_111100111000_111_1_111100111000;
      patterns[63944] = 29'b1_111100111001_000_1_111100111001;
      patterns[63945] = 29'b1_111100111001_001_1_111001111100;
      patterns[63946] = 29'b1_111100111001_010_1_111001110011;
      patterns[63947] = 29'b1_111100111001_011_1_110011100111;
      patterns[63948] = 29'b1_111100111001_100_1_111110011100;
      patterns[63949] = 29'b1_111100111001_101_0_111111001110;
      patterns[63950] = 29'b1_111100111001_110_1_111100111001;
      patterns[63951] = 29'b1_111100111001_111_1_111100111001;
      patterns[63952] = 29'b1_111100111010_000_1_111100111010;
      patterns[63953] = 29'b1_111100111010_001_1_111010111100;
      patterns[63954] = 29'b1_111100111010_010_1_111001110101;
      patterns[63955] = 29'b1_111100111010_011_1_110011101011;
      patterns[63956] = 29'b1_111100111010_100_0_111110011101;
      patterns[63957] = 29'b1_111100111010_101_1_011111001110;
      patterns[63958] = 29'b1_111100111010_110_1_111100111010;
      patterns[63959] = 29'b1_111100111010_111_1_111100111010;
      patterns[63960] = 29'b1_111100111011_000_1_111100111011;
      patterns[63961] = 29'b1_111100111011_001_1_111011111100;
      patterns[63962] = 29'b1_111100111011_010_1_111001110111;
      patterns[63963] = 29'b1_111100111011_011_1_110011101111;
      patterns[63964] = 29'b1_111100111011_100_1_111110011101;
      patterns[63965] = 29'b1_111100111011_101_1_111111001110;
      patterns[63966] = 29'b1_111100111011_110_1_111100111011;
      patterns[63967] = 29'b1_111100111011_111_1_111100111011;
      patterns[63968] = 29'b1_111100111100_000_1_111100111100;
      patterns[63969] = 29'b1_111100111100_001_1_111100111100;
      patterns[63970] = 29'b1_111100111100_010_1_111001111001;
      patterns[63971] = 29'b1_111100111100_011_1_110011110011;
      patterns[63972] = 29'b1_111100111100_100_0_111110011110;
      patterns[63973] = 29'b1_111100111100_101_0_011111001111;
      patterns[63974] = 29'b1_111100111100_110_1_111100111100;
      patterns[63975] = 29'b1_111100111100_111_1_111100111100;
      patterns[63976] = 29'b1_111100111101_000_1_111100111101;
      patterns[63977] = 29'b1_111100111101_001_1_111101111100;
      patterns[63978] = 29'b1_111100111101_010_1_111001111011;
      patterns[63979] = 29'b1_111100111101_011_1_110011110111;
      patterns[63980] = 29'b1_111100111101_100_1_111110011110;
      patterns[63981] = 29'b1_111100111101_101_0_111111001111;
      patterns[63982] = 29'b1_111100111101_110_1_111100111101;
      patterns[63983] = 29'b1_111100111101_111_1_111100111101;
      patterns[63984] = 29'b1_111100111110_000_1_111100111110;
      patterns[63985] = 29'b1_111100111110_001_1_111110111100;
      patterns[63986] = 29'b1_111100111110_010_1_111001111101;
      patterns[63987] = 29'b1_111100111110_011_1_110011111011;
      patterns[63988] = 29'b1_111100111110_100_0_111110011111;
      patterns[63989] = 29'b1_111100111110_101_1_011111001111;
      patterns[63990] = 29'b1_111100111110_110_1_111100111110;
      patterns[63991] = 29'b1_111100111110_111_1_111100111110;
      patterns[63992] = 29'b1_111100111111_000_1_111100111111;
      patterns[63993] = 29'b1_111100111111_001_1_111111111100;
      patterns[63994] = 29'b1_111100111111_010_1_111001111111;
      patterns[63995] = 29'b1_111100111111_011_1_110011111111;
      patterns[63996] = 29'b1_111100111111_100_1_111110011111;
      patterns[63997] = 29'b1_111100111111_101_1_111111001111;
      patterns[63998] = 29'b1_111100111111_110_1_111100111111;
      patterns[63999] = 29'b1_111100111111_111_1_111100111111;
      patterns[64000] = 29'b1_111101000000_000_1_111101000000;
      patterns[64001] = 29'b1_111101000000_001_1_000000111101;
      patterns[64002] = 29'b1_111101000000_010_1_111010000001;
      patterns[64003] = 29'b1_111101000000_011_1_110100000011;
      patterns[64004] = 29'b1_111101000000_100_0_111110100000;
      patterns[64005] = 29'b1_111101000000_101_0_011111010000;
      patterns[64006] = 29'b1_111101000000_110_1_111101000000;
      patterns[64007] = 29'b1_111101000000_111_1_111101000000;
      patterns[64008] = 29'b1_111101000001_000_1_111101000001;
      patterns[64009] = 29'b1_111101000001_001_1_000001111101;
      patterns[64010] = 29'b1_111101000001_010_1_111010000011;
      patterns[64011] = 29'b1_111101000001_011_1_110100000111;
      patterns[64012] = 29'b1_111101000001_100_1_111110100000;
      patterns[64013] = 29'b1_111101000001_101_0_111111010000;
      patterns[64014] = 29'b1_111101000001_110_1_111101000001;
      patterns[64015] = 29'b1_111101000001_111_1_111101000001;
      patterns[64016] = 29'b1_111101000010_000_1_111101000010;
      patterns[64017] = 29'b1_111101000010_001_1_000010111101;
      patterns[64018] = 29'b1_111101000010_010_1_111010000101;
      patterns[64019] = 29'b1_111101000010_011_1_110100001011;
      patterns[64020] = 29'b1_111101000010_100_0_111110100001;
      patterns[64021] = 29'b1_111101000010_101_1_011111010000;
      patterns[64022] = 29'b1_111101000010_110_1_111101000010;
      patterns[64023] = 29'b1_111101000010_111_1_111101000010;
      patterns[64024] = 29'b1_111101000011_000_1_111101000011;
      patterns[64025] = 29'b1_111101000011_001_1_000011111101;
      patterns[64026] = 29'b1_111101000011_010_1_111010000111;
      patterns[64027] = 29'b1_111101000011_011_1_110100001111;
      patterns[64028] = 29'b1_111101000011_100_1_111110100001;
      patterns[64029] = 29'b1_111101000011_101_1_111111010000;
      patterns[64030] = 29'b1_111101000011_110_1_111101000011;
      patterns[64031] = 29'b1_111101000011_111_1_111101000011;
      patterns[64032] = 29'b1_111101000100_000_1_111101000100;
      patterns[64033] = 29'b1_111101000100_001_1_000100111101;
      patterns[64034] = 29'b1_111101000100_010_1_111010001001;
      patterns[64035] = 29'b1_111101000100_011_1_110100010011;
      patterns[64036] = 29'b1_111101000100_100_0_111110100010;
      patterns[64037] = 29'b1_111101000100_101_0_011111010001;
      patterns[64038] = 29'b1_111101000100_110_1_111101000100;
      patterns[64039] = 29'b1_111101000100_111_1_111101000100;
      patterns[64040] = 29'b1_111101000101_000_1_111101000101;
      patterns[64041] = 29'b1_111101000101_001_1_000101111101;
      patterns[64042] = 29'b1_111101000101_010_1_111010001011;
      patterns[64043] = 29'b1_111101000101_011_1_110100010111;
      patterns[64044] = 29'b1_111101000101_100_1_111110100010;
      patterns[64045] = 29'b1_111101000101_101_0_111111010001;
      patterns[64046] = 29'b1_111101000101_110_1_111101000101;
      patterns[64047] = 29'b1_111101000101_111_1_111101000101;
      patterns[64048] = 29'b1_111101000110_000_1_111101000110;
      patterns[64049] = 29'b1_111101000110_001_1_000110111101;
      patterns[64050] = 29'b1_111101000110_010_1_111010001101;
      patterns[64051] = 29'b1_111101000110_011_1_110100011011;
      patterns[64052] = 29'b1_111101000110_100_0_111110100011;
      patterns[64053] = 29'b1_111101000110_101_1_011111010001;
      patterns[64054] = 29'b1_111101000110_110_1_111101000110;
      patterns[64055] = 29'b1_111101000110_111_1_111101000110;
      patterns[64056] = 29'b1_111101000111_000_1_111101000111;
      patterns[64057] = 29'b1_111101000111_001_1_000111111101;
      patterns[64058] = 29'b1_111101000111_010_1_111010001111;
      patterns[64059] = 29'b1_111101000111_011_1_110100011111;
      patterns[64060] = 29'b1_111101000111_100_1_111110100011;
      patterns[64061] = 29'b1_111101000111_101_1_111111010001;
      patterns[64062] = 29'b1_111101000111_110_1_111101000111;
      patterns[64063] = 29'b1_111101000111_111_1_111101000111;
      patterns[64064] = 29'b1_111101001000_000_1_111101001000;
      patterns[64065] = 29'b1_111101001000_001_1_001000111101;
      patterns[64066] = 29'b1_111101001000_010_1_111010010001;
      patterns[64067] = 29'b1_111101001000_011_1_110100100011;
      patterns[64068] = 29'b1_111101001000_100_0_111110100100;
      patterns[64069] = 29'b1_111101001000_101_0_011111010010;
      patterns[64070] = 29'b1_111101001000_110_1_111101001000;
      patterns[64071] = 29'b1_111101001000_111_1_111101001000;
      patterns[64072] = 29'b1_111101001001_000_1_111101001001;
      patterns[64073] = 29'b1_111101001001_001_1_001001111101;
      patterns[64074] = 29'b1_111101001001_010_1_111010010011;
      patterns[64075] = 29'b1_111101001001_011_1_110100100111;
      patterns[64076] = 29'b1_111101001001_100_1_111110100100;
      patterns[64077] = 29'b1_111101001001_101_0_111111010010;
      patterns[64078] = 29'b1_111101001001_110_1_111101001001;
      patterns[64079] = 29'b1_111101001001_111_1_111101001001;
      patterns[64080] = 29'b1_111101001010_000_1_111101001010;
      patterns[64081] = 29'b1_111101001010_001_1_001010111101;
      patterns[64082] = 29'b1_111101001010_010_1_111010010101;
      patterns[64083] = 29'b1_111101001010_011_1_110100101011;
      patterns[64084] = 29'b1_111101001010_100_0_111110100101;
      patterns[64085] = 29'b1_111101001010_101_1_011111010010;
      patterns[64086] = 29'b1_111101001010_110_1_111101001010;
      patterns[64087] = 29'b1_111101001010_111_1_111101001010;
      patterns[64088] = 29'b1_111101001011_000_1_111101001011;
      patterns[64089] = 29'b1_111101001011_001_1_001011111101;
      patterns[64090] = 29'b1_111101001011_010_1_111010010111;
      patterns[64091] = 29'b1_111101001011_011_1_110100101111;
      patterns[64092] = 29'b1_111101001011_100_1_111110100101;
      patterns[64093] = 29'b1_111101001011_101_1_111111010010;
      patterns[64094] = 29'b1_111101001011_110_1_111101001011;
      patterns[64095] = 29'b1_111101001011_111_1_111101001011;
      patterns[64096] = 29'b1_111101001100_000_1_111101001100;
      patterns[64097] = 29'b1_111101001100_001_1_001100111101;
      patterns[64098] = 29'b1_111101001100_010_1_111010011001;
      patterns[64099] = 29'b1_111101001100_011_1_110100110011;
      patterns[64100] = 29'b1_111101001100_100_0_111110100110;
      patterns[64101] = 29'b1_111101001100_101_0_011111010011;
      patterns[64102] = 29'b1_111101001100_110_1_111101001100;
      patterns[64103] = 29'b1_111101001100_111_1_111101001100;
      patterns[64104] = 29'b1_111101001101_000_1_111101001101;
      patterns[64105] = 29'b1_111101001101_001_1_001101111101;
      patterns[64106] = 29'b1_111101001101_010_1_111010011011;
      patterns[64107] = 29'b1_111101001101_011_1_110100110111;
      patterns[64108] = 29'b1_111101001101_100_1_111110100110;
      patterns[64109] = 29'b1_111101001101_101_0_111111010011;
      patterns[64110] = 29'b1_111101001101_110_1_111101001101;
      patterns[64111] = 29'b1_111101001101_111_1_111101001101;
      patterns[64112] = 29'b1_111101001110_000_1_111101001110;
      patterns[64113] = 29'b1_111101001110_001_1_001110111101;
      patterns[64114] = 29'b1_111101001110_010_1_111010011101;
      patterns[64115] = 29'b1_111101001110_011_1_110100111011;
      patterns[64116] = 29'b1_111101001110_100_0_111110100111;
      patterns[64117] = 29'b1_111101001110_101_1_011111010011;
      patterns[64118] = 29'b1_111101001110_110_1_111101001110;
      patterns[64119] = 29'b1_111101001110_111_1_111101001110;
      patterns[64120] = 29'b1_111101001111_000_1_111101001111;
      patterns[64121] = 29'b1_111101001111_001_1_001111111101;
      patterns[64122] = 29'b1_111101001111_010_1_111010011111;
      patterns[64123] = 29'b1_111101001111_011_1_110100111111;
      patterns[64124] = 29'b1_111101001111_100_1_111110100111;
      patterns[64125] = 29'b1_111101001111_101_1_111111010011;
      patterns[64126] = 29'b1_111101001111_110_1_111101001111;
      patterns[64127] = 29'b1_111101001111_111_1_111101001111;
      patterns[64128] = 29'b1_111101010000_000_1_111101010000;
      patterns[64129] = 29'b1_111101010000_001_1_010000111101;
      patterns[64130] = 29'b1_111101010000_010_1_111010100001;
      patterns[64131] = 29'b1_111101010000_011_1_110101000011;
      patterns[64132] = 29'b1_111101010000_100_0_111110101000;
      patterns[64133] = 29'b1_111101010000_101_0_011111010100;
      patterns[64134] = 29'b1_111101010000_110_1_111101010000;
      patterns[64135] = 29'b1_111101010000_111_1_111101010000;
      patterns[64136] = 29'b1_111101010001_000_1_111101010001;
      patterns[64137] = 29'b1_111101010001_001_1_010001111101;
      patterns[64138] = 29'b1_111101010001_010_1_111010100011;
      patterns[64139] = 29'b1_111101010001_011_1_110101000111;
      patterns[64140] = 29'b1_111101010001_100_1_111110101000;
      patterns[64141] = 29'b1_111101010001_101_0_111111010100;
      patterns[64142] = 29'b1_111101010001_110_1_111101010001;
      patterns[64143] = 29'b1_111101010001_111_1_111101010001;
      patterns[64144] = 29'b1_111101010010_000_1_111101010010;
      patterns[64145] = 29'b1_111101010010_001_1_010010111101;
      patterns[64146] = 29'b1_111101010010_010_1_111010100101;
      patterns[64147] = 29'b1_111101010010_011_1_110101001011;
      patterns[64148] = 29'b1_111101010010_100_0_111110101001;
      patterns[64149] = 29'b1_111101010010_101_1_011111010100;
      patterns[64150] = 29'b1_111101010010_110_1_111101010010;
      patterns[64151] = 29'b1_111101010010_111_1_111101010010;
      patterns[64152] = 29'b1_111101010011_000_1_111101010011;
      patterns[64153] = 29'b1_111101010011_001_1_010011111101;
      patterns[64154] = 29'b1_111101010011_010_1_111010100111;
      patterns[64155] = 29'b1_111101010011_011_1_110101001111;
      patterns[64156] = 29'b1_111101010011_100_1_111110101001;
      patterns[64157] = 29'b1_111101010011_101_1_111111010100;
      patterns[64158] = 29'b1_111101010011_110_1_111101010011;
      patterns[64159] = 29'b1_111101010011_111_1_111101010011;
      patterns[64160] = 29'b1_111101010100_000_1_111101010100;
      patterns[64161] = 29'b1_111101010100_001_1_010100111101;
      patterns[64162] = 29'b1_111101010100_010_1_111010101001;
      patterns[64163] = 29'b1_111101010100_011_1_110101010011;
      patterns[64164] = 29'b1_111101010100_100_0_111110101010;
      patterns[64165] = 29'b1_111101010100_101_0_011111010101;
      patterns[64166] = 29'b1_111101010100_110_1_111101010100;
      patterns[64167] = 29'b1_111101010100_111_1_111101010100;
      patterns[64168] = 29'b1_111101010101_000_1_111101010101;
      patterns[64169] = 29'b1_111101010101_001_1_010101111101;
      patterns[64170] = 29'b1_111101010101_010_1_111010101011;
      patterns[64171] = 29'b1_111101010101_011_1_110101010111;
      patterns[64172] = 29'b1_111101010101_100_1_111110101010;
      patterns[64173] = 29'b1_111101010101_101_0_111111010101;
      patterns[64174] = 29'b1_111101010101_110_1_111101010101;
      patterns[64175] = 29'b1_111101010101_111_1_111101010101;
      patterns[64176] = 29'b1_111101010110_000_1_111101010110;
      patterns[64177] = 29'b1_111101010110_001_1_010110111101;
      patterns[64178] = 29'b1_111101010110_010_1_111010101101;
      patterns[64179] = 29'b1_111101010110_011_1_110101011011;
      patterns[64180] = 29'b1_111101010110_100_0_111110101011;
      patterns[64181] = 29'b1_111101010110_101_1_011111010101;
      patterns[64182] = 29'b1_111101010110_110_1_111101010110;
      patterns[64183] = 29'b1_111101010110_111_1_111101010110;
      patterns[64184] = 29'b1_111101010111_000_1_111101010111;
      patterns[64185] = 29'b1_111101010111_001_1_010111111101;
      patterns[64186] = 29'b1_111101010111_010_1_111010101111;
      patterns[64187] = 29'b1_111101010111_011_1_110101011111;
      patterns[64188] = 29'b1_111101010111_100_1_111110101011;
      patterns[64189] = 29'b1_111101010111_101_1_111111010101;
      patterns[64190] = 29'b1_111101010111_110_1_111101010111;
      patterns[64191] = 29'b1_111101010111_111_1_111101010111;
      patterns[64192] = 29'b1_111101011000_000_1_111101011000;
      patterns[64193] = 29'b1_111101011000_001_1_011000111101;
      patterns[64194] = 29'b1_111101011000_010_1_111010110001;
      patterns[64195] = 29'b1_111101011000_011_1_110101100011;
      patterns[64196] = 29'b1_111101011000_100_0_111110101100;
      patterns[64197] = 29'b1_111101011000_101_0_011111010110;
      patterns[64198] = 29'b1_111101011000_110_1_111101011000;
      patterns[64199] = 29'b1_111101011000_111_1_111101011000;
      patterns[64200] = 29'b1_111101011001_000_1_111101011001;
      patterns[64201] = 29'b1_111101011001_001_1_011001111101;
      patterns[64202] = 29'b1_111101011001_010_1_111010110011;
      patterns[64203] = 29'b1_111101011001_011_1_110101100111;
      patterns[64204] = 29'b1_111101011001_100_1_111110101100;
      patterns[64205] = 29'b1_111101011001_101_0_111111010110;
      patterns[64206] = 29'b1_111101011001_110_1_111101011001;
      patterns[64207] = 29'b1_111101011001_111_1_111101011001;
      patterns[64208] = 29'b1_111101011010_000_1_111101011010;
      patterns[64209] = 29'b1_111101011010_001_1_011010111101;
      patterns[64210] = 29'b1_111101011010_010_1_111010110101;
      patterns[64211] = 29'b1_111101011010_011_1_110101101011;
      patterns[64212] = 29'b1_111101011010_100_0_111110101101;
      patterns[64213] = 29'b1_111101011010_101_1_011111010110;
      patterns[64214] = 29'b1_111101011010_110_1_111101011010;
      patterns[64215] = 29'b1_111101011010_111_1_111101011010;
      patterns[64216] = 29'b1_111101011011_000_1_111101011011;
      patterns[64217] = 29'b1_111101011011_001_1_011011111101;
      patterns[64218] = 29'b1_111101011011_010_1_111010110111;
      patterns[64219] = 29'b1_111101011011_011_1_110101101111;
      patterns[64220] = 29'b1_111101011011_100_1_111110101101;
      patterns[64221] = 29'b1_111101011011_101_1_111111010110;
      patterns[64222] = 29'b1_111101011011_110_1_111101011011;
      patterns[64223] = 29'b1_111101011011_111_1_111101011011;
      patterns[64224] = 29'b1_111101011100_000_1_111101011100;
      patterns[64225] = 29'b1_111101011100_001_1_011100111101;
      patterns[64226] = 29'b1_111101011100_010_1_111010111001;
      patterns[64227] = 29'b1_111101011100_011_1_110101110011;
      patterns[64228] = 29'b1_111101011100_100_0_111110101110;
      patterns[64229] = 29'b1_111101011100_101_0_011111010111;
      patterns[64230] = 29'b1_111101011100_110_1_111101011100;
      patterns[64231] = 29'b1_111101011100_111_1_111101011100;
      patterns[64232] = 29'b1_111101011101_000_1_111101011101;
      patterns[64233] = 29'b1_111101011101_001_1_011101111101;
      patterns[64234] = 29'b1_111101011101_010_1_111010111011;
      patterns[64235] = 29'b1_111101011101_011_1_110101110111;
      patterns[64236] = 29'b1_111101011101_100_1_111110101110;
      patterns[64237] = 29'b1_111101011101_101_0_111111010111;
      patterns[64238] = 29'b1_111101011101_110_1_111101011101;
      patterns[64239] = 29'b1_111101011101_111_1_111101011101;
      patterns[64240] = 29'b1_111101011110_000_1_111101011110;
      patterns[64241] = 29'b1_111101011110_001_1_011110111101;
      patterns[64242] = 29'b1_111101011110_010_1_111010111101;
      patterns[64243] = 29'b1_111101011110_011_1_110101111011;
      patterns[64244] = 29'b1_111101011110_100_0_111110101111;
      patterns[64245] = 29'b1_111101011110_101_1_011111010111;
      patterns[64246] = 29'b1_111101011110_110_1_111101011110;
      patterns[64247] = 29'b1_111101011110_111_1_111101011110;
      patterns[64248] = 29'b1_111101011111_000_1_111101011111;
      patterns[64249] = 29'b1_111101011111_001_1_011111111101;
      patterns[64250] = 29'b1_111101011111_010_1_111010111111;
      patterns[64251] = 29'b1_111101011111_011_1_110101111111;
      patterns[64252] = 29'b1_111101011111_100_1_111110101111;
      patterns[64253] = 29'b1_111101011111_101_1_111111010111;
      patterns[64254] = 29'b1_111101011111_110_1_111101011111;
      patterns[64255] = 29'b1_111101011111_111_1_111101011111;
      patterns[64256] = 29'b1_111101100000_000_1_111101100000;
      patterns[64257] = 29'b1_111101100000_001_1_100000111101;
      patterns[64258] = 29'b1_111101100000_010_1_111011000001;
      patterns[64259] = 29'b1_111101100000_011_1_110110000011;
      patterns[64260] = 29'b1_111101100000_100_0_111110110000;
      patterns[64261] = 29'b1_111101100000_101_0_011111011000;
      patterns[64262] = 29'b1_111101100000_110_1_111101100000;
      patterns[64263] = 29'b1_111101100000_111_1_111101100000;
      patterns[64264] = 29'b1_111101100001_000_1_111101100001;
      patterns[64265] = 29'b1_111101100001_001_1_100001111101;
      patterns[64266] = 29'b1_111101100001_010_1_111011000011;
      patterns[64267] = 29'b1_111101100001_011_1_110110000111;
      patterns[64268] = 29'b1_111101100001_100_1_111110110000;
      patterns[64269] = 29'b1_111101100001_101_0_111111011000;
      patterns[64270] = 29'b1_111101100001_110_1_111101100001;
      patterns[64271] = 29'b1_111101100001_111_1_111101100001;
      patterns[64272] = 29'b1_111101100010_000_1_111101100010;
      patterns[64273] = 29'b1_111101100010_001_1_100010111101;
      patterns[64274] = 29'b1_111101100010_010_1_111011000101;
      patterns[64275] = 29'b1_111101100010_011_1_110110001011;
      patterns[64276] = 29'b1_111101100010_100_0_111110110001;
      patterns[64277] = 29'b1_111101100010_101_1_011111011000;
      patterns[64278] = 29'b1_111101100010_110_1_111101100010;
      patterns[64279] = 29'b1_111101100010_111_1_111101100010;
      patterns[64280] = 29'b1_111101100011_000_1_111101100011;
      patterns[64281] = 29'b1_111101100011_001_1_100011111101;
      patterns[64282] = 29'b1_111101100011_010_1_111011000111;
      patterns[64283] = 29'b1_111101100011_011_1_110110001111;
      patterns[64284] = 29'b1_111101100011_100_1_111110110001;
      patterns[64285] = 29'b1_111101100011_101_1_111111011000;
      patterns[64286] = 29'b1_111101100011_110_1_111101100011;
      patterns[64287] = 29'b1_111101100011_111_1_111101100011;
      patterns[64288] = 29'b1_111101100100_000_1_111101100100;
      patterns[64289] = 29'b1_111101100100_001_1_100100111101;
      patterns[64290] = 29'b1_111101100100_010_1_111011001001;
      patterns[64291] = 29'b1_111101100100_011_1_110110010011;
      patterns[64292] = 29'b1_111101100100_100_0_111110110010;
      patterns[64293] = 29'b1_111101100100_101_0_011111011001;
      patterns[64294] = 29'b1_111101100100_110_1_111101100100;
      patterns[64295] = 29'b1_111101100100_111_1_111101100100;
      patterns[64296] = 29'b1_111101100101_000_1_111101100101;
      patterns[64297] = 29'b1_111101100101_001_1_100101111101;
      patterns[64298] = 29'b1_111101100101_010_1_111011001011;
      patterns[64299] = 29'b1_111101100101_011_1_110110010111;
      patterns[64300] = 29'b1_111101100101_100_1_111110110010;
      patterns[64301] = 29'b1_111101100101_101_0_111111011001;
      patterns[64302] = 29'b1_111101100101_110_1_111101100101;
      patterns[64303] = 29'b1_111101100101_111_1_111101100101;
      patterns[64304] = 29'b1_111101100110_000_1_111101100110;
      patterns[64305] = 29'b1_111101100110_001_1_100110111101;
      patterns[64306] = 29'b1_111101100110_010_1_111011001101;
      patterns[64307] = 29'b1_111101100110_011_1_110110011011;
      patterns[64308] = 29'b1_111101100110_100_0_111110110011;
      patterns[64309] = 29'b1_111101100110_101_1_011111011001;
      patterns[64310] = 29'b1_111101100110_110_1_111101100110;
      patterns[64311] = 29'b1_111101100110_111_1_111101100110;
      patterns[64312] = 29'b1_111101100111_000_1_111101100111;
      patterns[64313] = 29'b1_111101100111_001_1_100111111101;
      patterns[64314] = 29'b1_111101100111_010_1_111011001111;
      patterns[64315] = 29'b1_111101100111_011_1_110110011111;
      patterns[64316] = 29'b1_111101100111_100_1_111110110011;
      patterns[64317] = 29'b1_111101100111_101_1_111111011001;
      patterns[64318] = 29'b1_111101100111_110_1_111101100111;
      patterns[64319] = 29'b1_111101100111_111_1_111101100111;
      patterns[64320] = 29'b1_111101101000_000_1_111101101000;
      patterns[64321] = 29'b1_111101101000_001_1_101000111101;
      patterns[64322] = 29'b1_111101101000_010_1_111011010001;
      patterns[64323] = 29'b1_111101101000_011_1_110110100011;
      patterns[64324] = 29'b1_111101101000_100_0_111110110100;
      patterns[64325] = 29'b1_111101101000_101_0_011111011010;
      patterns[64326] = 29'b1_111101101000_110_1_111101101000;
      patterns[64327] = 29'b1_111101101000_111_1_111101101000;
      patterns[64328] = 29'b1_111101101001_000_1_111101101001;
      patterns[64329] = 29'b1_111101101001_001_1_101001111101;
      patterns[64330] = 29'b1_111101101001_010_1_111011010011;
      patterns[64331] = 29'b1_111101101001_011_1_110110100111;
      patterns[64332] = 29'b1_111101101001_100_1_111110110100;
      patterns[64333] = 29'b1_111101101001_101_0_111111011010;
      patterns[64334] = 29'b1_111101101001_110_1_111101101001;
      patterns[64335] = 29'b1_111101101001_111_1_111101101001;
      patterns[64336] = 29'b1_111101101010_000_1_111101101010;
      patterns[64337] = 29'b1_111101101010_001_1_101010111101;
      patterns[64338] = 29'b1_111101101010_010_1_111011010101;
      patterns[64339] = 29'b1_111101101010_011_1_110110101011;
      patterns[64340] = 29'b1_111101101010_100_0_111110110101;
      patterns[64341] = 29'b1_111101101010_101_1_011111011010;
      patterns[64342] = 29'b1_111101101010_110_1_111101101010;
      patterns[64343] = 29'b1_111101101010_111_1_111101101010;
      patterns[64344] = 29'b1_111101101011_000_1_111101101011;
      patterns[64345] = 29'b1_111101101011_001_1_101011111101;
      patterns[64346] = 29'b1_111101101011_010_1_111011010111;
      patterns[64347] = 29'b1_111101101011_011_1_110110101111;
      patterns[64348] = 29'b1_111101101011_100_1_111110110101;
      patterns[64349] = 29'b1_111101101011_101_1_111111011010;
      patterns[64350] = 29'b1_111101101011_110_1_111101101011;
      patterns[64351] = 29'b1_111101101011_111_1_111101101011;
      patterns[64352] = 29'b1_111101101100_000_1_111101101100;
      patterns[64353] = 29'b1_111101101100_001_1_101100111101;
      patterns[64354] = 29'b1_111101101100_010_1_111011011001;
      patterns[64355] = 29'b1_111101101100_011_1_110110110011;
      patterns[64356] = 29'b1_111101101100_100_0_111110110110;
      patterns[64357] = 29'b1_111101101100_101_0_011111011011;
      patterns[64358] = 29'b1_111101101100_110_1_111101101100;
      patterns[64359] = 29'b1_111101101100_111_1_111101101100;
      patterns[64360] = 29'b1_111101101101_000_1_111101101101;
      patterns[64361] = 29'b1_111101101101_001_1_101101111101;
      patterns[64362] = 29'b1_111101101101_010_1_111011011011;
      patterns[64363] = 29'b1_111101101101_011_1_110110110111;
      patterns[64364] = 29'b1_111101101101_100_1_111110110110;
      patterns[64365] = 29'b1_111101101101_101_0_111111011011;
      patterns[64366] = 29'b1_111101101101_110_1_111101101101;
      patterns[64367] = 29'b1_111101101101_111_1_111101101101;
      patterns[64368] = 29'b1_111101101110_000_1_111101101110;
      patterns[64369] = 29'b1_111101101110_001_1_101110111101;
      patterns[64370] = 29'b1_111101101110_010_1_111011011101;
      patterns[64371] = 29'b1_111101101110_011_1_110110111011;
      patterns[64372] = 29'b1_111101101110_100_0_111110110111;
      patterns[64373] = 29'b1_111101101110_101_1_011111011011;
      patterns[64374] = 29'b1_111101101110_110_1_111101101110;
      patterns[64375] = 29'b1_111101101110_111_1_111101101110;
      patterns[64376] = 29'b1_111101101111_000_1_111101101111;
      patterns[64377] = 29'b1_111101101111_001_1_101111111101;
      patterns[64378] = 29'b1_111101101111_010_1_111011011111;
      patterns[64379] = 29'b1_111101101111_011_1_110110111111;
      patterns[64380] = 29'b1_111101101111_100_1_111110110111;
      patterns[64381] = 29'b1_111101101111_101_1_111111011011;
      patterns[64382] = 29'b1_111101101111_110_1_111101101111;
      patterns[64383] = 29'b1_111101101111_111_1_111101101111;
      patterns[64384] = 29'b1_111101110000_000_1_111101110000;
      patterns[64385] = 29'b1_111101110000_001_1_110000111101;
      patterns[64386] = 29'b1_111101110000_010_1_111011100001;
      patterns[64387] = 29'b1_111101110000_011_1_110111000011;
      patterns[64388] = 29'b1_111101110000_100_0_111110111000;
      patterns[64389] = 29'b1_111101110000_101_0_011111011100;
      patterns[64390] = 29'b1_111101110000_110_1_111101110000;
      patterns[64391] = 29'b1_111101110000_111_1_111101110000;
      patterns[64392] = 29'b1_111101110001_000_1_111101110001;
      patterns[64393] = 29'b1_111101110001_001_1_110001111101;
      patterns[64394] = 29'b1_111101110001_010_1_111011100011;
      patterns[64395] = 29'b1_111101110001_011_1_110111000111;
      patterns[64396] = 29'b1_111101110001_100_1_111110111000;
      patterns[64397] = 29'b1_111101110001_101_0_111111011100;
      patterns[64398] = 29'b1_111101110001_110_1_111101110001;
      patterns[64399] = 29'b1_111101110001_111_1_111101110001;
      patterns[64400] = 29'b1_111101110010_000_1_111101110010;
      patterns[64401] = 29'b1_111101110010_001_1_110010111101;
      patterns[64402] = 29'b1_111101110010_010_1_111011100101;
      patterns[64403] = 29'b1_111101110010_011_1_110111001011;
      patterns[64404] = 29'b1_111101110010_100_0_111110111001;
      patterns[64405] = 29'b1_111101110010_101_1_011111011100;
      patterns[64406] = 29'b1_111101110010_110_1_111101110010;
      patterns[64407] = 29'b1_111101110010_111_1_111101110010;
      patterns[64408] = 29'b1_111101110011_000_1_111101110011;
      patterns[64409] = 29'b1_111101110011_001_1_110011111101;
      patterns[64410] = 29'b1_111101110011_010_1_111011100111;
      patterns[64411] = 29'b1_111101110011_011_1_110111001111;
      patterns[64412] = 29'b1_111101110011_100_1_111110111001;
      patterns[64413] = 29'b1_111101110011_101_1_111111011100;
      patterns[64414] = 29'b1_111101110011_110_1_111101110011;
      patterns[64415] = 29'b1_111101110011_111_1_111101110011;
      patterns[64416] = 29'b1_111101110100_000_1_111101110100;
      patterns[64417] = 29'b1_111101110100_001_1_110100111101;
      patterns[64418] = 29'b1_111101110100_010_1_111011101001;
      patterns[64419] = 29'b1_111101110100_011_1_110111010011;
      patterns[64420] = 29'b1_111101110100_100_0_111110111010;
      patterns[64421] = 29'b1_111101110100_101_0_011111011101;
      patterns[64422] = 29'b1_111101110100_110_1_111101110100;
      patterns[64423] = 29'b1_111101110100_111_1_111101110100;
      patterns[64424] = 29'b1_111101110101_000_1_111101110101;
      patterns[64425] = 29'b1_111101110101_001_1_110101111101;
      patterns[64426] = 29'b1_111101110101_010_1_111011101011;
      patterns[64427] = 29'b1_111101110101_011_1_110111010111;
      patterns[64428] = 29'b1_111101110101_100_1_111110111010;
      patterns[64429] = 29'b1_111101110101_101_0_111111011101;
      patterns[64430] = 29'b1_111101110101_110_1_111101110101;
      patterns[64431] = 29'b1_111101110101_111_1_111101110101;
      patterns[64432] = 29'b1_111101110110_000_1_111101110110;
      patterns[64433] = 29'b1_111101110110_001_1_110110111101;
      patterns[64434] = 29'b1_111101110110_010_1_111011101101;
      patterns[64435] = 29'b1_111101110110_011_1_110111011011;
      patterns[64436] = 29'b1_111101110110_100_0_111110111011;
      patterns[64437] = 29'b1_111101110110_101_1_011111011101;
      patterns[64438] = 29'b1_111101110110_110_1_111101110110;
      patterns[64439] = 29'b1_111101110110_111_1_111101110110;
      patterns[64440] = 29'b1_111101110111_000_1_111101110111;
      patterns[64441] = 29'b1_111101110111_001_1_110111111101;
      patterns[64442] = 29'b1_111101110111_010_1_111011101111;
      patterns[64443] = 29'b1_111101110111_011_1_110111011111;
      patterns[64444] = 29'b1_111101110111_100_1_111110111011;
      patterns[64445] = 29'b1_111101110111_101_1_111111011101;
      patterns[64446] = 29'b1_111101110111_110_1_111101110111;
      patterns[64447] = 29'b1_111101110111_111_1_111101110111;
      patterns[64448] = 29'b1_111101111000_000_1_111101111000;
      patterns[64449] = 29'b1_111101111000_001_1_111000111101;
      patterns[64450] = 29'b1_111101111000_010_1_111011110001;
      patterns[64451] = 29'b1_111101111000_011_1_110111100011;
      patterns[64452] = 29'b1_111101111000_100_0_111110111100;
      patterns[64453] = 29'b1_111101111000_101_0_011111011110;
      patterns[64454] = 29'b1_111101111000_110_1_111101111000;
      patterns[64455] = 29'b1_111101111000_111_1_111101111000;
      patterns[64456] = 29'b1_111101111001_000_1_111101111001;
      patterns[64457] = 29'b1_111101111001_001_1_111001111101;
      patterns[64458] = 29'b1_111101111001_010_1_111011110011;
      patterns[64459] = 29'b1_111101111001_011_1_110111100111;
      patterns[64460] = 29'b1_111101111001_100_1_111110111100;
      patterns[64461] = 29'b1_111101111001_101_0_111111011110;
      patterns[64462] = 29'b1_111101111001_110_1_111101111001;
      patterns[64463] = 29'b1_111101111001_111_1_111101111001;
      patterns[64464] = 29'b1_111101111010_000_1_111101111010;
      patterns[64465] = 29'b1_111101111010_001_1_111010111101;
      patterns[64466] = 29'b1_111101111010_010_1_111011110101;
      patterns[64467] = 29'b1_111101111010_011_1_110111101011;
      patterns[64468] = 29'b1_111101111010_100_0_111110111101;
      patterns[64469] = 29'b1_111101111010_101_1_011111011110;
      patterns[64470] = 29'b1_111101111010_110_1_111101111010;
      patterns[64471] = 29'b1_111101111010_111_1_111101111010;
      patterns[64472] = 29'b1_111101111011_000_1_111101111011;
      patterns[64473] = 29'b1_111101111011_001_1_111011111101;
      patterns[64474] = 29'b1_111101111011_010_1_111011110111;
      patterns[64475] = 29'b1_111101111011_011_1_110111101111;
      patterns[64476] = 29'b1_111101111011_100_1_111110111101;
      patterns[64477] = 29'b1_111101111011_101_1_111111011110;
      patterns[64478] = 29'b1_111101111011_110_1_111101111011;
      patterns[64479] = 29'b1_111101111011_111_1_111101111011;
      patterns[64480] = 29'b1_111101111100_000_1_111101111100;
      patterns[64481] = 29'b1_111101111100_001_1_111100111101;
      patterns[64482] = 29'b1_111101111100_010_1_111011111001;
      patterns[64483] = 29'b1_111101111100_011_1_110111110011;
      patterns[64484] = 29'b1_111101111100_100_0_111110111110;
      patterns[64485] = 29'b1_111101111100_101_0_011111011111;
      patterns[64486] = 29'b1_111101111100_110_1_111101111100;
      patterns[64487] = 29'b1_111101111100_111_1_111101111100;
      patterns[64488] = 29'b1_111101111101_000_1_111101111101;
      patterns[64489] = 29'b1_111101111101_001_1_111101111101;
      patterns[64490] = 29'b1_111101111101_010_1_111011111011;
      patterns[64491] = 29'b1_111101111101_011_1_110111110111;
      patterns[64492] = 29'b1_111101111101_100_1_111110111110;
      patterns[64493] = 29'b1_111101111101_101_0_111111011111;
      patterns[64494] = 29'b1_111101111101_110_1_111101111101;
      patterns[64495] = 29'b1_111101111101_111_1_111101111101;
      patterns[64496] = 29'b1_111101111110_000_1_111101111110;
      patterns[64497] = 29'b1_111101111110_001_1_111110111101;
      patterns[64498] = 29'b1_111101111110_010_1_111011111101;
      patterns[64499] = 29'b1_111101111110_011_1_110111111011;
      patterns[64500] = 29'b1_111101111110_100_0_111110111111;
      patterns[64501] = 29'b1_111101111110_101_1_011111011111;
      patterns[64502] = 29'b1_111101111110_110_1_111101111110;
      patterns[64503] = 29'b1_111101111110_111_1_111101111110;
      patterns[64504] = 29'b1_111101111111_000_1_111101111111;
      patterns[64505] = 29'b1_111101111111_001_1_111111111101;
      patterns[64506] = 29'b1_111101111111_010_1_111011111111;
      patterns[64507] = 29'b1_111101111111_011_1_110111111111;
      patterns[64508] = 29'b1_111101111111_100_1_111110111111;
      patterns[64509] = 29'b1_111101111111_101_1_111111011111;
      patterns[64510] = 29'b1_111101111111_110_1_111101111111;
      patterns[64511] = 29'b1_111101111111_111_1_111101111111;
      patterns[64512] = 29'b1_111110000000_000_1_111110000000;
      patterns[64513] = 29'b1_111110000000_001_1_000000111110;
      patterns[64514] = 29'b1_111110000000_010_1_111100000001;
      patterns[64515] = 29'b1_111110000000_011_1_111000000011;
      patterns[64516] = 29'b1_111110000000_100_0_111111000000;
      patterns[64517] = 29'b1_111110000000_101_0_011111100000;
      patterns[64518] = 29'b1_111110000000_110_1_111110000000;
      patterns[64519] = 29'b1_111110000000_111_1_111110000000;
      patterns[64520] = 29'b1_111110000001_000_1_111110000001;
      patterns[64521] = 29'b1_111110000001_001_1_000001111110;
      patterns[64522] = 29'b1_111110000001_010_1_111100000011;
      patterns[64523] = 29'b1_111110000001_011_1_111000000111;
      patterns[64524] = 29'b1_111110000001_100_1_111111000000;
      patterns[64525] = 29'b1_111110000001_101_0_111111100000;
      patterns[64526] = 29'b1_111110000001_110_1_111110000001;
      patterns[64527] = 29'b1_111110000001_111_1_111110000001;
      patterns[64528] = 29'b1_111110000010_000_1_111110000010;
      patterns[64529] = 29'b1_111110000010_001_1_000010111110;
      patterns[64530] = 29'b1_111110000010_010_1_111100000101;
      patterns[64531] = 29'b1_111110000010_011_1_111000001011;
      patterns[64532] = 29'b1_111110000010_100_0_111111000001;
      patterns[64533] = 29'b1_111110000010_101_1_011111100000;
      patterns[64534] = 29'b1_111110000010_110_1_111110000010;
      patterns[64535] = 29'b1_111110000010_111_1_111110000010;
      patterns[64536] = 29'b1_111110000011_000_1_111110000011;
      patterns[64537] = 29'b1_111110000011_001_1_000011111110;
      patterns[64538] = 29'b1_111110000011_010_1_111100000111;
      patterns[64539] = 29'b1_111110000011_011_1_111000001111;
      patterns[64540] = 29'b1_111110000011_100_1_111111000001;
      patterns[64541] = 29'b1_111110000011_101_1_111111100000;
      patterns[64542] = 29'b1_111110000011_110_1_111110000011;
      patterns[64543] = 29'b1_111110000011_111_1_111110000011;
      patterns[64544] = 29'b1_111110000100_000_1_111110000100;
      patterns[64545] = 29'b1_111110000100_001_1_000100111110;
      patterns[64546] = 29'b1_111110000100_010_1_111100001001;
      patterns[64547] = 29'b1_111110000100_011_1_111000010011;
      patterns[64548] = 29'b1_111110000100_100_0_111111000010;
      patterns[64549] = 29'b1_111110000100_101_0_011111100001;
      patterns[64550] = 29'b1_111110000100_110_1_111110000100;
      patterns[64551] = 29'b1_111110000100_111_1_111110000100;
      patterns[64552] = 29'b1_111110000101_000_1_111110000101;
      patterns[64553] = 29'b1_111110000101_001_1_000101111110;
      patterns[64554] = 29'b1_111110000101_010_1_111100001011;
      patterns[64555] = 29'b1_111110000101_011_1_111000010111;
      patterns[64556] = 29'b1_111110000101_100_1_111111000010;
      patterns[64557] = 29'b1_111110000101_101_0_111111100001;
      patterns[64558] = 29'b1_111110000101_110_1_111110000101;
      patterns[64559] = 29'b1_111110000101_111_1_111110000101;
      patterns[64560] = 29'b1_111110000110_000_1_111110000110;
      patterns[64561] = 29'b1_111110000110_001_1_000110111110;
      patterns[64562] = 29'b1_111110000110_010_1_111100001101;
      patterns[64563] = 29'b1_111110000110_011_1_111000011011;
      patterns[64564] = 29'b1_111110000110_100_0_111111000011;
      patterns[64565] = 29'b1_111110000110_101_1_011111100001;
      patterns[64566] = 29'b1_111110000110_110_1_111110000110;
      patterns[64567] = 29'b1_111110000110_111_1_111110000110;
      patterns[64568] = 29'b1_111110000111_000_1_111110000111;
      patterns[64569] = 29'b1_111110000111_001_1_000111111110;
      patterns[64570] = 29'b1_111110000111_010_1_111100001111;
      patterns[64571] = 29'b1_111110000111_011_1_111000011111;
      patterns[64572] = 29'b1_111110000111_100_1_111111000011;
      patterns[64573] = 29'b1_111110000111_101_1_111111100001;
      patterns[64574] = 29'b1_111110000111_110_1_111110000111;
      patterns[64575] = 29'b1_111110000111_111_1_111110000111;
      patterns[64576] = 29'b1_111110001000_000_1_111110001000;
      patterns[64577] = 29'b1_111110001000_001_1_001000111110;
      patterns[64578] = 29'b1_111110001000_010_1_111100010001;
      patterns[64579] = 29'b1_111110001000_011_1_111000100011;
      patterns[64580] = 29'b1_111110001000_100_0_111111000100;
      patterns[64581] = 29'b1_111110001000_101_0_011111100010;
      patterns[64582] = 29'b1_111110001000_110_1_111110001000;
      patterns[64583] = 29'b1_111110001000_111_1_111110001000;
      patterns[64584] = 29'b1_111110001001_000_1_111110001001;
      patterns[64585] = 29'b1_111110001001_001_1_001001111110;
      patterns[64586] = 29'b1_111110001001_010_1_111100010011;
      patterns[64587] = 29'b1_111110001001_011_1_111000100111;
      patterns[64588] = 29'b1_111110001001_100_1_111111000100;
      patterns[64589] = 29'b1_111110001001_101_0_111111100010;
      patterns[64590] = 29'b1_111110001001_110_1_111110001001;
      patterns[64591] = 29'b1_111110001001_111_1_111110001001;
      patterns[64592] = 29'b1_111110001010_000_1_111110001010;
      patterns[64593] = 29'b1_111110001010_001_1_001010111110;
      patterns[64594] = 29'b1_111110001010_010_1_111100010101;
      patterns[64595] = 29'b1_111110001010_011_1_111000101011;
      patterns[64596] = 29'b1_111110001010_100_0_111111000101;
      patterns[64597] = 29'b1_111110001010_101_1_011111100010;
      patterns[64598] = 29'b1_111110001010_110_1_111110001010;
      patterns[64599] = 29'b1_111110001010_111_1_111110001010;
      patterns[64600] = 29'b1_111110001011_000_1_111110001011;
      patterns[64601] = 29'b1_111110001011_001_1_001011111110;
      patterns[64602] = 29'b1_111110001011_010_1_111100010111;
      patterns[64603] = 29'b1_111110001011_011_1_111000101111;
      patterns[64604] = 29'b1_111110001011_100_1_111111000101;
      patterns[64605] = 29'b1_111110001011_101_1_111111100010;
      patterns[64606] = 29'b1_111110001011_110_1_111110001011;
      patterns[64607] = 29'b1_111110001011_111_1_111110001011;
      patterns[64608] = 29'b1_111110001100_000_1_111110001100;
      patterns[64609] = 29'b1_111110001100_001_1_001100111110;
      patterns[64610] = 29'b1_111110001100_010_1_111100011001;
      patterns[64611] = 29'b1_111110001100_011_1_111000110011;
      patterns[64612] = 29'b1_111110001100_100_0_111111000110;
      patterns[64613] = 29'b1_111110001100_101_0_011111100011;
      patterns[64614] = 29'b1_111110001100_110_1_111110001100;
      patterns[64615] = 29'b1_111110001100_111_1_111110001100;
      patterns[64616] = 29'b1_111110001101_000_1_111110001101;
      patterns[64617] = 29'b1_111110001101_001_1_001101111110;
      patterns[64618] = 29'b1_111110001101_010_1_111100011011;
      patterns[64619] = 29'b1_111110001101_011_1_111000110111;
      patterns[64620] = 29'b1_111110001101_100_1_111111000110;
      patterns[64621] = 29'b1_111110001101_101_0_111111100011;
      patterns[64622] = 29'b1_111110001101_110_1_111110001101;
      patterns[64623] = 29'b1_111110001101_111_1_111110001101;
      patterns[64624] = 29'b1_111110001110_000_1_111110001110;
      patterns[64625] = 29'b1_111110001110_001_1_001110111110;
      patterns[64626] = 29'b1_111110001110_010_1_111100011101;
      patterns[64627] = 29'b1_111110001110_011_1_111000111011;
      patterns[64628] = 29'b1_111110001110_100_0_111111000111;
      patterns[64629] = 29'b1_111110001110_101_1_011111100011;
      patterns[64630] = 29'b1_111110001110_110_1_111110001110;
      patterns[64631] = 29'b1_111110001110_111_1_111110001110;
      patterns[64632] = 29'b1_111110001111_000_1_111110001111;
      patterns[64633] = 29'b1_111110001111_001_1_001111111110;
      patterns[64634] = 29'b1_111110001111_010_1_111100011111;
      patterns[64635] = 29'b1_111110001111_011_1_111000111111;
      patterns[64636] = 29'b1_111110001111_100_1_111111000111;
      patterns[64637] = 29'b1_111110001111_101_1_111111100011;
      patterns[64638] = 29'b1_111110001111_110_1_111110001111;
      patterns[64639] = 29'b1_111110001111_111_1_111110001111;
      patterns[64640] = 29'b1_111110010000_000_1_111110010000;
      patterns[64641] = 29'b1_111110010000_001_1_010000111110;
      patterns[64642] = 29'b1_111110010000_010_1_111100100001;
      patterns[64643] = 29'b1_111110010000_011_1_111001000011;
      patterns[64644] = 29'b1_111110010000_100_0_111111001000;
      patterns[64645] = 29'b1_111110010000_101_0_011111100100;
      patterns[64646] = 29'b1_111110010000_110_1_111110010000;
      patterns[64647] = 29'b1_111110010000_111_1_111110010000;
      patterns[64648] = 29'b1_111110010001_000_1_111110010001;
      patterns[64649] = 29'b1_111110010001_001_1_010001111110;
      patterns[64650] = 29'b1_111110010001_010_1_111100100011;
      patterns[64651] = 29'b1_111110010001_011_1_111001000111;
      patterns[64652] = 29'b1_111110010001_100_1_111111001000;
      patterns[64653] = 29'b1_111110010001_101_0_111111100100;
      patterns[64654] = 29'b1_111110010001_110_1_111110010001;
      patterns[64655] = 29'b1_111110010001_111_1_111110010001;
      patterns[64656] = 29'b1_111110010010_000_1_111110010010;
      patterns[64657] = 29'b1_111110010010_001_1_010010111110;
      patterns[64658] = 29'b1_111110010010_010_1_111100100101;
      patterns[64659] = 29'b1_111110010010_011_1_111001001011;
      patterns[64660] = 29'b1_111110010010_100_0_111111001001;
      patterns[64661] = 29'b1_111110010010_101_1_011111100100;
      patterns[64662] = 29'b1_111110010010_110_1_111110010010;
      patterns[64663] = 29'b1_111110010010_111_1_111110010010;
      patterns[64664] = 29'b1_111110010011_000_1_111110010011;
      patterns[64665] = 29'b1_111110010011_001_1_010011111110;
      patterns[64666] = 29'b1_111110010011_010_1_111100100111;
      patterns[64667] = 29'b1_111110010011_011_1_111001001111;
      patterns[64668] = 29'b1_111110010011_100_1_111111001001;
      patterns[64669] = 29'b1_111110010011_101_1_111111100100;
      patterns[64670] = 29'b1_111110010011_110_1_111110010011;
      patterns[64671] = 29'b1_111110010011_111_1_111110010011;
      patterns[64672] = 29'b1_111110010100_000_1_111110010100;
      patterns[64673] = 29'b1_111110010100_001_1_010100111110;
      patterns[64674] = 29'b1_111110010100_010_1_111100101001;
      patterns[64675] = 29'b1_111110010100_011_1_111001010011;
      patterns[64676] = 29'b1_111110010100_100_0_111111001010;
      patterns[64677] = 29'b1_111110010100_101_0_011111100101;
      patterns[64678] = 29'b1_111110010100_110_1_111110010100;
      patterns[64679] = 29'b1_111110010100_111_1_111110010100;
      patterns[64680] = 29'b1_111110010101_000_1_111110010101;
      patterns[64681] = 29'b1_111110010101_001_1_010101111110;
      patterns[64682] = 29'b1_111110010101_010_1_111100101011;
      patterns[64683] = 29'b1_111110010101_011_1_111001010111;
      patterns[64684] = 29'b1_111110010101_100_1_111111001010;
      patterns[64685] = 29'b1_111110010101_101_0_111111100101;
      patterns[64686] = 29'b1_111110010101_110_1_111110010101;
      patterns[64687] = 29'b1_111110010101_111_1_111110010101;
      patterns[64688] = 29'b1_111110010110_000_1_111110010110;
      patterns[64689] = 29'b1_111110010110_001_1_010110111110;
      patterns[64690] = 29'b1_111110010110_010_1_111100101101;
      patterns[64691] = 29'b1_111110010110_011_1_111001011011;
      patterns[64692] = 29'b1_111110010110_100_0_111111001011;
      patterns[64693] = 29'b1_111110010110_101_1_011111100101;
      patterns[64694] = 29'b1_111110010110_110_1_111110010110;
      patterns[64695] = 29'b1_111110010110_111_1_111110010110;
      patterns[64696] = 29'b1_111110010111_000_1_111110010111;
      patterns[64697] = 29'b1_111110010111_001_1_010111111110;
      patterns[64698] = 29'b1_111110010111_010_1_111100101111;
      patterns[64699] = 29'b1_111110010111_011_1_111001011111;
      patterns[64700] = 29'b1_111110010111_100_1_111111001011;
      patterns[64701] = 29'b1_111110010111_101_1_111111100101;
      patterns[64702] = 29'b1_111110010111_110_1_111110010111;
      patterns[64703] = 29'b1_111110010111_111_1_111110010111;
      patterns[64704] = 29'b1_111110011000_000_1_111110011000;
      patterns[64705] = 29'b1_111110011000_001_1_011000111110;
      patterns[64706] = 29'b1_111110011000_010_1_111100110001;
      patterns[64707] = 29'b1_111110011000_011_1_111001100011;
      patterns[64708] = 29'b1_111110011000_100_0_111111001100;
      patterns[64709] = 29'b1_111110011000_101_0_011111100110;
      patterns[64710] = 29'b1_111110011000_110_1_111110011000;
      patterns[64711] = 29'b1_111110011000_111_1_111110011000;
      patterns[64712] = 29'b1_111110011001_000_1_111110011001;
      patterns[64713] = 29'b1_111110011001_001_1_011001111110;
      patterns[64714] = 29'b1_111110011001_010_1_111100110011;
      patterns[64715] = 29'b1_111110011001_011_1_111001100111;
      patterns[64716] = 29'b1_111110011001_100_1_111111001100;
      patterns[64717] = 29'b1_111110011001_101_0_111111100110;
      patterns[64718] = 29'b1_111110011001_110_1_111110011001;
      patterns[64719] = 29'b1_111110011001_111_1_111110011001;
      patterns[64720] = 29'b1_111110011010_000_1_111110011010;
      patterns[64721] = 29'b1_111110011010_001_1_011010111110;
      patterns[64722] = 29'b1_111110011010_010_1_111100110101;
      patterns[64723] = 29'b1_111110011010_011_1_111001101011;
      patterns[64724] = 29'b1_111110011010_100_0_111111001101;
      patterns[64725] = 29'b1_111110011010_101_1_011111100110;
      patterns[64726] = 29'b1_111110011010_110_1_111110011010;
      patterns[64727] = 29'b1_111110011010_111_1_111110011010;
      patterns[64728] = 29'b1_111110011011_000_1_111110011011;
      patterns[64729] = 29'b1_111110011011_001_1_011011111110;
      patterns[64730] = 29'b1_111110011011_010_1_111100110111;
      patterns[64731] = 29'b1_111110011011_011_1_111001101111;
      patterns[64732] = 29'b1_111110011011_100_1_111111001101;
      patterns[64733] = 29'b1_111110011011_101_1_111111100110;
      patterns[64734] = 29'b1_111110011011_110_1_111110011011;
      patterns[64735] = 29'b1_111110011011_111_1_111110011011;
      patterns[64736] = 29'b1_111110011100_000_1_111110011100;
      patterns[64737] = 29'b1_111110011100_001_1_011100111110;
      patterns[64738] = 29'b1_111110011100_010_1_111100111001;
      patterns[64739] = 29'b1_111110011100_011_1_111001110011;
      patterns[64740] = 29'b1_111110011100_100_0_111111001110;
      patterns[64741] = 29'b1_111110011100_101_0_011111100111;
      patterns[64742] = 29'b1_111110011100_110_1_111110011100;
      patterns[64743] = 29'b1_111110011100_111_1_111110011100;
      patterns[64744] = 29'b1_111110011101_000_1_111110011101;
      patterns[64745] = 29'b1_111110011101_001_1_011101111110;
      patterns[64746] = 29'b1_111110011101_010_1_111100111011;
      patterns[64747] = 29'b1_111110011101_011_1_111001110111;
      patterns[64748] = 29'b1_111110011101_100_1_111111001110;
      patterns[64749] = 29'b1_111110011101_101_0_111111100111;
      patterns[64750] = 29'b1_111110011101_110_1_111110011101;
      patterns[64751] = 29'b1_111110011101_111_1_111110011101;
      patterns[64752] = 29'b1_111110011110_000_1_111110011110;
      patterns[64753] = 29'b1_111110011110_001_1_011110111110;
      patterns[64754] = 29'b1_111110011110_010_1_111100111101;
      patterns[64755] = 29'b1_111110011110_011_1_111001111011;
      patterns[64756] = 29'b1_111110011110_100_0_111111001111;
      patterns[64757] = 29'b1_111110011110_101_1_011111100111;
      patterns[64758] = 29'b1_111110011110_110_1_111110011110;
      patterns[64759] = 29'b1_111110011110_111_1_111110011110;
      patterns[64760] = 29'b1_111110011111_000_1_111110011111;
      patterns[64761] = 29'b1_111110011111_001_1_011111111110;
      patterns[64762] = 29'b1_111110011111_010_1_111100111111;
      patterns[64763] = 29'b1_111110011111_011_1_111001111111;
      patterns[64764] = 29'b1_111110011111_100_1_111111001111;
      patterns[64765] = 29'b1_111110011111_101_1_111111100111;
      patterns[64766] = 29'b1_111110011111_110_1_111110011111;
      patterns[64767] = 29'b1_111110011111_111_1_111110011111;
      patterns[64768] = 29'b1_111110100000_000_1_111110100000;
      patterns[64769] = 29'b1_111110100000_001_1_100000111110;
      patterns[64770] = 29'b1_111110100000_010_1_111101000001;
      patterns[64771] = 29'b1_111110100000_011_1_111010000011;
      patterns[64772] = 29'b1_111110100000_100_0_111111010000;
      patterns[64773] = 29'b1_111110100000_101_0_011111101000;
      patterns[64774] = 29'b1_111110100000_110_1_111110100000;
      patterns[64775] = 29'b1_111110100000_111_1_111110100000;
      patterns[64776] = 29'b1_111110100001_000_1_111110100001;
      patterns[64777] = 29'b1_111110100001_001_1_100001111110;
      patterns[64778] = 29'b1_111110100001_010_1_111101000011;
      patterns[64779] = 29'b1_111110100001_011_1_111010000111;
      patterns[64780] = 29'b1_111110100001_100_1_111111010000;
      patterns[64781] = 29'b1_111110100001_101_0_111111101000;
      patterns[64782] = 29'b1_111110100001_110_1_111110100001;
      patterns[64783] = 29'b1_111110100001_111_1_111110100001;
      patterns[64784] = 29'b1_111110100010_000_1_111110100010;
      patterns[64785] = 29'b1_111110100010_001_1_100010111110;
      patterns[64786] = 29'b1_111110100010_010_1_111101000101;
      patterns[64787] = 29'b1_111110100010_011_1_111010001011;
      patterns[64788] = 29'b1_111110100010_100_0_111111010001;
      patterns[64789] = 29'b1_111110100010_101_1_011111101000;
      patterns[64790] = 29'b1_111110100010_110_1_111110100010;
      patterns[64791] = 29'b1_111110100010_111_1_111110100010;
      patterns[64792] = 29'b1_111110100011_000_1_111110100011;
      patterns[64793] = 29'b1_111110100011_001_1_100011111110;
      patterns[64794] = 29'b1_111110100011_010_1_111101000111;
      patterns[64795] = 29'b1_111110100011_011_1_111010001111;
      patterns[64796] = 29'b1_111110100011_100_1_111111010001;
      patterns[64797] = 29'b1_111110100011_101_1_111111101000;
      patterns[64798] = 29'b1_111110100011_110_1_111110100011;
      patterns[64799] = 29'b1_111110100011_111_1_111110100011;
      patterns[64800] = 29'b1_111110100100_000_1_111110100100;
      patterns[64801] = 29'b1_111110100100_001_1_100100111110;
      patterns[64802] = 29'b1_111110100100_010_1_111101001001;
      patterns[64803] = 29'b1_111110100100_011_1_111010010011;
      patterns[64804] = 29'b1_111110100100_100_0_111111010010;
      patterns[64805] = 29'b1_111110100100_101_0_011111101001;
      patterns[64806] = 29'b1_111110100100_110_1_111110100100;
      patterns[64807] = 29'b1_111110100100_111_1_111110100100;
      patterns[64808] = 29'b1_111110100101_000_1_111110100101;
      patterns[64809] = 29'b1_111110100101_001_1_100101111110;
      patterns[64810] = 29'b1_111110100101_010_1_111101001011;
      patterns[64811] = 29'b1_111110100101_011_1_111010010111;
      patterns[64812] = 29'b1_111110100101_100_1_111111010010;
      patterns[64813] = 29'b1_111110100101_101_0_111111101001;
      patterns[64814] = 29'b1_111110100101_110_1_111110100101;
      patterns[64815] = 29'b1_111110100101_111_1_111110100101;
      patterns[64816] = 29'b1_111110100110_000_1_111110100110;
      patterns[64817] = 29'b1_111110100110_001_1_100110111110;
      patterns[64818] = 29'b1_111110100110_010_1_111101001101;
      patterns[64819] = 29'b1_111110100110_011_1_111010011011;
      patterns[64820] = 29'b1_111110100110_100_0_111111010011;
      patterns[64821] = 29'b1_111110100110_101_1_011111101001;
      patterns[64822] = 29'b1_111110100110_110_1_111110100110;
      patterns[64823] = 29'b1_111110100110_111_1_111110100110;
      patterns[64824] = 29'b1_111110100111_000_1_111110100111;
      patterns[64825] = 29'b1_111110100111_001_1_100111111110;
      patterns[64826] = 29'b1_111110100111_010_1_111101001111;
      patterns[64827] = 29'b1_111110100111_011_1_111010011111;
      patterns[64828] = 29'b1_111110100111_100_1_111111010011;
      patterns[64829] = 29'b1_111110100111_101_1_111111101001;
      patterns[64830] = 29'b1_111110100111_110_1_111110100111;
      patterns[64831] = 29'b1_111110100111_111_1_111110100111;
      patterns[64832] = 29'b1_111110101000_000_1_111110101000;
      patterns[64833] = 29'b1_111110101000_001_1_101000111110;
      patterns[64834] = 29'b1_111110101000_010_1_111101010001;
      patterns[64835] = 29'b1_111110101000_011_1_111010100011;
      patterns[64836] = 29'b1_111110101000_100_0_111111010100;
      patterns[64837] = 29'b1_111110101000_101_0_011111101010;
      patterns[64838] = 29'b1_111110101000_110_1_111110101000;
      patterns[64839] = 29'b1_111110101000_111_1_111110101000;
      patterns[64840] = 29'b1_111110101001_000_1_111110101001;
      patterns[64841] = 29'b1_111110101001_001_1_101001111110;
      patterns[64842] = 29'b1_111110101001_010_1_111101010011;
      patterns[64843] = 29'b1_111110101001_011_1_111010100111;
      patterns[64844] = 29'b1_111110101001_100_1_111111010100;
      patterns[64845] = 29'b1_111110101001_101_0_111111101010;
      patterns[64846] = 29'b1_111110101001_110_1_111110101001;
      patterns[64847] = 29'b1_111110101001_111_1_111110101001;
      patterns[64848] = 29'b1_111110101010_000_1_111110101010;
      patterns[64849] = 29'b1_111110101010_001_1_101010111110;
      patterns[64850] = 29'b1_111110101010_010_1_111101010101;
      patterns[64851] = 29'b1_111110101010_011_1_111010101011;
      patterns[64852] = 29'b1_111110101010_100_0_111111010101;
      patterns[64853] = 29'b1_111110101010_101_1_011111101010;
      patterns[64854] = 29'b1_111110101010_110_1_111110101010;
      patterns[64855] = 29'b1_111110101010_111_1_111110101010;
      patterns[64856] = 29'b1_111110101011_000_1_111110101011;
      patterns[64857] = 29'b1_111110101011_001_1_101011111110;
      patterns[64858] = 29'b1_111110101011_010_1_111101010111;
      patterns[64859] = 29'b1_111110101011_011_1_111010101111;
      patterns[64860] = 29'b1_111110101011_100_1_111111010101;
      patterns[64861] = 29'b1_111110101011_101_1_111111101010;
      patterns[64862] = 29'b1_111110101011_110_1_111110101011;
      patterns[64863] = 29'b1_111110101011_111_1_111110101011;
      patterns[64864] = 29'b1_111110101100_000_1_111110101100;
      patterns[64865] = 29'b1_111110101100_001_1_101100111110;
      patterns[64866] = 29'b1_111110101100_010_1_111101011001;
      patterns[64867] = 29'b1_111110101100_011_1_111010110011;
      patterns[64868] = 29'b1_111110101100_100_0_111111010110;
      patterns[64869] = 29'b1_111110101100_101_0_011111101011;
      patterns[64870] = 29'b1_111110101100_110_1_111110101100;
      patterns[64871] = 29'b1_111110101100_111_1_111110101100;
      patterns[64872] = 29'b1_111110101101_000_1_111110101101;
      patterns[64873] = 29'b1_111110101101_001_1_101101111110;
      patterns[64874] = 29'b1_111110101101_010_1_111101011011;
      patterns[64875] = 29'b1_111110101101_011_1_111010110111;
      patterns[64876] = 29'b1_111110101101_100_1_111111010110;
      patterns[64877] = 29'b1_111110101101_101_0_111111101011;
      patterns[64878] = 29'b1_111110101101_110_1_111110101101;
      patterns[64879] = 29'b1_111110101101_111_1_111110101101;
      patterns[64880] = 29'b1_111110101110_000_1_111110101110;
      patterns[64881] = 29'b1_111110101110_001_1_101110111110;
      patterns[64882] = 29'b1_111110101110_010_1_111101011101;
      patterns[64883] = 29'b1_111110101110_011_1_111010111011;
      patterns[64884] = 29'b1_111110101110_100_0_111111010111;
      patterns[64885] = 29'b1_111110101110_101_1_011111101011;
      patterns[64886] = 29'b1_111110101110_110_1_111110101110;
      patterns[64887] = 29'b1_111110101110_111_1_111110101110;
      patterns[64888] = 29'b1_111110101111_000_1_111110101111;
      patterns[64889] = 29'b1_111110101111_001_1_101111111110;
      patterns[64890] = 29'b1_111110101111_010_1_111101011111;
      patterns[64891] = 29'b1_111110101111_011_1_111010111111;
      patterns[64892] = 29'b1_111110101111_100_1_111111010111;
      patterns[64893] = 29'b1_111110101111_101_1_111111101011;
      patterns[64894] = 29'b1_111110101111_110_1_111110101111;
      patterns[64895] = 29'b1_111110101111_111_1_111110101111;
      patterns[64896] = 29'b1_111110110000_000_1_111110110000;
      patterns[64897] = 29'b1_111110110000_001_1_110000111110;
      patterns[64898] = 29'b1_111110110000_010_1_111101100001;
      patterns[64899] = 29'b1_111110110000_011_1_111011000011;
      patterns[64900] = 29'b1_111110110000_100_0_111111011000;
      patterns[64901] = 29'b1_111110110000_101_0_011111101100;
      patterns[64902] = 29'b1_111110110000_110_1_111110110000;
      patterns[64903] = 29'b1_111110110000_111_1_111110110000;
      patterns[64904] = 29'b1_111110110001_000_1_111110110001;
      patterns[64905] = 29'b1_111110110001_001_1_110001111110;
      patterns[64906] = 29'b1_111110110001_010_1_111101100011;
      patterns[64907] = 29'b1_111110110001_011_1_111011000111;
      patterns[64908] = 29'b1_111110110001_100_1_111111011000;
      patterns[64909] = 29'b1_111110110001_101_0_111111101100;
      patterns[64910] = 29'b1_111110110001_110_1_111110110001;
      patterns[64911] = 29'b1_111110110001_111_1_111110110001;
      patterns[64912] = 29'b1_111110110010_000_1_111110110010;
      patterns[64913] = 29'b1_111110110010_001_1_110010111110;
      patterns[64914] = 29'b1_111110110010_010_1_111101100101;
      patterns[64915] = 29'b1_111110110010_011_1_111011001011;
      patterns[64916] = 29'b1_111110110010_100_0_111111011001;
      patterns[64917] = 29'b1_111110110010_101_1_011111101100;
      patterns[64918] = 29'b1_111110110010_110_1_111110110010;
      patterns[64919] = 29'b1_111110110010_111_1_111110110010;
      patterns[64920] = 29'b1_111110110011_000_1_111110110011;
      patterns[64921] = 29'b1_111110110011_001_1_110011111110;
      patterns[64922] = 29'b1_111110110011_010_1_111101100111;
      patterns[64923] = 29'b1_111110110011_011_1_111011001111;
      patterns[64924] = 29'b1_111110110011_100_1_111111011001;
      patterns[64925] = 29'b1_111110110011_101_1_111111101100;
      patterns[64926] = 29'b1_111110110011_110_1_111110110011;
      patterns[64927] = 29'b1_111110110011_111_1_111110110011;
      patterns[64928] = 29'b1_111110110100_000_1_111110110100;
      patterns[64929] = 29'b1_111110110100_001_1_110100111110;
      patterns[64930] = 29'b1_111110110100_010_1_111101101001;
      patterns[64931] = 29'b1_111110110100_011_1_111011010011;
      patterns[64932] = 29'b1_111110110100_100_0_111111011010;
      patterns[64933] = 29'b1_111110110100_101_0_011111101101;
      patterns[64934] = 29'b1_111110110100_110_1_111110110100;
      patterns[64935] = 29'b1_111110110100_111_1_111110110100;
      patterns[64936] = 29'b1_111110110101_000_1_111110110101;
      patterns[64937] = 29'b1_111110110101_001_1_110101111110;
      patterns[64938] = 29'b1_111110110101_010_1_111101101011;
      patterns[64939] = 29'b1_111110110101_011_1_111011010111;
      patterns[64940] = 29'b1_111110110101_100_1_111111011010;
      patterns[64941] = 29'b1_111110110101_101_0_111111101101;
      patterns[64942] = 29'b1_111110110101_110_1_111110110101;
      patterns[64943] = 29'b1_111110110101_111_1_111110110101;
      patterns[64944] = 29'b1_111110110110_000_1_111110110110;
      patterns[64945] = 29'b1_111110110110_001_1_110110111110;
      patterns[64946] = 29'b1_111110110110_010_1_111101101101;
      patterns[64947] = 29'b1_111110110110_011_1_111011011011;
      patterns[64948] = 29'b1_111110110110_100_0_111111011011;
      patterns[64949] = 29'b1_111110110110_101_1_011111101101;
      patterns[64950] = 29'b1_111110110110_110_1_111110110110;
      patterns[64951] = 29'b1_111110110110_111_1_111110110110;
      patterns[64952] = 29'b1_111110110111_000_1_111110110111;
      patterns[64953] = 29'b1_111110110111_001_1_110111111110;
      patterns[64954] = 29'b1_111110110111_010_1_111101101111;
      patterns[64955] = 29'b1_111110110111_011_1_111011011111;
      patterns[64956] = 29'b1_111110110111_100_1_111111011011;
      patterns[64957] = 29'b1_111110110111_101_1_111111101101;
      patterns[64958] = 29'b1_111110110111_110_1_111110110111;
      patterns[64959] = 29'b1_111110110111_111_1_111110110111;
      patterns[64960] = 29'b1_111110111000_000_1_111110111000;
      patterns[64961] = 29'b1_111110111000_001_1_111000111110;
      patterns[64962] = 29'b1_111110111000_010_1_111101110001;
      patterns[64963] = 29'b1_111110111000_011_1_111011100011;
      patterns[64964] = 29'b1_111110111000_100_0_111111011100;
      patterns[64965] = 29'b1_111110111000_101_0_011111101110;
      patterns[64966] = 29'b1_111110111000_110_1_111110111000;
      patterns[64967] = 29'b1_111110111000_111_1_111110111000;
      patterns[64968] = 29'b1_111110111001_000_1_111110111001;
      patterns[64969] = 29'b1_111110111001_001_1_111001111110;
      patterns[64970] = 29'b1_111110111001_010_1_111101110011;
      patterns[64971] = 29'b1_111110111001_011_1_111011100111;
      patterns[64972] = 29'b1_111110111001_100_1_111111011100;
      patterns[64973] = 29'b1_111110111001_101_0_111111101110;
      patterns[64974] = 29'b1_111110111001_110_1_111110111001;
      patterns[64975] = 29'b1_111110111001_111_1_111110111001;
      patterns[64976] = 29'b1_111110111010_000_1_111110111010;
      patterns[64977] = 29'b1_111110111010_001_1_111010111110;
      patterns[64978] = 29'b1_111110111010_010_1_111101110101;
      patterns[64979] = 29'b1_111110111010_011_1_111011101011;
      patterns[64980] = 29'b1_111110111010_100_0_111111011101;
      patterns[64981] = 29'b1_111110111010_101_1_011111101110;
      patterns[64982] = 29'b1_111110111010_110_1_111110111010;
      patterns[64983] = 29'b1_111110111010_111_1_111110111010;
      patterns[64984] = 29'b1_111110111011_000_1_111110111011;
      patterns[64985] = 29'b1_111110111011_001_1_111011111110;
      patterns[64986] = 29'b1_111110111011_010_1_111101110111;
      patterns[64987] = 29'b1_111110111011_011_1_111011101111;
      patterns[64988] = 29'b1_111110111011_100_1_111111011101;
      patterns[64989] = 29'b1_111110111011_101_1_111111101110;
      patterns[64990] = 29'b1_111110111011_110_1_111110111011;
      patterns[64991] = 29'b1_111110111011_111_1_111110111011;
      patterns[64992] = 29'b1_111110111100_000_1_111110111100;
      patterns[64993] = 29'b1_111110111100_001_1_111100111110;
      patterns[64994] = 29'b1_111110111100_010_1_111101111001;
      patterns[64995] = 29'b1_111110111100_011_1_111011110011;
      patterns[64996] = 29'b1_111110111100_100_0_111111011110;
      patterns[64997] = 29'b1_111110111100_101_0_011111101111;
      patterns[64998] = 29'b1_111110111100_110_1_111110111100;
      patterns[64999] = 29'b1_111110111100_111_1_111110111100;
      patterns[65000] = 29'b1_111110111101_000_1_111110111101;
      patterns[65001] = 29'b1_111110111101_001_1_111101111110;
      patterns[65002] = 29'b1_111110111101_010_1_111101111011;
      patterns[65003] = 29'b1_111110111101_011_1_111011110111;
      patterns[65004] = 29'b1_111110111101_100_1_111111011110;
      patterns[65005] = 29'b1_111110111101_101_0_111111101111;
      patterns[65006] = 29'b1_111110111101_110_1_111110111101;
      patterns[65007] = 29'b1_111110111101_111_1_111110111101;
      patterns[65008] = 29'b1_111110111110_000_1_111110111110;
      patterns[65009] = 29'b1_111110111110_001_1_111110111110;
      patterns[65010] = 29'b1_111110111110_010_1_111101111101;
      patterns[65011] = 29'b1_111110111110_011_1_111011111011;
      patterns[65012] = 29'b1_111110111110_100_0_111111011111;
      patterns[65013] = 29'b1_111110111110_101_1_011111101111;
      patterns[65014] = 29'b1_111110111110_110_1_111110111110;
      patterns[65015] = 29'b1_111110111110_111_1_111110111110;
      patterns[65016] = 29'b1_111110111111_000_1_111110111111;
      patterns[65017] = 29'b1_111110111111_001_1_111111111110;
      patterns[65018] = 29'b1_111110111111_010_1_111101111111;
      patterns[65019] = 29'b1_111110111111_011_1_111011111111;
      patterns[65020] = 29'b1_111110111111_100_1_111111011111;
      patterns[65021] = 29'b1_111110111111_101_1_111111101111;
      patterns[65022] = 29'b1_111110111111_110_1_111110111111;
      patterns[65023] = 29'b1_111110111111_111_1_111110111111;
      patterns[65024] = 29'b1_111111000000_000_1_111111000000;
      patterns[65025] = 29'b1_111111000000_001_1_000000111111;
      patterns[65026] = 29'b1_111111000000_010_1_111110000001;
      patterns[65027] = 29'b1_111111000000_011_1_111100000011;
      patterns[65028] = 29'b1_111111000000_100_0_111111100000;
      patterns[65029] = 29'b1_111111000000_101_0_011111110000;
      patterns[65030] = 29'b1_111111000000_110_1_111111000000;
      patterns[65031] = 29'b1_111111000000_111_1_111111000000;
      patterns[65032] = 29'b1_111111000001_000_1_111111000001;
      patterns[65033] = 29'b1_111111000001_001_1_000001111111;
      patterns[65034] = 29'b1_111111000001_010_1_111110000011;
      patterns[65035] = 29'b1_111111000001_011_1_111100000111;
      patterns[65036] = 29'b1_111111000001_100_1_111111100000;
      patterns[65037] = 29'b1_111111000001_101_0_111111110000;
      patterns[65038] = 29'b1_111111000001_110_1_111111000001;
      patterns[65039] = 29'b1_111111000001_111_1_111111000001;
      patterns[65040] = 29'b1_111111000010_000_1_111111000010;
      patterns[65041] = 29'b1_111111000010_001_1_000010111111;
      patterns[65042] = 29'b1_111111000010_010_1_111110000101;
      patterns[65043] = 29'b1_111111000010_011_1_111100001011;
      patterns[65044] = 29'b1_111111000010_100_0_111111100001;
      patterns[65045] = 29'b1_111111000010_101_1_011111110000;
      patterns[65046] = 29'b1_111111000010_110_1_111111000010;
      patterns[65047] = 29'b1_111111000010_111_1_111111000010;
      patterns[65048] = 29'b1_111111000011_000_1_111111000011;
      patterns[65049] = 29'b1_111111000011_001_1_000011111111;
      patterns[65050] = 29'b1_111111000011_010_1_111110000111;
      patterns[65051] = 29'b1_111111000011_011_1_111100001111;
      patterns[65052] = 29'b1_111111000011_100_1_111111100001;
      patterns[65053] = 29'b1_111111000011_101_1_111111110000;
      patterns[65054] = 29'b1_111111000011_110_1_111111000011;
      patterns[65055] = 29'b1_111111000011_111_1_111111000011;
      patterns[65056] = 29'b1_111111000100_000_1_111111000100;
      patterns[65057] = 29'b1_111111000100_001_1_000100111111;
      patterns[65058] = 29'b1_111111000100_010_1_111110001001;
      patterns[65059] = 29'b1_111111000100_011_1_111100010011;
      patterns[65060] = 29'b1_111111000100_100_0_111111100010;
      patterns[65061] = 29'b1_111111000100_101_0_011111110001;
      patterns[65062] = 29'b1_111111000100_110_1_111111000100;
      patterns[65063] = 29'b1_111111000100_111_1_111111000100;
      patterns[65064] = 29'b1_111111000101_000_1_111111000101;
      patterns[65065] = 29'b1_111111000101_001_1_000101111111;
      patterns[65066] = 29'b1_111111000101_010_1_111110001011;
      patterns[65067] = 29'b1_111111000101_011_1_111100010111;
      patterns[65068] = 29'b1_111111000101_100_1_111111100010;
      patterns[65069] = 29'b1_111111000101_101_0_111111110001;
      patterns[65070] = 29'b1_111111000101_110_1_111111000101;
      patterns[65071] = 29'b1_111111000101_111_1_111111000101;
      patterns[65072] = 29'b1_111111000110_000_1_111111000110;
      patterns[65073] = 29'b1_111111000110_001_1_000110111111;
      patterns[65074] = 29'b1_111111000110_010_1_111110001101;
      patterns[65075] = 29'b1_111111000110_011_1_111100011011;
      patterns[65076] = 29'b1_111111000110_100_0_111111100011;
      patterns[65077] = 29'b1_111111000110_101_1_011111110001;
      patterns[65078] = 29'b1_111111000110_110_1_111111000110;
      patterns[65079] = 29'b1_111111000110_111_1_111111000110;
      patterns[65080] = 29'b1_111111000111_000_1_111111000111;
      patterns[65081] = 29'b1_111111000111_001_1_000111111111;
      patterns[65082] = 29'b1_111111000111_010_1_111110001111;
      patterns[65083] = 29'b1_111111000111_011_1_111100011111;
      patterns[65084] = 29'b1_111111000111_100_1_111111100011;
      patterns[65085] = 29'b1_111111000111_101_1_111111110001;
      patterns[65086] = 29'b1_111111000111_110_1_111111000111;
      patterns[65087] = 29'b1_111111000111_111_1_111111000111;
      patterns[65088] = 29'b1_111111001000_000_1_111111001000;
      patterns[65089] = 29'b1_111111001000_001_1_001000111111;
      patterns[65090] = 29'b1_111111001000_010_1_111110010001;
      patterns[65091] = 29'b1_111111001000_011_1_111100100011;
      patterns[65092] = 29'b1_111111001000_100_0_111111100100;
      patterns[65093] = 29'b1_111111001000_101_0_011111110010;
      patterns[65094] = 29'b1_111111001000_110_1_111111001000;
      patterns[65095] = 29'b1_111111001000_111_1_111111001000;
      patterns[65096] = 29'b1_111111001001_000_1_111111001001;
      patterns[65097] = 29'b1_111111001001_001_1_001001111111;
      patterns[65098] = 29'b1_111111001001_010_1_111110010011;
      patterns[65099] = 29'b1_111111001001_011_1_111100100111;
      patterns[65100] = 29'b1_111111001001_100_1_111111100100;
      patterns[65101] = 29'b1_111111001001_101_0_111111110010;
      patterns[65102] = 29'b1_111111001001_110_1_111111001001;
      patterns[65103] = 29'b1_111111001001_111_1_111111001001;
      patterns[65104] = 29'b1_111111001010_000_1_111111001010;
      patterns[65105] = 29'b1_111111001010_001_1_001010111111;
      patterns[65106] = 29'b1_111111001010_010_1_111110010101;
      patterns[65107] = 29'b1_111111001010_011_1_111100101011;
      patterns[65108] = 29'b1_111111001010_100_0_111111100101;
      patterns[65109] = 29'b1_111111001010_101_1_011111110010;
      patterns[65110] = 29'b1_111111001010_110_1_111111001010;
      patterns[65111] = 29'b1_111111001010_111_1_111111001010;
      patterns[65112] = 29'b1_111111001011_000_1_111111001011;
      patterns[65113] = 29'b1_111111001011_001_1_001011111111;
      patterns[65114] = 29'b1_111111001011_010_1_111110010111;
      patterns[65115] = 29'b1_111111001011_011_1_111100101111;
      patterns[65116] = 29'b1_111111001011_100_1_111111100101;
      patterns[65117] = 29'b1_111111001011_101_1_111111110010;
      patterns[65118] = 29'b1_111111001011_110_1_111111001011;
      patterns[65119] = 29'b1_111111001011_111_1_111111001011;
      patterns[65120] = 29'b1_111111001100_000_1_111111001100;
      patterns[65121] = 29'b1_111111001100_001_1_001100111111;
      patterns[65122] = 29'b1_111111001100_010_1_111110011001;
      patterns[65123] = 29'b1_111111001100_011_1_111100110011;
      patterns[65124] = 29'b1_111111001100_100_0_111111100110;
      patterns[65125] = 29'b1_111111001100_101_0_011111110011;
      patterns[65126] = 29'b1_111111001100_110_1_111111001100;
      patterns[65127] = 29'b1_111111001100_111_1_111111001100;
      patterns[65128] = 29'b1_111111001101_000_1_111111001101;
      patterns[65129] = 29'b1_111111001101_001_1_001101111111;
      patterns[65130] = 29'b1_111111001101_010_1_111110011011;
      patterns[65131] = 29'b1_111111001101_011_1_111100110111;
      patterns[65132] = 29'b1_111111001101_100_1_111111100110;
      patterns[65133] = 29'b1_111111001101_101_0_111111110011;
      patterns[65134] = 29'b1_111111001101_110_1_111111001101;
      patterns[65135] = 29'b1_111111001101_111_1_111111001101;
      patterns[65136] = 29'b1_111111001110_000_1_111111001110;
      patterns[65137] = 29'b1_111111001110_001_1_001110111111;
      patterns[65138] = 29'b1_111111001110_010_1_111110011101;
      patterns[65139] = 29'b1_111111001110_011_1_111100111011;
      patterns[65140] = 29'b1_111111001110_100_0_111111100111;
      patterns[65141] = 29'b1_111111001110_101_1_011111110011;
      patterns[65142] = 29'b1_111111001110_110_1_111111001110;
      patterns[65143] = 29'b1_111111001110_111_1_111111001110;
      patterns[65144] = 29'b1_111111001111_000_1_111111001111;
      patterns[65145] = 29'b1_111111001111_001_1_001111111111;
      patterns[65146] = 29'b1_111111001111_010_1_111110011111;
      patterns[65147] = 29'b1_111111001111_011_1_111100111111;
      patterns[65148] = 29'b1_111111001111_100_1_111111100111;
      patterns[65149] = 29'b1_111111001111_101_1_111111110011;
      patterns[65150] = 29'b1_111111001111_110_1_111111001111;
      patterns[65151] = 29'b1_111111001111_111_1_111111001111;
      patterns[65152] = 29'b1_111111010000_000_1_111111010000;
      patterns[65153] = 29'b1_111111010000_001_1_010000111111;
      patterns[65154] = 29'b1_111111010000_010_1_111110100001;
      patterns[65155] = 29'b1_111111010000_011_1_111101000011;
      patterns[65156] = 29'b1_111111010000_100_0_111111101000;
      patterns[65157] = 29'b1_111111010000_101_0_011111110100;
      patterns[65158] = 29'b1_111111010000_110_1_111111010000;
      patterns[65159] = 29'b1_111111010000_111_1_111111010000;
      patterns[65160] = 29'b1_111111010001_000_1_111111010001;
      patterns[65161] = 29'b1_111111010001_001_1_010001111111;
      patterns[65162] = 29'b1_111111010001_010_1_111110100011;
      patterns[65163] = 29'b1_111111010001_011_1_111101000111;
      patterns[65164] = 29'b1_111111010001_100_1_111111101000;
      patterns[65165] = 29'b1_111111010001_101_0_111111110100;
      patterns[65166] = 29'b1_111111010001_110_1_111111010001;
      patterns[65167] = 29'b1_111111010001_111_1_111111010001;
      patterns[65168] = 29'b1_111111010010_000_1_111111010010;
      patterns[65169] = 29'b1_111111010010_001_1_010010111111;
      patterns[65170] = 29'b1_111111010010_010_1_111110100101;
      patterns[65171] = 29'b1_111111010010_011_1_111101001011;
      patterns[65172] = 29'b1_111111010010_100_0_111111101001;
      patterns[65173] = 29'b1_111111010010_101_1_011111110100;
      patterns[65174] = 29'b1_111111010010_110_1_111111010010;
      patterns[65175] = 29'b1_111111010010_111_1_111111010010;
      patterns[65176] = 29'b1_111111010011_000_1_111111010011;
      patterns[65177] = 29'b1_111111010011_001_1_010011111111;
      patterns[65178] = 29'b1_111111010011_010_1_111110100111;
      patterns[65179] = 29'b1_111111010011_011_1_111101001111;
      patterns[65180] = 29'b1_111111010011_100_1_111111101001;
      patterns[65181] = 29'b1_111111010011_101_1_111111110100;
      patterns[65182] = 29'b1_111111010011_110_1_111111010011;
      patterns[65183] = 29'b1_111111010011_111_1_111111010011;
      patterns[65184] = 29'b1_111111010100_000_1_111111010100;
      patterns[65185] = 29'b1_111111010100_001_1_010100111111;
      patterns[65186] = 29'b1_111111010100_010_1_111110101001;
      patterns[65187] = 29'b1_111111010100_011_1_111101010011;
      patterns[65188] = 29'b1_111111010100_100_0_111111101010;
      patterns[65189] = 29'b1_111111010100_101_0_011111110101;
      patterns[65190] = 29'b1_111111010100_110_1_111111010100;
      patterns[65191] = 29'b1_111111010100_111_1_111111010100;
      patterns[65192] = 29'b1_111111010101_000_1_111111010101;
      patterns[65193] = 29'b1_111111010101_001_1_010101111111;
      patterns[65194] = 29'b1_111111010101_010_1_111110101011;
      patterns[65195] = 29'b1_111111010101_011_1_111101010111;
      patterns[65196] = 29'b1_111111010101_100_1_111111101010;
      patterns[65197] = 29'b1_111111010101_101_0_111111110101;
      patterns[65198] = 29'b1_111111010101_110_1_111111010101;
      patterns[65199] = 29'b1_111111010101_111_1_111111010101;
      patterns[65200] = 29'b1_111111010110_000_1_111111010110;
      patterns[65201] = 29'b1_111111010110_001_1_010110111111;
      patterns[65202] = 29'b1_111111010110_010_1_111110101101;
      patterns[65203] = 29'b1_111111010110_011_1_111101011011;
      patterns[65204] = 29'b1_111111010110_100_0_111111101011;
      patterns[65205] = 29'b1_111111010110_101_1_011111110101;
      patterns[65206] = 29'b1_111111010110_110_1_111111010110;
      patterns[65207] = 29'b1_111111010110_111_1_111111010110;
      patterns[65208] = 29'b1_111111010111_000_1_111111010111;
      patterns[65209] = 29'b1_111111010111_001_1_010111111111;
      patterns[65210] = 29'b1_111111010111_010_1_111110101111;
      patterns[65211] = 29'b1_111111010111_011_1_111101011111;
      patterns[65212] = 29'b1_111111010111_100_1_111111101011;
      patterns[65213] = 29'b1_111111010111_101_1_111111110101;
      patterns[65214] = 29'b1_111111010111_110_1_111111010111;
      patterns[65215] = 29'b1_111111010111_111_1_111111010111;
      patterns[65216] = 29'b1_111111011000_000_1_111111011000;
      patterns[65217] = 29'b1_111111011000_001_1_011000111111;
      patterns[65218] = 29'b1_111111011000_010_1_111110110001;
      patterns[65219] = 29'b1_111111011000_011_1_111101100011;
      patterns[65220] = 29'b1_111111011000_100_0_111111101100;
      patterns[65221] = 29'b1_111111011000_101_0_011111110110;
      patterns[65222] = 29'b1_111111011000_110_1_111111011000;
      patterns[65223] = 29'b1_111111011000_111_1_111111011000;
      patterns[65224] = 29'b1_111111011001_000_1_111111011001;
      patterns[65225] = 29'b1_111111011001_001_1_011001111111;
      patterns[65226] = 29'b1_111111011001_010_1_111110110011;
      patterns[65227] = 29'b1_111111011001_011_1_111101100111;
      patterns[65228] = 29'b1_111111011001_100_1_111111101100;
      patterns[65229] = 29'b1_111111011001_101_0_111111110110;
      patterns[65230] = 29'b1_111111011001_110_1_111111011001;
      patterns[65231] = 29'b1_111111011001_111_1_111111011001;
      patterns[65232] = 29'b1_111111011010_000_1_111111011010;
      patterns[65233] = 29'b1_111111011010_001_1_011010111111;
      patterns[65234] = 29'b1_111111011010_010_1_111110110101;
      patterns[65235] = 29'b1_111111011010_011_1_111101101011;
      patterns[65236] = 29'b1_111111011010_100_0_111111101101;
      patterns[65237] = 29'b1_111111011010_101_1_011111110110;
      patterns[65238] = 29'b1_111111011010_110_1_111111011010;
      patterns[65239] = 29'b1_111111011010_111_1_111111011010;
      patterns[65240] = 29'b1_111111011011_000_1_111111011011;
      patterns[65241] = 29'b1_111111011011_001_1_011011111111;
      patterns[65242] = 29'b1_111111011011_010_1_111110110111;
      patterns[65243] = 29'b1_111111011011_011_1_111101101111;
      patterns[65244] = 29'b1_111111011011_100_1_111111101101;
      patterns[65245] = 29'b1_111111011011_101_1_111111110110;
      patterns[65246] = 29'b1_111111011011_110_1_111111011011;
      patterns[65247] = 29'b1_111111011011_111_1_111111011011;
      patterns[65248] = 29'b1_111111011100_000_1_111111011100;
      patterns[65249] = 29'b1_111111011100_001_1_011100111111;
      patterns[65250] = 29'b1_111111011100_010_1_111110111001;
      patterns[65251] = 29'b1_111111011100_011_1_111101110011;
      patterns[65252] = 29'b1_111111011100_100_0_111111101110;
      patterns[65253] = 29'b1_111111011100_101_0_011111110111;
      patterns[65254] = 29'b1_111111011100_110_1_111111011100;
      patterns[65255] = 29'b1_111111011100_111_1_111111011100;
      patterns[65256] = 29'b1_111111011101_000_1_111111011101;
      patterns[65257] = 29'b1_111111011101_001_1_011101111111;
      patterns[65258] = 29'b1_111111011101_010_1_111110111011;
      patterns[65259] = 29'b1_111111011101_011_1_111101110111;
      patterns[65260] = 29'b1_111111011101_100_1_111111101110;
      patterns[65261] = 29'b1_111111011101_101_0_111111110111;
      patterns[65262] = 29'b1_111111011101_110_1_111111011101;
      patterns[65263] = 29'b1_111111011101_111_1_111111011101;
      patterns[65264] = 29'b1_111111011110_000_1_111111011110;
      patterns[65265] = 29'b1_111111011110_001_1_011110111111;
      patterns[65266] = 29'b1_111111011110_010_1_111110111101;
      patterns[65267] = 29'b1_111111011110_011_1_111101111011;
      patterns[65268] = 29'b1_111111011110_100_0_111111101111;
      patterns[65269] = 29'b1_111111011110_101_1_011111110111;
      patterns[65270] = 29'b1_111111011110_110_1_111111011110;
      patterns[65271] = 29'b1_111111011110_111_1_111111011110;
      patterns[65272] = 29'b1_111111011111_000_1_111111011111;
      patterns[65273] = 29'b1_111111011111_001_1_011111111111;
      patterns[65274] = 29'b1_111111011111_010_1_111110111111;
      patterns[65275] = 29'b1_111111011111_011_1_111101111111;
      patterns[65276] = 29'b1_111111011111_100_1_111111101111;
      patterns[65277] = 29'b1_111111011111_101_1_111111110111;
      patterns[65278] = 29'b1_111111011111_110_1_111111011111;
      patterns[65279] = 29'b1_111111011111_111_1_111111011111;
      patterns[65280] = 29'b1_111111100000_000_1_111111100000;
      patterns[65281] = 29'b1_111111100000_001_1_100000111111;
      patterns[65282] = 29'b1_111111100000_010_1_111111000001;
      patterns[65283] = 29'b1_111111100000_011_1_111110000011;
      patterns[65284] = 29'b1_111111100000_100_0_111111110000;
      patterns[65285] = 29'b1_111111100000_101_0_011111111000;
      patterns[65286] = 29'b1_111111100000_110_1_111111100000;
      patterns[65287] = 29'b1_111111100000_111_1_111111100000;
      patterns[65288] = 29'b1_111111100001_000_1_111111100001;
      patterns[65289] = 29'b1_111111100001_001_1_100001111111;
      patterns[65290] = 29'b1_111111100001_010_1_111111000011;
      patterns[65291] = 29'b1_111111100001_011_1_111110000111;
      patterns[65292] = 29'b1_111111100001_100_1_111111110000;
      patterns[65293] = 29'b1_111111100001_101_0_111111111000;
      patterns[65294] = 29'b1_111111100001_110_1_111111100001;
      patterns[65295] = 29'b1_111111100001_111_1_111111100001;
      patterns[65296] = 29'b1_111111100010_000_1_111111100010;
      patterns[65297] = 29'b1_111111100010_001_1_100010111111;
      patterns[65298] = 29'b1_111111100010_010_1_111111000101;
      patterns[65299] = 29'b1_111111100010_011_1_111110001011;
      patterns[65300] = 29'b1_111111100010_100_0_111111110001;
      patterns[65301] = 29'b1_111111100010_101_1_011111111000;
      patterns[65302] = 29'b1_111111100010_110_1_111111100010;
      patterns[65303] = 29'b1_111111100010_111_1_111111100010;
      patterns[65304] = 29'b1_111111100011_000_1_111111100011;
      patterns[65305] = 29'b1_111111100011_001_1_100011111111;
      patterns[65306] = 29'b1_111111100011_010_1_111111000111;
      patterns[65307] = 29'b1_111111100011_011_1_111110001111;
      patterns[65308] = 29'b1_111111100011_100_1_111111110001;
      patterns[65309] = 29'b1_111111100011_101_1_111111111000;
      patterns[65310] = 29'b1_111111100011_110_1_111111100011;
      patterns[65311] = 29'b1_111111100011_111_1_111111100011;
      patterns[65312] = 29'b1_111111100100_000_1_111111100100;
      patterns[65313] = 29'b1_111111100100_001_1_100100111111;
      patterns[65314] = 29'b1_111111100100_010_1_111111001001;
      patterns[65315] = 29'b1_111111100100_011_1_111110010011;
      patterns[65316] = 29'b1_111111100100_100_0_111111110010;
      patterns[65317] = 29'b1_111111100100_101_0_011111111001;
      patterns[65318] = 29'b1_111111100100_110_1_111111100100;
      patterns[65319] = 29'b1_111111100100_111_1_111111100100;
      patterns[65320] = 29'b1_111111100101_000_1_111111100101;
      patterns[65321] = 29'b1_111111100101_001_1_100101111111;
      patterns[65322] = 29'b1_111111100101_010_1_111111001011;
      patterns[65323] = 29'b1_111111100101_011_1_111110010111;
      patterns[65324] = 29'b1_111111100101_100_1_111111110010;
      patterns[65325] = 29'b1_111111100101_101_0_111111111001;
      patterns[65326] = 29'b1_111111100101_110_1_111111100101;
      patterns[65327] = 29'b1_111111100101_111_1_111111100101;
      patterns[65328] = 29'b1_111111100110_000_1_111111100110;
      patterns[65329] = 29'b1_111111100110_001_1_100110111111;
      patterns[65330] = 29'b1_111111100110_010_1_111111001101;
      patterns[65331] = 29'b1_111111100110_011_1_111110011011;
      patterns[65332] = 29'b1_111111100110_100_0_111111110011;
      patterns[65333] = 29'b1_111111100110_101_1_011111111001;
      patterns[65334] = 29'b1_111111100110_110_1_111111100110;
      patterns[65335] = 29'b1_111111100110_111_1_111111100110;
      patterns[65336] = 29'b1_111111100111_000_1_111111100111;
      patterns[65337] = 29'b1_111111100111_001_1_100111111111;
      patterns[65338] = 29'b1_111111100111_010_1_111111001111;
      patterns[65339] = 29'b1_111111100111_011_1_111110011111;
      patterns[65340] = 29'b1_111111100111_100_1_111111110011;
      patterns[65341] = 29'b1_111111100111_101_1_111111111001;
      patterns[65342] = 29'b1_111111100111_110_1_111111100111;
      patterns[65343] = 29'b1_111111100111_111_1_111111100111;
      patterns[65344] = 29'b1_111111101000_000_1_111111101000;
      patterns[65345] = 29'b1_111111101000_001_1_101000111111;
      patterns[65346] = 29'b1_111111101000_010_1_111111010001;
      patterns[65347] = 29'b1_111111101000_011_1_111110100011;
      patterns[65348] = 29'b1_111111101000_100_0_111111110100;
      patterns[65349] = 29'b1_111111101000_101_0_011111111010;
      patterns[65350] = 29'b1_111111101000_110_1_111111101000;
      patterns[65351] = 29'b1_111111101000_111_1_111111101000;
      patterns[65352] = 29'b1_111111101001_000_1_111111101001;
      patterns[65353] = 29'b1_111111101001_001_1_101001111111;
      patterns[65354] = 29'b1_111111101001_010_1_111111010011;
      patterns[65355] = 29'b1_111111101001_011_1_111110100111;
      patterns[65356] = 29'b1_111111101001_100_1_111111110100;
      patterns[65357] = 29'b1_111111101001_101_0_111111111010;
      patterns[65358] = 29'b1_111111101001_110_1_111111101001;
      patterns[65359] = 29'b1_111111101001_111_1_111111101001;
      patterns[65360] = 29'b1_111111101010_000_1_111111101010;
      patterns[65361] = 29'b1_111111101010_001_1_101010111111;
      patterns[65362] = 29'b1_111111101010_010_1_111111010101;
      patterns[65363] = 29'b1_111111101010_011_1_111110101011;
      patterns[65364] = 29'b1_111111101010_100_0_111111110101;
      patterns[65365] = 29'b1_111111101010_101_1_011111111010;
      patterns[65366] = 29'b1_111111101010_110_1_111111101010;
      patterns[65367] = 29'b1_111111101010_111_1_111111101010;
      patterns[65368] = 29'b1_111111101011_000_1_111111101011;
      patterns[65369] = 29'b1_111111101011_001_1_101011111111;
      patterns[65370] = 29'b1_111111101011_010_1_111111010111;
      patterns[65371] = 29'b1_111111101011_011_1_111110101111;
      patterns[65372] = 29'b1_111111101011_100_1_111111110101;
      patterns[65373] = 29'b1_111111101011_101_1_111111111010;
      patterns[65374] = 29'b1_111111101011_110_1_111111101011;
      patterns[65375] = 29'b1_111111101011_111_1_111111101011;
      patterns[65376] = 29'b1_111111101100_000_1_111111101100;
      patterns[65377] = 29'b1_111111101100_001_1_101100111111;
      patterns[65378] = 29'b1_111111101100_010_1_111111011001;
      patterns[65379] = 29'b1_111111101100_011_1_111110110011;
      patterns[65380] = 29'b1_111111101100_100_0_111111110110;
      patterns[65381] = 29'b1_111111101100_101_0_011111111011;
      patterns[65382] = 29'b1_111111101100_110_1_111111101100;
      patterns[65383] = 29'b1_111111101100_111_1_111111101100;
      patterns[65384] = 29'b1_111111101101_000_1_111111101101;
      patterns[65385] = 29'b1_111111101101_001_1_101101111111;
      patterns[65386] = 29'b1_111111101101_010_1_111111011011;
      patterns[65387] = 29'b1_111111101101_011_1_111110110111;
      patterns[65388] = 29'b1_111111101101_100_1_111111110110;
      patterns[65389] = 29'b1_111111101101_101_0_111111111011;
      patterns[65390] = 29'b1_111111101101_110_1_111111101101;
      patterns[65391] = 29'b1_111111101101_111_1_111111101101;
      patterns[65392] = 29'b1_111111101110_000_1_111111101110;
      patterns[65393] = 29'b1_111111101110_001_1_101110111111;
      patterns[65394] = 29'b1_111111101110_010_1_111111011101;
      patterns[65395] = 29'b1_111111101110_011_1_111110111011;
      patterns[65396] = 29'b1_111111101110_100_0_111111110111;
      patterns[65397] = 29'b1_111111101110_101_1_011111111011;
      patterns[65398] = 29'b1_111111101110_110_1_111111101110;
      patterns[65399] = 29'b1_111111101110_111_1_111111101110;
      patterns[65400] = 29'b1_111111101111_000_1_111111101111;
      patterns[65401] = 29'b1_111111101111_001_1_101111111111;
      patterns[65402] = 29'b1_111111101111_010_1_111111011111;
      patterns[65403] = 29'b1_111111101111_011_1_111110111111;
      patterns[65404] = 29'b1_111111101111_100_1_111111110111;
      patterns[65405] = 29'b1_111111101111_101_1_111111111011;
      patterns[65406] = 29'b1_111111101111_110_1_111111101111;
      patterns[65407] = 29'b1_111111101111_111_1_111111101111;
      patterns[65408] = 29'b1_111111110000_000_1_111111110000;
      patterns[65409] = 29'b1_111111110000_001_1_110000111111;
      patterns[65410] = 29'b1_111111110000_010_1_111111100001;
      patterns[65411] = 29'b1_111111110000_011_1_111111000011;
      patterns[65412] = 29'b1_111111110000_100_0_111111111000;
      patterns[65413] = 29'b1_111111110000_101_0_011111111100;
      patterns[65414] = 29'b1_111111110000_110_1_111111110000;
      patterns[65415] = 29'b1_111111110000_111_1_111111110000;
      patterns[65416] = 29'b1_111111110001_000_1_111111110001;
      patterns[65417] = 29'b1_111111110001_001_1_110001111111;
      patterns[65418] = 29'b1_111111110001_010_1_111111100011;
      patterns[65419] = 29'b1_111111110001_011_1_111111000111;
      patterns[65420] = 29'b1_111111110001_100_1_111111111000;
      patterns[65421] = 29'b1_111111110001_101_0_111111111100;
      patterns[65422] = 29'b1_111111110001_110_1_111111110001;
      patterns[65423] = 29'b1_111111110001_111_1_111111110001;
      patterns[65424] = 29'b1_111111110010_000_1_111111110010;
      patterns[65425] = 29'b1_111111110010_001_1_110010111111;
      patterns[65426] = 29'b1_111111110010_010_1_111111100101;
      patterns[65427] = 29'b1_111111110010_011_1_111111001011;
      patterns[65428] = 29'b1_111111110010_100_0_111111111001;
      patterns[65429] = 29'b1_111111110010_101_1_011111111100;
      patterns[65430] = 29'b1_111111110010_110_1_111111110010;
      patterns[65431] = 29'b1_111111110010_111_1_111111110010;
      patterns[65432] = 29'b1_111111110011_000_1_111111110011;
      patterns[65433] = 29'b1_111111110011_001_1_110011111111;
      patterns[65434] = 29'b1_111111110011_010_1_111111100111;
      patterns[65435] = 29'b1_111111110011_011_1_111111001111;
      patterns[65436] = 29'b1_111111110011_100_1_111111111001;
      patterns[65437] = 29'b1_111111110011_101_1_111111111100;
      patterns[65438] = 29'b1_111111110011_110_1_111111110011;
      patterns[65439] = 29'b1_111111110011_111_1_111111110011;
      patterns[65440] = 29'b1_111111110100_000_1_111111110100;
      patterns[65441] = 29'b1_111111110100_001_1_110100111111;
      patterns[65442] = 29'b1_111111110100_010_1_111111101001;
      patterns[65443] = 29'b1_111111110100_011_1_111111010011;
      patterns[65444] = 29'b1_111111110100_100_0_111111111010;
      patterns[65445] = 29'b1_111111110100_101_0_011111111101;
      patterns[65446] = 29'b1_111111110100_110_1_111111110100;
      patterns[65447] = 29'b1_111111110100_111_1_111111110100;
      patterns[65448] = 29'b1_111111110101_000_1_111111110101;
      patterns[65449] = 29'b1_111111110101_001_1_110101111111;
      patterns[65450] = 29'b1_111111110101_010_1_111111101011;
      patterns[65451] = 29'b1_111111110101_011_1_111111010111;
      patterns[65452] = 29'b1_111111110101_100_1_111111111010;
      patterns[65453] = 29'b1_111111110101_101_0_111111111101;
      patterns[65454] = 29'b1_111111110101_110_1_111111110101;
      patterns[65455] = 29'b1_111111110101_111_1_111111110101;
      patterns[65456] = 29'b1_111111110110_000_1_111111110110;
      patterns[65457] = 29'b1_111111110110_001_1_110110111111;
      patterns[65458] = 29'b1_111111110110_010_1_111111101101;
      patterns[65459] = 29'b1_111111110110_011_1_111111011011;
      patterns[65460] = 29'b1_111111110110_100_0_111111111011;
      patterns[65461] = 29'b1_111111110110_101_1_011111111101;
      patterns[65462] = 29'b1_111111110110_110_1_111111110110;
      patterns[65463] = 29'b1_111111110110_111_1_111111110110;
      patterns[65464] = 29'b1_111111110111_000_1_111111110111;
      patterns[65465] = 29'b1_111111110111_001_1_110111111111;
      patterns[65466] = 29'b1_111111110111_010_1_111111101111;
      patterns[65467] = 29'b1_111111110111_011_1_111111011111;
      patterns[65468] = 29'b1_111111110111_100_1_111111111011;
      patterns[65469] = 29'b1_111111110111_101_1_111111111101;
      patterns[65470] = 29'b1_111111110111_110_1_111111110111;
      patterns[65471] = 29'b1_111111110111_111_1_111111110111;
      patterns[65472] = 29'b1_111111111000_000_1_111111111000;
      patterns[65473] = 29'b1_111111111000_001_1_111000111111;
      patterns[65474] = 29'b1_111111111000_010_1_111111110001;
      patterns[65475] = 29'b1_111111111000_011_1_111111100011;
      patterns[65476] = 29'b1_111111111000_100_0_111111111100;
      patterns[65477] = 29'b1_111111111000_101_0_011111111110;
      patterns[65478] = 29'b1_111111111000_110_1_111111111000;
      patterns[65479] = 29'b1_111111111000_111_1_111111111000;
      patterns[65480] = 29'b1_111111111001_000_1_111111111001;
      patterns[65481] = 29'b1_111111111001_001_1_111001111111;
      patterns[65482] = 29'b1_111111111001_010_1_111111110011;
      patterns[65483] = 29'b1_111111111001_011_1_111111100111;
      patterns[65484] = 29'b1_111111111001_100_1_111111111100;
      patterns[65485] = 29'b1_111111111001_101_0_111111111110;
      patterns[65486] = 29'b1_111111111001_110_1_111111111001;
      patterns[65487] = 29'b1_111111111001_111_1_111111111001;
      patterns[65488] = 29'b1_111111111010_000_1_111111111010;
      patterns[65489] = 29'b1_111111111010_001_1_111010111111;
      patterns[65490] = 29'b1_111111111010_010_1_111111110101;
      patterns[65491] = 29'b1_111111111010_011_1_111111101011;
      patterns[65492] = 29'b1_111111111010_100_0_111111111101;
      patterns[65493] = 29'b1_111111111010_101_1_011111111110;
      patterns[65494] = 29'b1_111111111010_110_1_111111111010;
      patterns[65495] = 29'b1_111111111010_111_1_111111111010;
      patterns[65496] = 29'b1_111111111011_000_1_111111111011;
      patterns[65497] = 29'b1_111111111011_001_1_111011111111;
      patterns[65498] = 29'b1_111111111011_010_1_111111110111;
      patterns[65499] = 29'b1_111111111011_011_1_111111101111;
      patterns[65500] = 29'b1_111111111011_100_1_111111111101;
      patterns[65501] = 29'b1_111111111011_101_1_111111111110;
      patterns[65502] = 29'b1_111111111011_110_1_111111111011;
      patterns[65503] = 29'b1_111111111011_111_1_111111111011;
      patterns[65504] = 29'b1_111111111100_000_1_111111111100;
      patterns[65505] = 29'b1_111111111100_001_1_111100111111;
      patterns[65506] = 29'b1_111111111100_010_1_111111111001;
      patterns[65507] = 29'b1_111111111100_011_1_111111110011;
      patterns[65508] = 29'b1_111111111100_100_0_111111111110;
      patterns[65509] = 29'b1_111111111100_101_0_011111111111;
      patterns[65510] = 29'b1_111111111100_110_1_111111111100;
      patterns[65511] = 29'b1_111111111100_111_1_111111111100;
      patterns[65512] = 29'b1_111111111101_000_1_111111111101;
      patterns[65513] = 29'b1_111111111101_001_1_111101111111;
      patterns[65514] = 29'b1_111111111101_010_1_111111111011;
      patterns[65515] = 29'b1_111111111101_011_1_111111110111;
      patterns[65516] = 29'b1_111111111101_100_1_111111111110;
      patterns[65517] = 29'b1_111111111101_101_0_111111111111;
      patterns[65518] = 29'b1_111111111101_110_1_111111111101;
      patterns[65519] = 29'b1_111111111101_111_1_111111111101;
      patterns[65520] = 29'b1_111111111110_000_1_111111111110;
      patterns[65521] = 29'b1_111111111110_001_1_111110111111;
      patterns[65522] = 29'b1_111111111110_010_1_111111111101;
      patterns[65523] = 29'b1_111111111110_011_1_111111111011;
      patterns[65524] = 29'b1_111111111110_100_0_111111111111;
      patterns[65525] = 29'b1_111111111110_101_1_011111111111;
      patterns[65526] = 29'b1_111111111110_110_1_111111111110;
      patterns[65527] = 29'b1_111111111110_111_1_111111111110;
      patterns[65528] = 29'b1_111111111111_000_1_111111111111;
      patterns[65529] = 29'b1_111111111111_001_1_111111111111;
      patterns[65530] = 29'b1_111111111111_010_1_111111111111;
      patterns[65531] = 29'b1_111111111111_011_1_111111111111;
      patterns[65532] = 29'b1_111111111111_100_1_111111111111;
      patterns[65533] = 29'b1_111111111111_101_1_111111111111;
      patterns[65534] = 29'b1_111111111111_110_1_111111111111;
      patterns[65535] = 29'b1_111111111111_111_1_111111111111;

      for (i = 0; i < 65536; i = i + 1)
      begin
        LI = patterns[i][28];
        AI = patterns[i][27:16];
        OP = patterns[i][15:13];
        #10;
        if (patterns[i][12] !== 1'hx)
        begin
          if (LO !== patterns[i][12])
          begin
            $display("%d:LO: (assertion error). Expected %h, found %h", i, patterns[i][12], LO);
            $finish;
          end
        end
        if (patterns[i][11:0] !== 12'hx)
        begin
          if (AO !== patterns[i][11:0])
          begin
            $display("%d:AO: (assertion error). Expected %h, found %h", i, patterns[i][11:0], AO);
            $finish;
          end
        end
      end

      $display("All tests passed.");
    end
    endmodule
