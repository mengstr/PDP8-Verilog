//  A testbench for UART-RX_simple_tb
`timescale 1us/1ns

module UART-RX_simple_tb;
    reg RX;
    reg clk16;
    reg CDP;
    reg en;
    wire [7:0] DATA;
    wire DP;
    wire busy;

  \UART-RX  \UART-RX 0 (
    .RX(RX),
    .clk16(clk16),
    .CDP(CDP),
    .en(en),
    .DATA(DATA),
    .DP(DP),
    .busy(busy)
  );

    reg [11:0] patterns[0:992];
    integer i;

    initial begin
      patterns[0] = 12'b0_0_0_xxxxxxxx_x;
      patterns[1] = 12'b0_1_0_xxxxxxxx_x;
      patterns[2] = 12'b0_0_0_xxxxxxxx_0;
      patterns[3] = 12'b0_0_0_xxxxxxxx_x;
      patterns[4] = 12'b0_1_0_xxxxxxxx_x;
      patterns[5] = 12'b0_0_0_xxxxxxxx_0;
      patterns[6] = 12'b0_0_0_xxxxxxxx_x;
      patterns[7] = 12'b0_1_0_xxxxxxxx_x;
      patterns[8] = 12'b0_0_0_xxxxxxxx_0;
      patterns[9] = 12'b0_0_0_xxxxxxxx_x;
      patterns[10] = 12'b0_1_0_xxxxxxxx_x;
      patterns[11] = 12'b0_0_0_xxxxxxxx_0;
      patterns[12] = 12'b0_0_0_xxxxxxxx_x;
      patterns[13] = 12'b0_1_0_xxxxxxxx_x;
      patterns[14] = 12'b0_0_0_xxxxxxxx_0;
      patterns[15] = 12'b0_0_1_xxxxxxxx_x;
      patterns[16] = 12'b0_1_1_xxxxxxxx_x;
      patterns[17] = 12'b0_0_1_xxxxxxxx_0;
      patterns[18] = 12'b0_0_1_xxxxxxxx_x;
      patterns[19] = 12'b0_1_1_xxxxxxxx_x;
      patterns[20] = 12'b0_0_1_xxxxxxxx_0;
      patterns[21] = 12'b0_0_1_xxxxxxxx_x;
      patterns[22] = 12'b0_1_1_xxxxxxxx_x;
      patterns[23] = 12'b0_0_1_xxxxxxxx_0;
      patterns[24] = 12'b0_0_1_xxxxxxxx_x;
      patterns[25] = 12'b0_1_1_xxxxxxxx_x;
      patterns[26] = 12'b0_0_1_xxxxxxxx_0;
      patterns[27] = 12'b0_0_1_xxxxxxxx_x;
      patterns[28] = 12'b0_1_1_xxxxxxxx_x;
      patterns[29] = 12'b0_0_1_xxxxxxxx_0;
      patterns[30] = 12'b0_0_1_xxxxxxxx_x;
      patterns[31] = 12'b0_1_1_xxxxxxxx_x;
      patterns[32] = 12'b0_0_1_xxxxxxxx_0;
      patterns[33] = 12'b0_0_1_xxxxxxxx_x;
      patterns[34] = 12'b0_1_1_xxxxxxxx_x;
      patterns[35] = 12'b0_0_1_xxxxxxxx_0;
      patterns[36] = 12'b0_0_1_xxxxxxxx_x;
      patterns[37] = 12'b0_1_1_xxxxxxxx_x;
      patterns[38] = 12'b0_0_1_xxxxxxxx_0;
      patterns[39] = 12'b0_0_1_xxxxxxxx_x;
      patterns[40] = 12'b0_1_1_xxxxxxxx_x;
      patterns[41] = 12'b0_0_1_xxxxxxxx_0;
      patterns[42] = 12'b0_0_1_xxxxxxxx_x;
      patterns[43] = 12'b0_1_1_xxxxxxxx_x;
      patterns[44] = 12'b0_0_1_xxxxxxxx_0;
      patterns[45] = 12'b0_0_1_xxxxxxxx_x;
      patterns[46] = 12'b0_1_1_xxxxxxxx_x;
      patterns[47] = 12'b0_0_1_xxxxxxxx_0;
      patterns[48] = 12'b0_0_1_xxxxxxxx_x;
      patterns[49] = 12'b0_1_1_xxxxxxxx_x;
      patterns[50] = 12'b0_0_1_xxxxxxxx_0;
      patterns[51] = 12'b0_0_1_xxxxxxxx_x;
      patterns[52] = 12'b0_1_1_xxxxxxxx_x;
      patterns[53] = 12'b0_0_1_xxxxxxxx_0;
      patterns[54] = 12'b0_0_1_xxxxxxxx_x;
      patterns[55] = 12'b0_1_1_xxxxxxxx_x;
      patterns[56] = 12'b0_0_1_xxxxxxxx_0;
      patterns[57] = 12'b0_0_1_xxxxxxxx_x;
      patterns[58] = 12'b0_1_1_xxxxxxxx_x;
      patterns[59] = 12'b0_0_1_xxxxxxxx_0;
      patterns[60] = 12'b0_0_1_xxxxxxxx_x;
      patterns[61] = 12'b0_1_1_xxxxxxxx_x;
      patterns[62] = 12'b0_0_1_xxxxxxxx_0;
      patterns[63] = 12'b0_0_0_xxxxxxxx_x;
      patterns[64] = 12'b0_1_0_xxxxxxxx_x;
      patterns[65] = 12'b0_0_0_xxxxxxxx_0;
      patterns[66] = 12'b0_0_0_xxxxxxxx_x;
      patterns[67] = 12'b0_1_0_xxxxxxxx_x;
      patterns[68] = 12'b0_0_0_xxxxxxxx_0;
      patterns[69] = 12'b0_0_0_xxxxxxxx_x;
      patterns[70] = 12'b0_1_0_xxxxxxxx_x;
      patterns[71] = 12'b0_0_0_xxxxxxxx_0;
      patterns[72] = 12'b0_0_0_xxxxxxxx_x;
      patterns[73] = 12'b0_1_0_xxxxxxxx_x;
      patterns[74] = 12'b0_0_0_xxxxxxxx_0;
      patterns[75] = 12'b0_0_0_xxxxxxxx_x;
      patterns[76] = 12'b0_1_0_xxxxxxxx_x;
      patterns[77] = 12'b0_0_0_xxxxxxxx_0;
      patterns[78] = 12'b0_0_0_xxxxxxxx_x;
      patterns[79] = 12'b0_1_0_xxxxxxxx_x;
      patterns[80] = 12'b0_0_0_xxxxxxxx_0;
      patterns[81] = 12'b0_0_0_xxxxxxxx_x;
      patterns[82] = 12'b0_1_0_xxxxxxxx_x;
      patterns[83] = 12'b0_0_0_xxxxxxxx_0;
      patterns[84] = 12'b0_0_0_xxxxxxxx_x;
      patterns[85] = 12'b0_1_0_xxxxxxxx_x;
      patterns[86] = 12'b0_0_0_xxxxxxxx_0;
      patterns[87] = 12'b0_0_0_xxxxxxxx_x;
      patterns[88] = 12'b0_1_0_xxxxxxxx_x;
      patterns[89] = 12'b0_0_0_xxxxxxxx_0;
      patterns[90] = 12'b0_0_0_xxxxxxxx_x;
      patterns[91] = 12'b0_1_0_xxxxxxxx_x;
      patterns[92] = 12'b0_0_0_xxxxxxxx_0;
      patterns[93] = 12'b0_0_0_xxxxxxxx_x;
      patterns[94] = 12'b0_1_0_xxxxxxxx_x;
      patterns[95] = 12'b0_0_0_xxxxxxxx_0;
      patterns[96] = 12'b0_0_0_xxxxxxxx_x;
      patterns[97] = 12'b0_1_0_xxxxxxxx_x;
      patterns[98] = 12'b0_0_0_xxxxxxxx_0;
      patterns[99] = 12'b0_0_0_xxxxxxxx_x;
      patterns[100] = 12'b0_1_0_xxxxxxxx_x;
      patterns[101] = 12'b0_0_0_xxxxxxxx_0;
      patterns[102] = 12'b0_0_0_xxxxxxxx_x;
      patterns[103] = 12'b0_1_0_xxxxxxxx_x;
      patterns[104] = 12'b0_0_0_xxxxxxxx_0;
      patterns[105] = 12'b0_0_0_xxxxxxxx_x;
      patterns[106] = 12'b0_1_0_xxxxxxxx_x;
      patterns[107] = 12'b0_0_0_xxxxxxxx_0;
      patterns[108] = 12'b0_0_0_xxxxxxxx_x;
      patterns[109] = 12'b0_1_0_xxxxxxxx_x;
      patterns[110] = 12'b0_0_0_xxxxxxxx_0;
      patterns[111] = 12'b0_0_1_xxxxxxxx_x;
      patterns[112] = 12'b0_1_1_xxxxxxxx_x;
      patterns[113] = 12'b0_0_1_xxxxxxxx_0;
      patterns[114] = 12'b0_0_1_xxxxxxxx_x;
      patterns[115] = 12'b0_1_1_xxxxxxxx_x;
      patterns[116] = 12'b0_0_1_xxxxxxxx_0;
      patterns[117] = 12'b0_0_1_xxxxxxxx_x;
      patterns[118] = 12'b0_1_1_xxxxxxxx_x;
      patterns[119] = 12'b0_0_1_xxxxxxxx_0;
      patterns[120] = 12'b0_0_1_xxxxxxxx_x;
      patterns[121] = 12'b0_1_1_xxxxxxxx_x;
      patterns[122] = 12'b0_0_1_xxxxxxxx_0;
      patterns[123] = 12'b0_0_1_xxxxxxxx_x;
      patterns[124] = 12'b0_1_1_xxxxxxxx_x;
      patterns[125] = 12'b0_0_1_xxxxxxxx_0;
      patterns[126] = 12'b0_0_1_xxxxxxxx_x;
      patterns[127] = 12'b0_1_1_xxxxxxxx_x;
      patterns[128] = 12'b0_0_1_xxxxxxxx_0;
      patterns[129] = 12'b0_0_1_xxxxxxxx_x;
      patterns[130] = 12'b0_1_1_xxxxxxxx_x;
      patterns[131] = 12'b0_0_1_xxxxxxxx_0;
      patterns[132] = 12'b0_0_1_xxxxxxxx_x;
      patterns[133] = 12'b0_1_1_xxxxxxxx_x;
      patterns[134] = 12'b0_0_1_xxxxxxxx_0;
      patterns[135] = 12'b0_0_1_xxxxxxxx_x;
      patterns[136] = 12'b0_1_1_xxxxxxxx_x;
      patterns[137] = 12'b0_0_1_xxxxxxxx_0;
      patterns[138] = 12'b0_0_1_xxxxxxxx_x;
      patterns[139] = 12'b0_1_1_xxxxxxxx_x;
      patterns[140] = 12'b0_0_1_xxxxxxxx_0;
      patterns[141] = 12'b0_0_1_xxxxxxxx_x;
      patterns[142] = 12'b0_1_1_xxxxxxxx_x;
      patterns[143] = 12'b0_0_1_xxxxxxxx_0;
      patterns[144] = 12'b0_0_1_xxxxxxxx_x;
      patterns[145] = 12'b0_1_1_xxxxxxxx_x;
      patterns[146] = 12'b0_0_1_xxxxxxxx_0;
      patterns[147] = 12'b0_0_1_xxxxxxxx_x;
      patterns[148] = 12'b0_1_1_xxxxxxxx_x;
      patterns[149] = 12'b0_0_1_xxxxxxxx_0;
      patterns[150] = 12'b0_0_1_xxxxxxxx_x;
      patterns[151] = 12'b0_1_1_xxxxxxxx_x;
      patterns[152] = 12'b0_0_1_xxxxxxxx_0;
      patterns[153] = 12'b0_0_1_xxxxxxxx_x;
      patterns[154] = 12'b0_1_1_xxxxxxxx_x;
      patterns[155] = 12'b0_0_1_xxxxxxxx_0;
      patterns[156] = 12'b0_0_1_xxxxxxxx_x;
      patterns[157] = 12'b0_1_1_xxxxxxxx_x;
      patterns[158] = 12'b0_0_1_xxxxxxxx_0;
      patterns[159] = 12'b0_0_0_xxxxxxxx_x;
      patterns[160] = 12'b0_1_0_xxxxxxxx_x;
      patterns[161] = 12'b0_0_0_xxxxxxxx_0;
      patterns[162] = 12'b0_0_0_xxxxxxxx_x;
      patterns[163] = 12'b0_1_0_xxxxxxxx_x;
      patterns[164] = 12'b0_0_0_xxxxxxxx_0;
      patterns[165] = 12'b0_0_0_xxxxxxxx_x;
      patterns[166] = 12'b0_1_0_xxxxxxxx_x;
      patterns[167] = 12'b0_0_0_xxxxxxxx_0;
      patterns[168] = 12'b0_0_0_xxxxxxxx_x;
      patterns[169] = 12'b0_1_0_xxxxxxxx_x;
      patterns[170] = 12'b0_0_0_xxxxxxxx_0;
      patterns[171] = 12'b0_0_0_xxxxxxxx_x;
      patterns[172] = 12'b0_1_0_xxxxxxxx_x;
      patterns[173] = 12'b0_0_0_xxxxxxxx_0;
      patterns[174] = 12'b0_0_0_xxxxxxxx_x;
      patterns[175] = 12'b0_1_0_xxxxxxxx_x;
      patterns[176] = 12'b0_0_0_xxxxxxxx_0;
      patterns[177] = 12'b0_0_0_xxxxxxxx_x;
      patterns[178] = 12'b0_1_0_xxxxxxxx_x;
      patterns[179] = 12'b0_0_0_xxxxxxxx_0;
      patterns[180] = 12'b0_0_0_xxxxxxxx_x;
      patterns[181] = 12'b0_1_0_xxxxxxxx_x;
      patterns[182] = 12'b0_0_0_xxxxxxxx_0;
      patterns[183] = 12'b0_0_0_xxxxxxxx_x;
      patterns[184] = 12'b0_1_0_xxxxxxxx_x;
      patterns[185] = 12'b0_0_0_xxxxxxxx_0;
      patterns[186] = 12'b0_0_0_xxxxxxxx_x;
      patterns[187] = 12'b0_1_0_xxxxxxxx_x;
      patterns[188] = 12'b0_0_0_xxxxxxxx_0;
      patterns[189] = 12'b0_0_0_xxxxxxxx_x;
      patterns[190] = 12'b0_1_0_xxxxxxxx_x;
      patterns[191] = 12'b0_0_0_xxxxxxxx_0;
      patterns[192] = 12'b0_0_0_xxxxxxxx_x;
      patterns[193] = 12'b0_1_0_xxxxxxxx_x;
      patterns[194] = 12'b0_0_0_xxxxxxxx_0;
      patterns[195] = 12'b0_0_0_xxxxxxxx_x;
      patterns[196] = 12'b0_1_0_xxxxxxxx_x;
      patterns[197] = 12'b0_0_0_xxxxxxxx_0;
      patterns[198] = 12'b0_0_0_xxxxxxxx_x;
      patterns[199] = 12'b0_1_0_xxxxxxxx_x;
      patterns[200] = 12'b0_0_0_xxxxxxxx_0;
      patterns[201] = 12'b0_0_0_xxxxxxxx_x;
      patterns[202] = 12'b0_1_0_xxxxxxxx_x;
      patterns[203] = 12'b0_0_0_xxxxxxxx_0;
      patterns[204] = 12'b0_0_0_xxxxxxxx_x;
      patterns[205] = 12'b0_1_0_xxxxxxxx_x;
      patterns[206] = 12'b0_0_0_xxxxxxxx_0;
      patterns[207] = 12'b0_0_1_xxxxxxxx_x;
      patterns[208] = 12'b0_1_1_xxxxxxxx_x;
      patterns[209] = 12'b0_0_1_xxxxxxxx_0;
      patterns[210] = 12'b0_0_1_xxxxxxxx_x;
      patterns[211] = 12'b0_1_1_xxxxxxxx_x;
      patterns[212] = 12'b0_0_1_xxxxxxxx_0;
      patterns[213] = 12'b0_0_1_xxxxxxxx_x;
      patterns[214] = 12'b0_1_1_xxxxxxxx_x;
      patterns[215] = 12'b0_0_1_xxxxxxxx_0;
      patterns[216] = 12'b0_0_1_xxxxxxxx_x;
      patterns[217] = 12'b0_1_1_xxxxxxxx_x;
      patterns[218] = 12'b0_0_1_xxxxxxxx_0;
      patterns[219] = 12'b0_0_1_xxxxxxxx_x;
      patterns[220] = 12'b0_1_1_xxxxxxxx_x;
      patterns[221] = 12'b0_0_1_xxxxxxxx_0;
      patterns[222] = 12'b0_0_1_xxxxxxxx_x;
      patterns[223] = 12'b0_1_1_xxxxxxxx_x;
      patterns[224] = 12'b0_0_1_xxxxxxxx_0;
      patterns[225] = 12'b0_0_1_xxxxxxxx_x;
      patterns[226] = 12'b0_1_1_xxxxxxxx_x;
      patterns[227] = 12'b0_0_1_xxxxxxxx_0;
      patterns[228] = 12'b0_0_1_xxxxxxxx_x;
      patterns[229] = 12'b0_1_1_xxxxxxxx_x;
      patterns[230] = 12'b0_0_1_xxxxxxxx_0;
      patterns[231] = 12'b0_0_1_xxxxxxxx_x;
      patterns[232] = 12'b0_1_1_xxxxxxxx_x;
      patterns[233] = 12'b0_0_1_xxxxxxxx_0;
      patterns[234] = 12'b0_0_1_xxxxxxxx_x;
      patterns[235] = 12'b0_1_1_xxxxxxxx_x;
      patterns[236] = 12'b0_0_1_xxxxxxxx_0;
      patterns[237] = 12'b0_0_1_xxxxxxxx_x;
      patterns[238] = 12'b0_1_1_xxxxxxxx_x;
      patterns[239] = 12'b0_0_1_xxxxxxxx_0;
      patterns[240] = 12'b0_0_1_xxxxxxxx_x;
      patterns[241] = 12'b0_1_1_xxxxxxxx_x;
      patterns[242] = 12'b0_0_1_xxxxxxxx_0;
      patterns[243] = 12'b0_0_1_xxxxxxxx_x;
      patterns[244] = 12'b0_1_1_xxxxxxxx_x;
      patterns[245] = 12'b0_0_1_xxxxxxxx_0;
      patterns[246] = 12'b0_0_1_xxxxxxxx_x;
      patterns[247] = 12'b0_1_1_xxxxxxxx_x;
      patterns[248] = 12'b0_0_1_xxxxxxxx_0;
      patterns[249] = 12'b0_0_1_xxxxxxxx_x;
      patterns[250] = 12'b0_1_1_xxxxxxxx_x;
      patterns[251] = 12'b0_0_1_xxxxxxxx_0;
      patterns[252] = 12'b0_0_1_xxxxxxxx_x;
      patterns[253] = 12'b0_1_1_xxxxxxxx_x;
      patterns[254] = 12'b0_0_1_xxxxxxxx_0;
      patterns[255] = 12'b0_0_0_xxxxxxxx_x;
      patterns[256] = 12'b0_1_0_xxxxxxxx_x;
      patterns[257] = 12'b0_0_0_xxxxxxxx_0;
      patterns[258] = 12'b0_0_0_xxxxxxxx_x;
      patterns[259] = 12'b0_1_0_xxxxxxxx_x;
      patterns[260] = 12'b0_0_0_xxxxxxxx_0;
      patterns[261] = 12'b0_0_0_xxxxxxxx_x;
      patterns[262] = 12'b0_1_0_xxxxxxxx_x;
      patterns[263] = 12'b0_0_0_xxxxxxxx_0;
      patterns[264] = 12'b0_0_0_xxxxxxxx_x;
      patterns[265] = 12'b0_1_0_xxxxxxxx_x;
      patterns[266] = 12'b0_0_0_xxxxxxxx_0;
      patterns[267] = 12'b0_0_0_xxxxxxxx_x;
      patterns[268] = 12'b0_1_0_xxxxxxxx_x;
      patterns[269] = 12'b0_0_0_xxxxxxxx_0;
      patterns[270] = 12'b0_0_0_xxxxxxxx_x;
      patterns[271] = 12'b0_1_0_xxxxxxxx_x;
      patterns[272] = 12'b0_0_0_xxxxxxxx_0;
      patterns[273] = 12'b0_0_0_xxxxxxxx_x;
      patterns[274] = 12'b0_1_0_xxxxxxxx_x;
      patterns[275] = 12'b0_0_0_xxxxxxxx_0;
      patterns[276] = 12'b0_0_0_xxxxxxxx_x;
      patterns[277] = 12'b0_1_0_xxxxxxxx_x;
      patterns[278] = 12'b0_0_0_xxxxxxxx_0;
      patterns[279] = 12'b0_0_0_xxxxxxxx_x;
      patterns[280] = 12'b0_1_0_xxxxxxxx_x;
      patterns[281] = 12'b0_0_0_xxxxxxxx_0;
      patterns[282] = 12'b0_0_0_xxxxxxxx_x;
      patterns[283] = 12'b0_1_0_xxxxxxxx_x;
      patterns[284] = 12'b0_0_0_xxxxxxxx_0;
      patterns[285] = 12'b0_0_0_xxxxxxxx_x;
      patterns[286] = 12'b0_1_0_xxxxxxxx_x;
      patterns[287] = 12'b0_0_0_xxxxxxxx_0;
      patterns[288] = 12'b0_0_0_xxxxxxxx_x;
      patterns[289] = 12'b0_1_0_xxxxxxxx_x;
      patterns[290] = 12'b0_0_0_xxxxxxxx_0;
      patterns[291] = 12'b0_0_0_xxxxxxxx_x;
      patterns[292] = 12'b0_1_0_xxxxxxxx_x;
      patterns[293] = 12'b0_0_0_xxxxxxxx_0;
      patterns[294] = 12'b0_0_0_xxxxxxxx_x;
      patterns[295] = 12'b0_1_0_xxxxxxxx_x;
      patterns[296] = 12'b0_0_0_xxxxxxxx_0;
      patterns[297] = 12'b0_0_0_xxxxxxxx_x;
      patterns[298] = 12'b0_1_0_xxxxxxxx_x;
      patterns[299] = 12'b0_0_0_xxxxxxxx_0;
      patterns[300] = 12'b0_0_0_xxxxxxxx_x;
      patterns[301] = 12'b0_1_0_xxxxxxxx_x;
      patterns[302] = 12'b0_0_0_xxxxxxxx_0;
      patterns[303] = 12'b0_0_1_xxxxxxxx_x;
      patterns[304] = 12'b0_1_1_xxxxxxxx_x;
      patterns[305] = 12'b0_0_1_xxxxxxxx_0;
      patterns[306] = 12'b0_0_1_xxxxxxxx_x;
      patterns[307] = 12'b0_1_1_xxxxxxxx_x;
      patterns[308] = 12'b0_0_1_xxxxxxxx_0;
      patterns[309] = 12'b0_0_1_xxxxxxxx_x;
      patterns[310] = 12'b0_1_1_xxxxxxxx_x;
      patterns[311] = 12'b0_0_1_xxxxxxxx_0;
      patterns[312] = 12'b0_0_1_xxxxxxxx_x;
      patterns[313] = 12'b0_1_1_xxxxxxxx_x;
      patterns[314] = 12'b0_0_1_xxxxxxxx_0;
      patterns[315] = 12'b0_0_1_xxxxxxxx_x;
      patterns[316] = 12'b0_1_1_xxxxxxxx_x;
      patterns[317] = 12'b0_0_1_xxxxxxxx_0;
      patterns[318] = 12'b0_0_1_xxxxxxxx_x;
      patterns[319] = 12'b0_1_1_xxxxxxxx_x;
      patterns[320] = 12'b0_0_1_xxxxxxxx_0;
      patterns[321] = 12'b0_0_1_xxxxxxxx_x;
      patterns[322] = 12'b0_1_1_xxxxxxxx_x;
      patterns[323] = 12'b0_0_1_xxxxxxxx_0;
      patterns[324] = 12'b0_0_1_xxxxxxxx_x;
      patterns[325] = 12'b0_1_1_xxxxxxxx_x;
      patterns[326] = 12'b0_0_1_xxxxxxxx_0;
      patterns[327] = 12'b0_0_1_xxxxxxxx_x;
      patterns[328] = 12'b0_1_1_xxxxxxxx_x;
      patterns[329] = 12'b0_0_1_xxxxxxxx_0;
      patterns[330] = 12'b0_0_1_xxxxxxxx_x;
      patterns[331] = 12'b0_1_1_xxxxxxxx_x;
      patterns[332] = 12'b0_0_1_xxxxxxxx_0;
      patterns[333] = 12'b0_0_1_xxxxxxxx_x;
      patterns[334] = 12'b0_1_1_xxxxxxxx_x;
      patterns[335] = 12'b0_0_1_xxxxxxxx_0;
      patterns[336] = 12'b0_0_1_xxxxxxxx_x;
      patterns[337] = 12'b0_1_1_xxxxxxxx_x;
      patterns[338] = 12'b0_0_1_xxxxxxxx_0;
      patterns[339] = 12'b0_0_1_xxxxxxxx_x;
      patterns[340] = 12'b0_1_1_xxxxxxxx_x;
      patterns[341] = 12'b0_0_1_xxxxxxxx_0;
      patterns[342] = 12'b0_0_1_xxxxxxxx_x;
      patterns[343] = 12'b0_1_1_xxxxxxxx_x;
      patterns[344] = 12'b0_0_1_xxxxxxxx_0;
      patterns[345] = 12'b0_0_1_xxxxxxxx_x;
      patterns[346] = 12'b0_1_1_xxxxxxxx_x;
      patterns[347] = 12'b0_0_1_xxxxxxxx_0;
      patterns[348] = 12'b0_0_1_xxxxxxxx_x;
      patterns[349] = 12'b0_1_1_xxxxxxxx_x;
      patterns[350] = 12'b0_0_1_xxxxxxxx_0;
      patterns[351] = 12'b0_0_0_xxxxxxxx_x;
      patterns[352] = 12'b0_1_0_xxxxxxxx_x;
      patterns[353] = 12'b0_0_0_xxxxxxxx_0;
      patterns[354] = 12'b0_0_0_xxxxxxxx_x;
      patterns[355] = 12'b0_1_0_xxxxxxxx_x;
      patterns[356] = 12'b0_0_0_xxxxxxxx_0;
      patterns[357] = 12'b0_0_0_xxxxxxxx_x;
      patterns[358] = 12'b0_1_0_xxxxxxxx_x;
      patterns[359] = 12'b0_0_0_xxxxxxxx_0;
      patterns[360] = 12'b0_0_0_xxxxxxxx_x;
      patterns[361] = 12'b0_1_0_xxxxxxxx_x;
      patterns[362] = 12'b0_0_0_xxxxxxxx_0;
      patterns[363] = 12'b0_0_0_xxxxxxxx_x;
      patterns[364] = 12'b0_1_0_xxxxxxxx_x;
      patterns[365] = 12'b0_0_0_xxxxxxxx_0;
      patterns[366] = 12'b0_0_0_xxxxxxxx_x;
      patterns[367] = 12'b0_1_0_xxxxxxxx_x;
      patterns[368] = 12'b0_0_0_xxxxxxxx_0;
      patterns[369] = 12'b0_0_0_xxxxxxxx_x;
      patterns[370] = 12'b0_1_0_xxxxxxxx_x;
      patterns[371] = 12'b0_0_0_xxxxxxxx_0;
      patterns[372] = 12'b0_0_0_xxxxxxxx_x;
      patterns[373] = 12'b0_1_0_xxxxxxxx_x;
      patterns[374] = 12'b0_0_0_xxxxxxxx_0;
      patterns[375] = 12'b0_0_0_xxxxxxxx_x;
      patterns[376] = 12'b0_1_0_xxxxxxxx_x;
      patterns[377] = 12'b0_0_0_xxxxxxxx_0;
      patterns[378] = 12'b0_0_0_xxxxxxxx_x;
      patterns[379] = 12'b0_1_0_xxxxxxxx_x;
      patterns[380] = 12'b0_0_0_xxxxxxxx_0;
      patterns[381] = 12'b0_0_0_xxxxxxxx_x;
      patterns[382] = 12'b0_1_0_xxxxxxxx_x;
      patterns[383] = 12'b0_0_0_xxxxxxxx_0;
      patterns[384] = 12'b0_0_0_xxxxxxxx_x;
      patterns[385] = 12'b0_1_0_xxxxxxxx_x;
      patterns[386] = 12'b0_0_0_xxxxxxxx_0;
      patterns[387] = 12'b0_0_0_xxxxxxxx_x;
      patterns[388] = 12'b0_1_0_xxxxxxxx_x;
      patterns[389] = 12'b0_0_0_xxxxxxxx_0;
      patterns[390] = 12'b0_0_0_xxxxxxxx_x;
      patterns[391] = 12'b0_1_0_xxxxxxxx_x;
      patterns[392] = 12'b0_0_0_xxxxxxxx_0;
      patterns[393] = 12'b0_0_0_xxxxxxxx_x;
      patterns[394] = 12'b0_1_0_xxxxxxxx_x;
      patterns[395] = 12'b0_0_0_xxxxxxxx_0;
      patterns[396] = 12'b0_0_0_xxxxxxxx_x;
      patterns[397] = 12'b0_1_0_xxxxxxxx_x;
      patterns[398] = 12'b0_0_0_xxxxxxxx_0;
      patterns[399] = 12'b0_0_1_xxxxxxxx_x;
      patterns[400] = 12'b0_1_1_xxxxxxxx_x;
      patterns[401] = 12'b0_0_1_xxxxxxxx_x;
      patterns[402] = 12'b0_0_1_xxxxxxxx_x;
      patterns[403] = 12'b0_1_1_xxxxxxxx_x;
      patterns[404] = 12'b0_0_1_xxxxxxxx_x;
      patterns[405] = 12'b0_0_1_xxxxxxxx_x;
      patterns[406] = 12'b0_1_1_xxxxxxxx_x;
      patterns[407] = 12'b0_0_1_xxxxxxxx_x;
      patterns[408] = 12'b0_0_1_xxxxxxxx_x;
      patterns[409] = 12'b0_1_1_xxxxxxxx_x;
      patterns[410] = 12'b0_0_1_xxxxxxxx_x;
      patterns[411] = 12'b0_0_1_xxxxxxxx_x;
      patterns[412] = 12'b0_1_1_xxxxxxxx_x;
      patterns[413] = 12'b0_0_1_xxxxxxxx_x;
      patterns[414] = 12'b0_0_1_xxxxxxxx_x;
      patterns[415] = 12'b0_1_1_xxxxxxxx_x;
      patterns[416] = 12'b0_0_1_xxxxxxxx_x;
      patterns[417] = 12'b0_0_1_xxxxxxxx_x;
      patterns[418] = 12'b0_1_1_xxxxxxxx_x;
      patterns[419] = 12'b0_0_1_xxxxxxxx_x;
      patterns[420] = 12'b0_0_1_xxxxxxxx_x;
      patterns[421] = 12'b0_1_1_xxxxxxxx_x;
      patterns[422] = 12'b0_0_1_xxxxxxxx_x;
      patterns[423] = 12'b0_0_1_xxxxxxxx_x;
      patterns[424] = 12'b0_1_1_xxxxxxxx_x;
      patterns[425] = 12'b0_0_1_xxxxxxxx_x;
      patterns[426] = 12'b0_0_1_xxxxxxxx_x;
      patterns[427] = 12'b0_1_1_xxxxxxxx_x;
      patterns[428] = 12'b0_0_1_xxxxxxxx_x;
      patterns[429] = 12'b0_0_1_xxxxxxxx_x;
      patterns[430] = 12'b0_1_1_xxxxxxxx_x;
      patterns[431] = 12'b0_0_1_xxxxxxxx_x;
      patterns[432] = 12'b0_0_1_xxxxxxxx_x;
      patterns[433] = 12'b0_1_1_xxxxxxxx_x;
      patterns[434] = 12'b0_0_1_xxxxxxxx_x;
      patterns[435] = 12'b0_0_1_xxxxxxxx_x;
      patterns[436] = 12'b0_1_1_xxxxxxxx_x;
      patterns[437] = 12'b0_0_1_xxxxxxxx_x;
      patterns[438] = 12'b0_0_1_xxxxxxxx_x;
      patterns[439] = 12'b0_1_1_xxxxxxxx_x;
      patterns[440] = 12'b0_0_1_xxxxxxxx_x;
      patterns[441] = 12'b0_0_1_xxxxxxxx_x;
      patterns[442] = 12'b0_1_1_xxxxxxxx_x;
      patterns[443] = 12'b0_0_1_xxxxxxxx_x;
      patterns[444] = 12'b0_0_1_xxxxxxxx_x;
      patterns[445] = 12'b0_1_1_xxxxxxxx_x;
      patterns[446] = 12'b0_0_1_xxxxxxxx_x;
      patterns[447] = 12'b0_0_0_xxxxxxxx_x;
      patterns[448] = 12'b0_1_0_xxxxxxxx_x;
      patterns[449] = 12'b0_0_0_10101010_1;
      patterns[450] = 12'b0_0_0_xxxxxxxx_x;
      patterns[451] = 12'b0_1_0_xxxxxxxx_x;
      patterns[452] = 12'b0_0_0_10101010_1;
      patterns[453] = 12'b0_0_0_xxxxxxxx_x;
      patterns[454] = 12'b0_1_0_xxxxxxxx_x;
      patterns[455] = 12'b0_0_0_10101010_1;
      patterns[456] = 12'b0_0_0_xxxxxxxx_x;
      patterns[457] = 12'b0_1_0_xxxxxxxx_x;
      patterns[458] = 12'b0_0_0_10101010_1;
      patterns[459] = 12'b0_0_0_xxxxxxxx_x;
      patterns[460] = 12'b0_1_0_xxxxxxxx_x;
      patterns[461] = 12'b0_0_0_10101010_1;
      patterns[462] = 12'b0_0_0_xxxxxxxx_x;
      patterns[463] = 12'b0_1_0_xxxxxxxx_x;
      patterns[464] = 12'b0_0_0_10101010_1;
      patterns[465] = 12'b0_0_0_xxxxxxxx_x;
      patterns[466] = 12'b0_1_0_xxxxxxxx_x;
      patterns[467] = 12'b0_0_0_10101010_1;
      patterns[468] = 12'b0_0_0_xxxxxxxx_x;
      patterns[469] = 12'b0_1_0_xxxxxxxx_x;
      patterns[470] = 12'b0_0_0_10101010_1;
      patterns[471] = 12'b0_0_0_xxxxxxxx_x;
      patterns[472] = 12'b0_1_0_xxxxxxxx_x;
      patterns[473] = 12'b0_0_0_10101010_1;
      patterns[474] = 12'b0_0_0_xxxxxxxx_x;
      patterns[475] = 12'b0_1_0_xxxxxxxx_x;
      patterns[476] = 12'b0_0_0_10101010_1;
      patterns[477] = 12'b0_0_0_xxxxxxxx_x;
      patterns[478] = 12'b0_1_0_xxxxxxxx_x;
      patterns[479] = 12'b0_0_0_10101010_1;
      patterns[480] = 12'b0_0_0_xxxxxxxx_x;
      patterns[481] = 12'b0_1_0_xxxxxxxx_x;
      patterns[482] = 12'b0_0_0_10101010_1;
      patterns[483] = 12'b0_0_0_xxxxxxxx_x;
      patterns[484] = 12'b0_1_0_xxxxxxxx_x;
      patterns[485] = 12'b0_0_0_10101010_1;
      patterns[486] = 12'b0_0_0_xxxxxxxx_x;
      patterns[487] = 12'b0_1_0_xxxxxxxx_x;
      patterns[488] = 12'b0_0_0_10101010_1;
      patterns[489] = 12'b0_0_0_xxxxxxxx_x;
      patterns[490] = 12'b0_1_0_xxxxxxxx_x;
      patterns[491] = 12'b0_0_0_10101010_1;
      patterns[492] = 12'b0_0_0_xxxxxxxx_x;
      patterns[493] = 12'b0_1_0_xxxxxxxx_x;
      patterns[494] = 12'b0_0_0_10101010_1;
      patterns[495] = 12'b1_0_0_xxxxxxxx_x;
      patterns[496] = 12'b1_1_0_xxxxxxxx_x;
      patterns[497] = 12'b1_0_0_xxxxxxxx_0;
      patterns[498] = 12'b0_0_0_xxxxxxxx_x;
      patterns[499] = 12'b0_1_0_xxxxxxxx_x;
      patterns[500] = 12'b0_0_0_xxxxxxxx_0;
      patterns[501] = 12'b0_0_0_xxxxxxxx_x;
      patterns[502] = 12'b0_1_0_xxxxxxxx_x;
      patterns[503] = 12'b0_0_0_xxxxxxxx_0;
      patterns[504] = 12'b0_0_0_xxxxxxxx_x;
      patterns[505] = 12'b0_1_0_xxxxxxxx_x;
      patterns[506] = 12'b0_0_0_xxxxxxxx_0;
      patterns[507] = 12'b0_0_0_xxxxxxxx_x;
      patterns[508] = 12'b0_1_0_xxxxxxxx_x;
      patterns[509] = 12'b0_0_0_xxxxxxxx_0;
      patterns[510] = 12'b0_0_0_xxxxxxxx_x;
      patterns[511] = 12'b0_1_0_xxxxxxxx_x;
      patterns[512] = 12'b0_0_0_xxxxxxxx_0;
      patterns[513] = 12'b0_0_1_xxxxxxxx_x;
      patterns[514] = 12'b0_1_1_xxxxxxxx_x;
      patterns[515] = 12'b0_0_1_xxxxxxxx_0;
      patterns[516] = 12'b0_0_1_xxxxxxxx_x;
      patterns[517] = 12'b0_1_1_xxxxxxxx_x;
      patterns[518] = 12'b0_0_1_xxxxxxxx_0;
      patterns[519] = 12'b0_0_1_xxxxxxxx_x;
      patterns[520] = 12'b0_1_1_xxxxxxxx_x;
      patterns[521] = 12'b0_0_1_xxxxxxxx_0;
      patterns[522] = 12'b0_0_1_xxxxxxxx_x;
      patterns[523] = 12'b0_1_1_xxxxxxxx_x;
      patterns[524] = 12'b0_0_1_xxxxxxxx_0;
      patterns[525] = 12'b0_0_1_xxxxxxxx_x;
      patterns[526] = 12'b0_1_1_xxxxxxxx_x;
      patterns[527] = 12'b0_0_1_xxxxxxxx_0;
      patterns[528] = 12'b0_0_1_xxxxxxxx_x;
      patterns[529] = 12'b0_1_1_xxxxxxxx_x;
      patterns[530] = 12'b0_0_1_xxxxxxxx_0;
      patterns[531] = 12'b0_0_1_xxxxxxxx_x;
      patterns[532] = 12'b0_1_1_xxxxxxxx_x;
      patterns[533] = 12'b0_0_1_xxxxxxxx_0;
      patterns[534] = 12'b0_0_1_xxxxxxxx_x;
      patterns[535] = 12'b0_1_1_xxxxxxxx_x;
      patterns[536] = 12'b0_0_1_xxxxxxxx_0;
      patterns[537] = 12'b0_0_1_xxxxxxxx_x;
      patterns[538] = 12'b0_1_1_xxxxxxxx_x;
      patterns[539] = 12'b0_0_1_xxxxxxxx_0;
      patterns[540] = 12'b0_0_1_xxxxxxxx_x;
      patterns[541] = 12'b0_1_1_xxxxxxxx_x;
      patterns[542] = 12'b0_0_1_xxxxxxxx_0;
      patterns[543] = 12'b0_0_1_xxxxxxxx_x;
      patterns[544] = 12'b0_1_1_xxxxxxxx_x;
      patterns[545] = 12'b0_0_1_xxxxxxxx_0;
      patterns[546] = 12'b0_0_1_xxxxxxxx_x;
      patterns[547] = 12'b0_1_1_xxxxxxxx_x;
      patterns[548] = 12'b0_0_1_xxxxxxxx_0;
      patterns[549] = 12'b0_0_1_xxxxxxxx_x;
      patterns[550] = 12'b0_1_1_xxxxxxxx_x;
      patterns[551] = 12'b0_0_1_xxxxxxxx_0;
      patterns[552] = 12'b0_0_1_xxxxxxxx_x;
      patterns[553] = 12'b0_1_1_xxxxxxxx_x;
      patterns[554] = 12'b0_0_1_xxxxxxxx_0;
      patterns[555] = 12'b0_0_1_xxxxxxxx_x;
      patterns[556] = 12'b0_1_1_xxxxxxxx_x;
      patterns[557] = 12'b0_0_1_xxxxxxxx_0;
      patterns[558] = 12'b0_0_1_xxxxxxxx_x;
      patterns[559] = 12'b0_1_1_xxxxxxxx_x;
      patterns[560] = 12'b0_0_1_xxxxxxxx_0;
      patterns[561] = 12'b0_0_1_xxxxxxxx_x;
      patterns[562] = 12'b0_1_1_xxxxxxxx_x;
      patterns[563] = 12'b0_0_1_xxxxxxxx_0;
      patterns[564] = 12'b0_0_1_xxxxxxxx_x;
      patterns[565] = 12'b0_1_1_xxxxxxxx_x;
      patterns[566] = 12'b0_0_1_xxxxxxxx_0;
      patterns[567] = 12'b0_0_1_xxxxxxxx_x;
      patterns[568] = 12'b0_1_1_xxxxxxxx_x;
      patterns[569] = 12'b0_0_1_xxxxxxxx_0;
      patterns[570] = 12'b0_0_1_xxxxxxxx_x;
      patterns[571] = 12'b0_1_1_xxxxxxxx_x;
      patterns[572] = 12'b0_0_1_xxxxxxxx_0;
      patterns[573] = 12'b0_0_1_xxxxxxxx_x;
      patterns[574] = 12'b0_1_1_xxxxxxxx_x;
      patterns[575] = 12'b0_0_1_xxxxxxxx_0;
      patterns[576] = 12'b0_0_1_xxxxxxxx_x;
      patterns[577] = 12'b0_1_1_xxxxxxxx_x;
      patterns[578] = 12'b0_0_1_xxxxxxxx_0;
      patterns[579] = 12'b0_0_1_xxxxxxxx_x;
      patterns[580] = 12'b0_1_1_xxxxxxxx_x;
      patterns[581] = 12'b0_0_1_xxxxxxxx_0;
      patterns[582] = 12'b0_0_1_xxxxxxxx_x;
      patterns[583] = 12'b0_1_1_xxxxxxxx_x;
      patterns[584] = 12'b0_0_1_xxxxxxxx_0;
      patterns[585] = 12'b0_0_1_xxxxxxxx_x;
      patterns[586] = 12'b0_1_1_xxxxxxxx_x;
      patterns[587] = 12'b0_0_1_xxxxxxxx_0;
      patterns[588] = 12'b0_0_1_xxxxxxxx_x;
      patterns[589] = 12'b0_1_1_xxxxxxxx_x;
      patterns[590] = 12'b0_0_1_xxxxxxxx_0;
      patterns[591] = 12'b0_0_1_xxxxxxxx_x;
      patterns[592] = 12'b0_1_1_xxxxxxxx_x;
      patterns[593] = 12'b0_0_1_xxxxxxxx_0;
      patterns[594] = 12'b0_0_1_xxxxxxxx_x;
      patterns[595] = 12'b0_1_1_xxxxxxxx_x;
      patterns[596] = 12'b0_0_1_xxxxxxxx_0;
      patterns[597] = 12'b0_0_1_xxxxxxxx_x;
      patterns[598] = 12'b0_1_1_xxxxxxxx_x;
      patterns[599] = 12'b0_0_1_xxxxxxxx_0;
      patterns[600] = 12'b0_0_1_xxxxxxxx_x;
      patterns[601] = 12'b0_1_1_xxxxxxxx_x;
      patterns[602] = 12'b0_0_1_xxxxxxxx_0;
      patterns[603] = 12'b0_0_1_xxxxxxxx_x;
      patterns[604] = 12'b0_1_1_xxxxxxxx_x;
      patterns[605] = 12'b0_0_1_xxxxxxxx_0;
      patterns[606] = 12'b0_0_1_xxxxxxxx_x;
      patterns[607] = 12'b0_1_1_xxxxxxxx_x;
      patterns[608] = 12'b0_0_1_xxxxxxxx_0;
      patterns[609] = 12'b0_0_0_xxxxxxxx_x;
      patterns[610] = 12'b0_1_0_xxxxxxxx_x;
      patterns[611] = 12'b0_0_0_xxxxxxxx_0;
      patterns[612] = 12'b0_0_0_xxxxxxxx_x;
      patterns[613] = 12'b0_1_0_xxxxxxxx_x;
      patterns[614] = 12'b0_0_0_xxxxxxxx_0;
      patterns[615] = 12'b0_0_0_xxxxxxxx_x;
      patterns[616] = 12'b0_1_0_xxxxxxxx_x;
      patterns[617] = 12'b0_0_0_xxxxxxxx_0;
      patterns[618] = 12'b0_0_0_xxxxxxxx_x;
      patterns[619] = 12'b0_1_0_xxxxxxxx_x;
      patterns[620] = 12'b0_0_0_xxxxxxxx_0;
      patterns[621] = 12'b0_0_0_xxxxxxxx_x;
      patterns[622] = 12'b0_1_0_xxxxxxxx_x;
      patterns[623] = 12'b0_0_0_xxxxxxxx_0;
      patterns[624] = 12'b0_0_0_xxxxxxxx_x;
      patterns[625] = 12'b0_1_0_xxxxxxxx_x;
      patterns[626] = 12'b0_0_0_xxxxxxxx_0;
      patterns[627] = 12'b0_0_0_xxxxxxxx_x;
      patterns[628] = 12'b0_1_0_xxxxxxxx_x;
      patterns[629] = 12'b0_0_0_xxxxxxxx_0;
      patterns[630] = 12'b0_0_0_xxxxxxxx_x;
      patterns[631] = 12'b0_1_0_xxxxxxxx_x;
      patterns[632] = 12'b0_0_0_xxxxxxxx_0;
      patterns[633] = 12'b0_0_0_xxxxxxxx_x;
      patterns[634] = 12'b0_1_0_xxxxxxxx_x;
      patterns[635] = 12'b0_0_0_xxxxxxxx_0;
      patterns[636] = 12'b0_0_0_xxxxxxxx_x;
      patterns[637] = 12'b0_1_0_xxxxxxxx_x;
      patterns[638] = 12'b0_0_0_xxxxxxxx_0;
      patterns[639] = 12'b0_0_0_xxxxxxxx_x;
      patterns[640] = 12'b0_1_0_xxxxxxxx_x;
      patterns[641] = 12'b0_0_0_xxxxxxxx_0;
      patterns[642] = 12'b0_0_0_xxxxxxxx_x;
      patterns[643] = 12'b0_1_0_xxxxxxxx_x;
      patterns[644] = 12'b0_0_0_xxxxxxxx_0;
      patterns[645] = 12'b0_0_0_xxxxxxxx_x;
      patterns[646] = 12'b0_1_0_xxxxxxxx_x;
      patterns[647] = 12'b0_0_0_xxxxxxxx_0;
      patterns[648] = 12'b0_0_0_xxxxxxxx_x;
      patterns[649] = 12'b0_1_0_xxxxxxxx_x;
      patterns[650] = 12'b0_0_0_xxxxxxxx_0;
      patterns[651] = 12'b0_0_0_xxxxxxxx_x;
      patterns[652] = 12'b0_1_0_xxxxxxxx_x;
      patterns[653] = 12'b0_0_0_xxxxxxxx_0;
      patterns[654] = 12'b0_0_0_xxxxxxxx_x;
      patterns[655] = 12'b0_1_0_xxxxxxxx_x;
      patterns[656] = 12'b0_0_0_xxxxxxxx_0;
      patterns[657] = 12'b0_0_1_xxxxxxxx_x;
      patterns[658] = 12'b0_1_1_xxxxxxxx_x;
      patterns[659] = 12'b0_0_1_xxxxxxxx_0;
      patterns[660] = 12'b0_0_1_xxxxxxxx_x;
      patterns[661] = 12'b0_1_1_xxxxxxxx_x;
      patterns[662] = 12'b0_0_1_xxxxxxxx_0;
      patterns[663] = 12'b0_0_1_xxxxxxxx_x;
      patterns[664] = 12'b0_1_1_xxxxxxxx_x;
      patterns[665] = 12'b0_0_1_xxxxxxxx_0;
      patterns[666] = 12'b0_0_1_xxxxxxxx_x;
      patterns[667] = 12'b0_1_1_xxxxxxxx_x;
      patterns[668] = 12'b0_0_1_xxxxxxxx_0;
      patterns[669] = 12'b0_0_1_xxxxxxxx_x;
      patterns[670] = 12'b0_1_1_xxxxxxxx_x;
      patterns[671] = 12'b0_0_1_xxxxxxxx_0;
      patterns[672] = 12'b0_0_1_xxxxxxxx_x;
      patterns[673] = 12'b0_1_1_xxxxxxxx_x;
      patterns[674] = 12'b0_0_1_xxxxxxxx_0;
      patterns[675] = 12'b0_0_1_xxxxxxxx_x;
      patterns[676] = 12'b0_1_1_xxxxxxxx_x;
      patterns[677] = 12'b0_0_1_xxxxxxxx_0;
      patterns[678] = 12'b0_0_1_xxxxxxxx_x;
      patterns[679] = 12'b0_1_1_xxxxxxxx_x;
      patterns[680] = 12'b0_0_1_xxxxxxxx_0;
      patterns[681] = 12'b0_0_1_xxxxxxxx_x;
      patterns[682] = 12'b0_1_1_xxxxxxxx_x;
      patterns[683] = 12'b0_0_1_xxxxxxxx_0;
      patterns[684] = 12'b0_0_1_xxxxxxxx_x;
      patterns[685] = 12'b0_1_1_xxxxxxxx_x;
      patterns[686] = 12'b0_0_1_xxxxxxxx_0;
      patterns[687] = 12'b0_0_1_xxxxxxxx_x;
      patterns[688] = 12'b0_1_1_xxxxxxxx_x;
      patterns[689] = 12'b0_0_1_xxxxxxxx_0;
      patterns[690] = 12'b0_0_1_xxxxxxxx_x;
      patterns[691] = 12'b0_1_1_xxxxxxxx_x;
      patterns[692] = 12'b0_0_1_xxxxxxxx_0;
      patterns[693] = 12'b0_0_1_xxxxxxxx_x;
      patterns[694] = 12'b0_1_1_xxxxxxxx_x;
      patterns[695] = 12'b0_0_1_xxxxxxxx_0;
      patterns[696] = 12'b0_0_1_xxxxxxxx_x;
      patterns[697] = 12'b0_1_1_xxxxxxxx_x;
      patterns[698] = 12'b0_0_1_xxxxxxxx_0;
      patterns[699] = 12'b0_0_1_xxxxxxxx_x;
      patterns[700] = 12'b0_1_1_xxxxxxxx_x;
      patterns[701] = 12'b0_0_1_xxxxxxxx_0;
      patterns[702] = 12'b0_0_1_xxxxxxxx_x;
      patterns[703] = 12'b0_1_1_xxxxxxxx_x;
      patterns[704] = 12'b0_0_1_xxxxxxxx_0;
      patterns[705] = 12'b0_0_0_xxxxxxxx_x;
      patterns[706] = 12'b0_1_0_xxxxxxxx_x;
      patterns[707] = 12'b0_0_0_xxxxxxxx_0;
      patterns[708] = 12'b0_0_0_xxxxxxxx_x;
      patterns[709] = 12'b0_1_0_xxxxxxxx_x;
      patterns[710] = 12'b0_0_0_xxxxxxxx_0;
      patterns[711] = 12'b0_0_0_xxxxxxxx_x;
      patterns[712] = 12'b0_1_0_xxxxxxxx_x;
      patterns[713] = 12'b0_0_0_xxxxxxxx_0;
      patterns[714] = 12'b0_0_0_xxxxxxxx_x;
      patterns[715] = 12'b0_1_0_xxxxxxxx_x;
      patterns[716] = 12'b0_0_0_xxxxxxxx_0;
      patterns[717] = 12'b0_0_0_xxxxxxxx_x;
      patterns[718] = 12'b0_1_0_xxxxxxxx_x;
      patterns[719] = 12'b0_0_0_xxxxxxxx_0;
      patterns[720] = 12'b0_0_0_xxxxxxxx_x;
      patterns[721] = 12'b0_1_0_xxxxxxxx_x;
      patterns[722] = 12'b0_0_0_xxxxxxxx_0;
      patterns[723] = 12'b0_0_0_xxxxxxxx_x;
      patterns[724] = 12'b0_1_0_xxxxxxxx_x;
      patterns[725] = 12'b0_0_0_xxxxxxxx_0;
      patterns[726] = 12'b0_0_0_xxxxxxxx_x;
      patterns[727] = 12'b0_1_0_xxxxxxxx_x;
      patterns[728] = 12'b0_0_0_xxxxxxxx_0;
      patterns[729] = 12'b0_0_0_xxxxxxxx_x;
      patterns[730] = 12'b0_1_0_xxxxxxxx_x;
      patterns[731] = 12'b0_0_0_xxxxxxxx_0;
      patterns[732] = 12'b0_0_0_xxxxxxxx_x;
      patterns[733] = 12'b0_1_0_xxxxxxxx_x;
      patterns[734] = 12'b0_0_0_xxxxxxxx_0;
      patterns[735] = 12'b0_0_0_xxxxxxxx_x;
      patterns[736] = 12'b0_1_0_xxxxxxxx_x;
      patterns[737] = 12'b0_0_0_xxxxxxxx_0;
      patterns[738] = 12'b0_0_0_xxxxxxxx_x;
      patterns[739] = 12'b0_1_0_xxxxxxxx_x;
      patterns[740] = 12'b0_0_0_xxxxxxxx_0;
      patterns[741] = 12'b0_0_0_xxxxxxxx_x;
      patterns[742] = 12'b0_1_0_xxxxxxxx_x;
      patterns[743] = 12'b0_0_0_xxxxxxxx_0;
      patterns[744] = 12'b0_0_0_xxxxxxxx_x;
      patterns[745] = 12'b0_1_0_xxxxxxxx_x;
      patterns[746] = 12'b0_0_0_xxxxxxxx_0;
      patterns[747] = 12'b0_0_0_xxxxxxxx_x;
      patterns[748] = 12'b0_1_0_xxxxxxxx_x;
      patterns[749] = 12'b0_0_0_xxxxxxxx_0;
      patterns[750] = 12'b0_0_0_xxxxxxxx_x;
      patterns[751] = 12'b0_1_0_xxxxxxxx_x;
      patterns[752] = 12'b0_0_0_xxxxxxxx_0;
      patterns[753] = 12'b0_0_1_xxxxxxxx_x;
      patterns[754] = 12'b0_1_1_xxxxxxxx_x;
      patterns[755] = 12'b0_0_1_xxxxxxxx_0;
      patterns[756] = 12'b0_0_1_xxxxxxxx_x;
      patterns[757] = 12'b0_1_1_xxxxxxxx_x;
      patterns[758] = 12'b0_0_1_xxxxxxxx_0;
      patterns[759] = 12'b0_0_1_xxxxxxxx_x;
      patterns[760] = 12'b0_1_1_xxxxxxxx_x;
      patterns[761] = 12'b0_0_1_xxxxxxxx_0;
      patterns[762] = 12'b0_0_1_xxxxxxxx_x;
      patterns[763] = 12'b0_1_1_xxxxxxxx_x;
      patterns[764] = 12'b0_0_1_xxxxxxxx_0;
      patterns[765] = 12'b0_0_1_xxxxxxxx_x;
      patterns[766] = 12'b0_1_1_xxxxxxxx_x;
      patterns[767] = 12'b0_0_1_xxxxxxxx_0;
      patterns[768] = 12'b0_0_1_xxxxxxxx_x;
      patterns[769] = 12'b0_1_1_xxxxxxxx_x;
      patterns[770] = 12'b0_0_1_xxxxxxxx_0;
      patterns[771] = 12'b0_0_1_xxxxxxxx_x;
      patterns[772] = 12'b0_1_1_xxxxxxxx_x;
      patterns[773] = 12'b0_0_1_xxxxxxxx_0;
      patterns[774] = 12'b0_0_1_xxxxxxxx_x;
      patterns[775] = 12'b0_1_1_xxxxxxxx_x;
      patterns[776] = 12'b0_0_1_xxxxxxxx_0;
      patterns[777] = 12'b0_0_1_xxxxxxxx_x;
      patterns[778] = 12'b0_1_1_xxxxxxxx_x;
      patterns[779] = 12'b0_0_1_xxxxxxxx_0;
      patterns[780] = 12'b0_0_1_xxxxxxxx_x;
      patterns[781] = 12'b0_1_1_xxxxxxxx_x;
      patterns[782] = 12'b0_0_1_xxxxxxxx_0;
      patterns[783] = 12'b0_0_1_xxxxxxxx_x;
      patterns[784] = 12'b0_1_1_xxxxxxxx_x;
      patterns[785] = 12'b0_0_1_xxxxxxxx_0;
      patterns[786] = 12'b0_0_1_xxxxxxxx_x;
      patterns[787] = 12'b0_1_1_xxxxxxxx_x;
      patterns[788] = 12'b0_0_1_xxxxxxxx_0;
      patterns[789] = 12'b0_0_1_xxxxxxxx_x;
      patterns[790] = 12'b0_1_1_xxxxxxxx_x;
      patterns[791] = 12'b0_0_1_xxxxxxxx_0;
      patterns[792] = 12'b0_0_1_xxxxxxxx_x;
      patterns[793] = 12'b0_1_1_xxxxxxxx_x;
      patterns[794] = 12'b0_0_1_xxxxxxxx_0;
      patterns[795] = 12'b0_0_1_xxxxxxxx_x;
      patterns[796] = 12'b0_1_1_xxxxxxxx_x;
      patterns[797] = 12'b0_0_1_xxxxxxxx_0;
      patterns[798] = 12'b0_0_1_xxxxxxxx_x;
      patterns[799] = 12'b0_1_1_xxxxxxxx_x;
      patterns[800] = 12'b0_0_1_xxxxxxxx_0;
      patterns[801] = 12'b0_0_0_xxxxxxxx_x;
      patterns[802] = 12'b0_1_0_xxxxxxxx_x;
      patterns[803] = 12'b0_0_0_xxxxxxxx_0;
      patterns[804] = 12'b0_0_0_xxxxxxxx_x;
      patterns[805] = 12'b0_1_0_xxxxxxxx_x;
      patterns[806] = 12'b0_0_0_xxxxxxxx_0;
      patterns[807] = 12'b0_0_0_xxxxxxxx_x;
      patterns[808] = 12'b0_1_0_xxxxxxxx_x;
      patterns[809] = 12'b0_0_0_xxxxxxxx_0;
      patterns[810] = 12'b0_0_0_xxxxxxxx_x;
      patterns[811] = 12'b0_1_0_xxxxxxxx_x;
      patterns[812] = 12'b0_0_0_xxxxxxxx_0;
      patterns[813] = 12'b0_0_0_xxxxxxxx_x;
      patterns[814] = 12'b0_1_0_xxxxxxxx_x;
      patterns[815] = 12'b0_0_0_xxxxxxxx_0;
      patterns[816] = 12'b0_0_0_xxxxxxxx_x;
      patterns[817] = 12'b0_1_0_xxxxxxxx_x;
      patterns[818] = 12'b0_0_0_xxxxxxxx_0;
      patterns[819] = 12'b0_0_0_xxxxxxxx_x;
      patterns[820] = 12'b0_1_0_xxxxxxxx_x;
      patterns[821] = 12'b0_0_0_xxxxxxxx_0;
      patterns[822] = 12'b0_0_0_xxxxxxxx_x;
      patterns[823] = 12'b0_1_0_xxxxxxxx_x;
      patterns[824] = 12'b0_0_0_xxxxxxxx_0;
      patterns[825] = 12'b0_0_0_xxxxxxxx_x;
      patterns[826] = 12'b0_1_0_xxxxxxxx_x;
      patterns[827] = 12'b0_0_0_xxxxxxxx_0;
      patterns[828] = 12'b0_0_0_xxxxxxxx_x;
      patterns[829] = 12'b0_1_0_xxxxxxxx_x;
      patterns[830] = 12'b0_0_0_xxxxxxxx_0;
      patterns[831] = 12'b0_0_0_xxxxxxxx_x;
      patterns[832] = 12'b0_1_0_xxxxxxxx_x;
      patterns[833] = 12'b0_0_0_xxxxxxxx_0;
      patterns[834] = 12'b0_0_0_xxxxxxxx_x;
      patterns[835] = 12'b0_1_0_xxxxxxxx_x;
      patterns[836] = 12'b0_0_0_xxxxxxxx_0;
      patterns[837] = 12'b0_0_0_xxxxxxxx_x;
      patterns[838] = 12'b0_1_0_xxxxxxxx_x;
      patterns[839] = 12'b0_0_0_xxxxxxxx_0;
      patterns[840] = 12'b0_0_0_xxxxxxxx_x;
      patterns[841] = 12'b0_1_0_xxxxxxxx_x;
      patterns[842] = 12'b0_0_0_xxxxxxxx_0;
      patterns[843] = 12'b0_0_0_xxxxxxxx_x;
      patterns[844] = 12'b0_1_0_xxxxxxxx_x;
      patterns[845] = 12'b0_0_0_xxxxxxxx_0;
      patterns[846] = 12'b0_0_0_xxxxxxxx_x;
      patterns[847] = 12'b0_1_0_xxxxxxxx_x;
      patterns[848] = 12'b0_0_0_xxxxxxxx_0;
      patterns[849] = 12'b0_0_1_xxxxxxxx_x;
      patterns[850] = 12'b0_1_1_xxxxxxxx_x;
      patterns[851] = 12'b0_0_1_xxxxxxxx_0;
      patterns[852] = 12'b0_0_1_xxxxxxxx_x;
      patterns[853] = 12'b0_1_1_xxxxxxxx_x;
      patterns[854] = 12'b0_0_1_xxxxxxxx_0;
      patterns[855] = 12'b0_0_1_xxxxxxxx_x;
      patterns[856] = 12'b0_1_1_xxxxxxxx_x;
      patterns[857] = 12'b0_0_1_xxxxxxxx_0;
      patterns[858] = 12'b0_0_1_xxxxxxxx_x;
      patterns[859] = 12'b0_1_1_xxxxxxxx_x;
      patterns[860] = 12'b0_0_1_xxxxxxxx_0;
      patterns[861] = 12'b0_0_1_xxxxxxxx_x;
      patterns[862] = 12'b0_1_1_xxxxxxxx_x;
      patterns[863] = 12'b0_0_1_xxxxxxxx_0;
      patterns[864] = 12'b0_0_1_xxxxxxxx_x;
      patterns[865] = 12'b0_1_1_xxxxxxxx_x;
      patterns[866] = 12'b0_0_1_xxxxxxxx_0;
      patterns[867] = 12'b0_0_1_xxxxxxxx_x;
      patterns[868] = 12'b0_1_1_xxxxxxxx_x;
      patterns[869] = 12'b0_0_1_xxxxxxxx_0;
      patterns[870] = 12'b0_0_1_xxxxxxxx_x;
      patterns[871] = 12'b0_1_1_xxxxxxxx_x;
      patterns[872] = 12'b0_0_1_xxxxxxxx_0;
      patterns[873] = 12'b0_0_1_xxxxxxxx_x;
      patterns[874] = 12'b0_1_1_xxxxxxxx_x;
      patterns[875] = 12'b0_0_1_xxxxxxxx_0;
      patterns[876] = 12'b0_0_1_xxxxxxxx_x;
      patterns[877] = 12'b0_1_1_xxxxxxxx_x;
      patterns[878] = 12'b0_0_1_xxxxxxxx_0;
      patterns[879] = 12'b0_0_1_xxxxxxxx_x;
      patterns[880] = 12'b0_1_1_xxxxxxxx_x;
      patterns[881] = 12'b0_0_1_xxxxxxxx_0;
      patterns[882] = 12'b0_0_1_xxxxxxxx_x;
      patterns[883] = 12'b0_1_1_xxxxxxxx_x;
      patterns[884] = 12'b0_0_1_xxxxxxxx_0;
      patterns[885] = 12'b0_0_1_xxxxxxxx_x;
      patterns[886] = 12'b0_1_1_xxxxxxxx_x;
      patterns[887] = 12'b0_0_1_xxxxxxxx_0;
      patterns[888] = 12'b0_0_1_xxxxxxxx_x;
      patterns[889] = 12'b0_1_1_xxxxxxxx_x;
      patterns[890] = 12'b0_0_1_xxxxxxxx_0;
      patterns[891] = 12'b0_0_1_xxxxxxxx_x;
      patterns[892] = 12'b0_1_1_xxxxxxxx_x;
      patterns[893] = 12'b0_0_1_xxxxxxxx_0;
      patterns[894] = 12'b0_0_1_xxxxxxxx_x;
      patterns[895] = 12'b0_1_1_xxxxxxxx_x;
      patterns[896] = 12'b0_0_1_xxxxxxxx_0;
      patterns[897] = 12'b0_0_0_xxxxxxxx_x;
      patterns[898] = 12'b0_1_0_xxxxxxxx_x;
      patterns[899] = 12'b0_0_0_xxxxxxxx_x;
      patterns[900] = 12'b0_0_0_xxxxxxxx_x;
      patterns[901] = 12'b0_1_0_xxxxxxxx_x;
      patterns[902] = 12'b0_0_0_xxxxxxxx_x;
      patterns[903] = 12'b0_0_0_xxxxxxxx_x;
      patterns[904] = 12'b0_1_0_xxxxxxxx_x;
      patterns[905] = 12'b0_0_0_xxxxxxxx_x;
      patterns[906] = 12'b0_0_0_xxxxxxxx_x;
      patterns[907] = 12'b0_1_0_xxxxxxxx_x;
      patterns[908] = 12'b0_0_0_xxxxxxxx_x;
      patterns[909] = 12'b0_0_0_xxxxxxxx_x;
      patterns[910] = 12'b0_1_0_xxxxxxxx_x;
      patterns[911] = 12'b0_0_0_xxxxxxxx_x;
      patterns[912] = 12'b0_0_0_xxxxxxxx_x;
      patterns[913] = 12'b0_1_0_xxxxxxxx_x;
      patterns[914] = 12'b0_0_0_xxxxxxxx_x;
      patterns[915] = 12'b0_0_0_xxxxxxxx_x;
      patterns[916] = 12'b0_1_0_xxxxxxxx_x;
      patterns[917] = 12'b0_0_0_xxxxxxxx_x;
      patterns[918] = 12'b0_0_0_xxxxxxxx_x;
      patterns[919] = 12'b0_1_0_xxxxxxxx_x;
      patterns[920] = 12'b0_0_0_xxxxxxxx_x;
      patterns[921] = 12'b0_0_0_xxxxxxxx_x;
      patterns[922] = 12'b0_1_0_xxxxxxxx_x;
      patterns[923] = 12'b0_0_0_xxxxxxxx_x;
      patterns[924] = 12'b0_0_0_xxxxxxxx_x;
      patterns[925] = 12'b0_1_0_xxxxxxxx_x;
      patterns[926] = 12'b0_0_0_xxxxxxxx_x;
      patterns[927] = 12'b0_0_0_xxxxxxxx_x;
      patterns[928] = 12'b0_1_0_xxxxxxxx_x;
      patterns[929] = 12'b0_0_0_xxxxxxxx_x;
      patterns[930] = 12'b0_0_0_xxxxxxxx_x;
      patterns[931] = 12'b0_1_0_xxxxxxxx_x;
      patterns[932] = 12'b0_0_0_xxxxxxxx_x;
      patterns[933] = 12'b0_0_0_xxxxxxxx_x;
      patterns[934] = 12'b0_1_0_xxxxxxxx_x;
      patterns[935] = 12'b0_0_0_xxxxxxxx_x;
      patterns[936] = 12'b0_0_0_xxxxxxxx_x;
      patterns[937] = 12'b0_1_0_xxxxxxxx_x;
      patterns[938] = 12'b0_0_0_xxxxxxxx_x;
      patterns[939] = 12'b0_0_0_xxxxxxxx_x;
      patterns[940] = 12'b0_1_0_xxxxxxxx_x;
      patterns[941] = 12'b0_0_0_xxxxxxxx_x;
      patterns[942] = 12'b0_0_0_xxxxxxxx_x;
      patterns[943] = 12'b0_1_0_xxxxxxxx_x;
      patterns[944] = 12'b0_0_0_xxxxxxxx_x;
      patterns[945] = 12'b0_0_0_xxxxxxxx_x;
      patterns[946] = 12'b0_1_0_xxxxxxxx_x;
      patterns[947] = 12'b0_0_0_01010101_1;
      patterns[948] = 12'b0_0_0_xxxxxxxx_x;
      patterns[949] = 12'b0_1_0_xxxxxxxx_x;
      patterns[950] = 12'b0_0_0_01010101_1;
      patterns[951] = 12'b0_0_0_xxxxxxxx_x;
      patterns[952] = 12'b0_1_0_xxxxxxxx_x;
      patterns[953] = 12'b0_0_0_01010101_1;
      patterns[954] = 12'b0_0_0_xxxxxxxx_x;
      patterns[955] = 12'b0_1_0_xxxxxxxx_x;
      patterns[956] = 12'b0_0_0_01010101_1;
      patterns[957] = 12'b0_0_0_xxxxxxxx_x;
      patterns[958] = 12'b0_1_0_xxxxxxxx_x;
      patterns[959] = 12'b0_0_0_01010101_1;
      patterns[960] = 12'b0_0_0_xxxxxxxx_x;
      patterns[961] = 12'b0_1_0_xxxxxxxx_x;
      patterns[962] = 12'b0_0_0_01010101_1;
      patterns[963] = 12'b0_0_0_xxxxxxxx_x;
      patterns[964] = 12'b0_1_0_xxxxxxxx_x;
      patterns[965] = 12'b0_0_0_01010101_1;
      patterns[966] = 12'b0_0_0_xxxxxxxx_x;
      patterns[967] = 12'b0_1_0_xxxxxxxx_x;
      patterns[968] = 12'b0_0_0_01010101_1;
      patterns[969] = 12'b0_0_0_xxxxxxxx_x;
      patterns[970] = 12'b0_1_0_xxxxxxxx_x;
      patterns[971] = 12'b0_0_0_01010101_1;
      patterns[972] = 12'b0_0_0_xxxxxxxx_x;
      patterns[973] = 12'b0_1_0_xxxxxxxx_x;
      patterns[974] = 12'b0_0_0_01010101_1;
      patterns[975] = 12'b0_0_0_xxxxxxxx_x;
      patterns[976] = 12'b0_1_0_xxxxxxxx_x;
      patterns[977] = 12'b0_0_0_01010101_1;
      patterns[978] = 12'b0_0_0_xxxxxxxx_x;
      patterns[979] = 12'b0_1_0_xxxxxxxx_x;
      patterns[980] = 12'b0_0_0_01010101_1;
      patterns[981] = 12'b0_0_0_xxxxxxxx_x;
      patterns[982] = 12'b0_1_0_xxxxxxxx_x;
      patterns[983] = 12'b0_0_0_01010101_1;
      patterns[984] = 12'b0_0_0_xxxxxxxx_x;
      patterns[985] = 12'b0_1_0_xxxxxxxx_x;
      patterns[986] = 12'b0_0_0_01010101_1;
      patterns[987] = 12'b0_0_0_xxxxxxxx_x;
      patterns[988] = 12'b0_1_0_xxxxxxxx_x;
      patterns[989] = 12'b0_0_0_01010101_1;
      patterns[990] = 12'b0_0_0_xxxxxxxx_x;
      patterns[991] = 12'b0_1_0_xxxxxxxx_x;
      patterns[992] = 12'b0_0_0_01010101_1;

      for (i = 0; i < 993; i = i + 1)
      begin
        CDP = patterns[i][11];
        clk16 = patterns[i][10];
        RX = patterns[i][9];
        #10;
        if (patterns[i][8:1] !== 8'hx)
        begin
          if (DATA !== patterns[i][8:1])
          begin
            $display("%d:DATA: (assertion error). Expected %h, found %h", i, patterns[i][8:1], DATA);
            $finish;
          end
        end
        if (patterns[i][0] !== 1'hx)
        begin
          if (DP !== patterns[i][0])
          begin
            $display("%d:DP: (assertion error). Expected %h, found %h", i, patterns[i][0], DP);
            $finish;
          end
        end
      end

      $display("All tests passed.");
    end
    endmodule
