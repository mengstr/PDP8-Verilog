`timescale 1us/1ns

module IOTBASEDECODER_tb();
endmodule

